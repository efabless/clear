magic
tech sky130A
magscale 1 2
timestamp 1656242383
<< viali >>
rect 9321 20553 9355 20587
rect 10977 20553 11011 20587
rect 12817 20553 12851 20587
rect 13369 20553 13403 20587
rect 14289 20553 14323 20587
rect 15393 20553 15427 20587
rect 16865 20553 16899 20587
rect 18521 20553 18555 20587
rect 19441 20553 19475 20587
rect 10517 20485 10551 20519
rect 10701 20485 10735 20519
rect 2237 20417 2271 20451
rect 3801 20417 3835 20451
rect 4997 20417 5031 20451
rect 5549 20417 5583 20451
rect 9965 20417 9999 20451
rect 11161 20417 11195 20451
rect 11805 20417 11839 20451
rect 12633 20417 12667 20451
rect 13185 20417 13219 20451
rect 14105 20417 14139 20451
rect 14657 20417 14691 20451
rect 15209 20417 15243 20451
rect 15761 20417 15795 20451
rect 16681 20417 16715 20451
rect 17233 20417 17267 20451
rect 17785 20417 17819 20451
rect 18337 20417 18371 20451
rect 19257 20417 19291 20451
rect 21106 20417 21140 20451
rect 1961 20349 1995 20383
rect 3157 20349 3191 20383
rect 3433 20349 3467 20383
rect 4077 20349 4111 20383
rect 6561 20349 6595 20383
rect 6837 20349 6871 20383
rect 7665 20349 7699 20383
rect 7941 20349 7975 20383
rect 9413 20349 9447 20383
rect 9597 20349 9631 20383
rect 11529 20349 11563 20383
rect 21373 20349 21407 20383
rect 10149 20281 10183 20315
rect 14841 20281 14875 20315
rect 15945 20281 15979 20315
rect 17417 20281 17451 20315
rect 5089 20213 5123 20247
rect 5641 20213 5675 20247
rect 8953 20213 8987 20247
rect 17969 20213 18003 20247
rect 19993 20213 20027 20247
rect 3433 20009 3467 20043
rect 3893 20009 3927 20043
rect 5273 20009 5307 20043
rect 12725 20009 12759 20043
rect 13645 20009 13679 20043
rect 18337 20009 18371 20043
rect 18705 20009 18739 20043
rect 1777 19941 1811 19975
rect 5733 19941 5767 19975
rect 16037 19941 16071 19975
rect 17785 19941 17819 19975
rect 1593 19805 1627 19839
rect 2237 19805 2271 19839
rect 2697 19805 2731 19839
rect 4169 19805 4203 19839
rect 4629 19805 4663 19839
rect 5089 19805 5123 19839
rect 5549 19805 5583 19839
rect 6009 19805 6043 19839
rect 6285 19805 6319 19839
rect 10609 19805 10643 19839
rect 10885 19805 10919 19839
rect 12541 19805 12575 19839
rect 13461 19805 13495 19839
rect 15485 19805 15519 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 17325 19805 17359 19839
rect 17601 19805 17635 19839
rect 18153 19805 18187 19839
rect 18889 19805 18923 19839
rect 19533 19805 19567 19839
rect 21373 19805 21407 19839
rect 2421 19737 2455 19771
rect 7297 19737 7331 19771
rect 7849 19737 7883 19771
rect 8401 19737 8435 19771
rect 8585 19737 8619 19771
rect 10342 19737 10376 19771
rect 11152 19737 11186 19771
rect 13093 19737 13127 19771
rect 15218 19737 15252 19771
rect 19800 19737 19834 19771
rect 2881 19669 2915 19703
rect 4353 19669 4387 19703
rect 4813 19669 4847 19703
rect 7389 19669 7423 19703
rect 7941 19669 7975 19703
rect 9229 19669 9263 19703
rect 12265 19669 12299 19703
rect 14105 19669 14139 19703
rect 16681 19669 16715 19703
rect 17141 19669 17175 19703
rect 20913 19669 20947 19703
rect 21189 19669 21223 19703
rect 1593 19465 1627 19499
rect 4997 19465 5031 19499
rect 5733 19465 5767 19499
rect 6377 19465 6411 19499
rect 6837 19465 6871 19499
rect 8125 19465 8159 19499
rect 11161 19465 11195 19499
rect 11713 19465 11747 19499
rect 12173 19465 12207 19499
rect 12633 19465 12667 19499
rect 14657 19465 14691 19499
rect 18429 19465 18463 19499
rect 18705 19465 18739 19499
rect 4169 19397 4203 19431
rect 10026 19397 10060 19431
rect 15770 19397 15804 19431
rect 19818 19397 19852 19431
rect 1409 19329 1443 19363
rect 4813 19329 4847 19363
rect 5641 19329 5675 19363
rect 6745 19329 6779 19363
rect 7665 19329 7699 19363
rect 9249 19329 9283 19363
rect 11529 19329 11563 19363
rect 11989 19329 12023 19363
rect 12449 19329 12483 19363
rect 14114 19329 14148 19363
rect 16037 19329 16071 19363
rect 17049 19329 17083 19363
rect 17316 19329 17350 19363
rect 20361 19329 20395 19363
rect 2329 19261 2363 19295
rect 2697 19261 2731 19295
rect 3801 19261 3835 19295
rect 5825 19261 5859 19295
rect 7021 19261 7055 19295
rect 9505 19261 9539 19295
rect 9781 19261 9815 19295
rect 14381 19261 14415 19295
rect 20085 19261 20119 19295
rect 20729 19261 20763 19295
rect 3065 19193 3099 19227
rect 3433 19193 3467 19227
rect 1961 19125 1995 19159
rect 4445 19125 4479 19159
rect 5273 19125 5307 19159
rect 7849 19125 7883 19159
rect 13001 19125 13035 19159
rect 16681 19125 16715 19159
rect 1593 18921 1627 18955
rect 3433 18921 3467 18955
rect 6469 18921 6503 18955
rect 11161 18921 11195 18955
rect 1961 18853 1995 18887
rect 3065 18853 3099 18887
rect 6745 18853 6779 18887
rect 8953 18853 8987 18887
rect 2329 18785 2363 18819
rect 4813 18785 4847 18819
rect 16865 18785 16899 18819
rect 20637 18785 20671 18819
rect 4445 18717 4479 18751
rect 5825 18717 5859 18751
rect 6285 18717 6319 18751
rect 6929 18717 6963 18751
rect 8585 18717 8619 18751
rect 10333 18717 10367 18751
rect 10609 18717 10643 18751
rect 10977 18717 11011 18751
rect 12550 18717 12584 18751
rect 12817 18717 12851 18751
rect 13737 18717 13771 18751
rect 14197 18717 14231 18751
rect 14473 18717 14507 18751
rect 14729 18717 14763 18751
rect 16589 18717 16623 18751
rect 18889 18717 18923 18751
rect 21097 18717 21131 18751
rect 2697 18649 2731 18683
rect 3985 18649 4019 18683
rect 5089 18649 5123 18683
rect 5457 18649 5491 18683
rect 8340 18649 8374 18683
rect 10066 18649 10100 18683
rect 17132 18649 17166 18683
rect 20392 18649 20426 18683
rect 6009 18581 6043 18615
rect 7205 18581 7239 18615
rect 11437 18581 11471 18615
rect 13093 18581 13127 18615
rect 13553 18581 13587 18615
rect 15853 18581 15887 18615
rect 16405 18581 16439 18615
rect 18245 18581 18279 18615
rect 18705 18581 18739 18615
rect 19257 18581 19291 18615
rect 21281 18581 21315 18615
rect 1409 18377 1443 18411
rect 1777 18377 1811 18411
rect 2237 18377 2271 18411
rect 3065 18377 3099 18411
rect 3801 18377 3835 18411
rect 5273 18377 5307 18411
rect 5917 18377 5951 18411
rect 6561 18377 6595 18411
rect 7021 18377 7055 18411
rect 7849 18377 7883 18411
rect 8769 18377 8803 18411
rect 12265 18377 12299 18411
rect 15669 18377 15703 18411
rect 2697 18309 2731 18343
rect 3433 18309 3467 18343
rect 5641 18309 5675 18343
rect 21128 18309 21162 18343
rect 4169 18241 4203 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 7941 18241 7975 18275
rect 8585 18241 8619 18275
rect 10158 18241 10192 18275
rect 10425 18241 10459 18275
rect 10701 18241 10735 18275
rect 11621 18241 11655 18275
rect 12081 18241 12115 18275
rect 13654 18241 13688 18275
rect 13921 18241 13955 18275
rect 14289 18241 14323 18275
rect 14545 18241 14579 18275
rect 16037 18241 16071 18275
rect 16681 18241 16715 18275
rect 16937 18241 16971 18275
rect 18337 18241 18371 18275
rect 18593 18241 18627 18275
rect 21373 18241 21407 18275
rect 4905 18173 4939 18207
rect 8125 18173 8159 18207
rect 4537 18105 4571 18139
rect 11805 18105 11839 18139
rect 19717 18105 19751 18139
rect 7481 18037 7515 18071
rect 9045 18037 9079 18071
rect 11069 18037 11103 18071
rect 12541 18037 12575 18071
rect 16221 18037 16255 18071
rect 18061 18037 18095 18071
rect 19993 18037 20027 18071
rect 4169 17833 4203 17867
rect 4445 17833 4479 17867
rect 5549 17833 5583 17867
rect 5917 17833 5951 17867
rect 7021 17833 7055 17867
rect 7941 17833 7975 17867
rect 14841 17833 14875 17867
rect 4905 17765 4939 17799
rect 6745 17765 6779 17799
rect 8401 17765 8435 17799
rect 13737 17765 13771 17799
rect 14289 17765 14323 17799
rect 17141 17765 17175 17799
rect 2053 17697 2087 17731
rect 1685 17629 1719 17663
rect 7205 17629 7239 17663
rect 7757 17629 7791 17663
rect 8217 17629 8251 17663
rect 9781 17629 9815 17663
rect 11529 17629 11563 17663
rect 11805 17629 11839 17663
rect 13553 17629 13587 17663
rect 14105 17629 14139 17663
rect 14657 17629 14691 17663
rect 15117 17629 15151 17663
rect 18521 17629 18555 17663
rect 18797 17629 18831 17663
rect 19625 17629 19659 17663
rect 21373 17629 21407 17663
rect 10026 17561 10060 17595
rect 12050 17561 12084 17595
rect 15373 17561 15407 17595
rect 18254 17561 18288 17595
rect 21128 17561 21162 17595
rect 1501 17493 1535 17527
rect 5181 17493 5215 17527
rect 6285 17493 6319 17527
rect 9045 17493 9079 17527
rect 9413 17493 9447 17527
rect 11161 17493 11195 17527
rect 13185 17493 13219 17527
rect 16497 17493 16531 17527
rect 16865 17493 16899 17527
rect 19441 17493 19475 17527
rect 19993 17493 20027 17527
rect 5549 17289 5583 17323
rect 6929 17289 6963 17323
rect 13461 17289 13495 17323
rect 16221 17289 16255 17323
rect 16865 17289 16899 17323
rect 17969 17289 18003 17323
rect 18429 17289 18463 17323
rect 4997 17153 5031 17187
rect 5641 17153 5675 17187
rect 8033 17153 8067 17187
rect 10158 17153 10192 17187
rect 10425 17153 10459 17187
rect 10701 17153 10735 17187
rect 11069 17153 11103 17187
rect 11713 17153 11747 17187
rect 12081 17153 12115 17187
rect 12449 17153 12483 17187
rect 12817 17153 12851 17187
rect 13277 17153 13311 17187
rect 14850 17153 14884 17187
rect 15117 17153 15151 17187
rect 15577 17153 15611 17187
rect 16037 17153 16071 17187
rect 16681 17153 16715 17187
rect 17233 17153 17267 17187
rect 17785 17153 17819 17187
rect 18613 17153 18647 17187
rect 20013 17153 20047 17187
rect 20545 17153 20579 17187
rect 21097 17153 21131 17187
rect 5457 17085 5491 17119
rect 7665 17085 7699 17119
rect 20269 17085 20303 17119
rect 6469 17017 6503 17051
rect 7205 17017 7239 17051
rect 8309 17017 8343 17051
rect 8677 17017 8711 17051
rect 13001 17017 13035 17051
rect 15761 17017 15795 17051
rect 6009 16949 6043 16983
rect 9045 16949 9079 16983
rect 13737 16949 13771 16983
rect 17417 16949 17451 16983
rect 18889 16949 18923 16983
rect 20729 16949 20763 16983
rect 21281 16949 21315 16983
rect 5365 16745 5399 16779
rect 6009 16745 6043 16779
rect 6837 16745 6871 16779
rect 7665 16745 7699 16779
rect 13737 16745 13771 16779
rect 15485 16677 15519 16711
rect 17141 16677 17175 16711
rect 5641 16609 5675 16643
rect 7205 16609 7239 16643
rect 8125 16609 8159 16643
rect 8217 16609 8251 16643
rect 8953 16609 8987 16643
rect 12449 16609 12483 16643
rect 13277 16609 13311 16643
rect 15761 16609 15795 16643
rect 18889 16609 18923 16643
rect 19257 16609 19291 16643
rect 10701 16541 10735 16575
rect 10968 16541 11002 16575
rect 13553 16541 13587 16575
rect 14105 16541 14139 16575
rect 16017 16541 16051 16575
rect 19513 16541 19547 16575
rect 21097 16541 21131 16575
rect 9198 16473 9232 16507
rect 14350 16473 14384 16507
rect 18622 16473 18656 16507
rect 4537 16405 4571 16439
rect 6377 16405 6411 16439
rect 8033 16405 8067 16439
rect 10333 16405 10367 16439
rect 12081 16405 12115 16439
rect 12817 16405 12851 16439
rect 17509 16405 17543 16439
rect 20637 16405 20671 16439
rect 21281 16405 21315 16439
rect 4169 16201 4203 16235
rect 5273 16201 5307 16235
rect 6653 16201 6687 16235
rect 14933 16201 14967 16235
rect 16129 16201 16163 16235
rect 18061 16201 18095 16235
rect 10342 16133 10376 16167
rect 18766 16133 18800 16167
rect 5181 16065 5215 16099
rect 6745 16065 6779 16099
rect 7573 16065 7607 16099
rect 7829 16065 7863 16099
rect 10609 16065 10643 16099
rect 13010 16065 13044 16099
rect 13277 16065 13311 16099
rect 13553 16065 13587 16099
rect 13820 16065 13854 16099
rect 15209 16065 15243 16099
rect 15853 16065 15887 16099
rect 16313 16065 16347 16099
rect 16681 16065 16715 16099
rect 16948 16065 16982 16099
rect 18521 16065 18555 16099
rect 20545 16065 20579 16099
rect 21097 16065 21131 16099
rect 3985 15997 4019 16031
rect 4077 15997 4111 16031
rect 5457 15997 5491 16031
rect 6561 15997 6595 16031
rect 11897 15929 11931 15963
rect 15393 15929 15427 15963
rect 15669 15929 15703 15963
rect 20177 15929 20211 15963
rect 4537 15861 4571 15895
rect 4813 15861 4847 15895
rect 6009 15861 6043 15895
rect 7113 15861 7147 15895
rect 8953 15861 8987 15895
rect 9229 15861 9263 15895
rect 10977 15861 11011 15895
rect 11621 15861 11655 15895
rect 19901 15861 19935 15895
rect 20729 15861 20763 15895
rect 21281 15861 21315 15895
rect 8953 15657 8987 15691
rect 9321 15657 9355 15691
rect 17693 15657 17727 15691
rect 18245 15657 18279 15691
rect 18705 15657 18739 15691
rect 19625 15657 19659 15691
rect 5825 15589 5859 15623
rect 9781 15589 9815 15623
rect 12081 15589 12115 15623
rect 5273 15521 5307 15555
rect 6745 15521 6779 15555
rect 7205 15521 7239 15555
rect 11161 15521 11195 15555
rect 13461 15521 13495 15555
rect 15577 15521 15611 15555
rect 15853 15521 15887 15555
rect 5457 15453 5491 15487
rect 6469 15453 6503 15487
rect 17509 15453 17543 15487
rect 18429 15453 18463 15487
rect 18889 15453 18923 15487
rect 19441 15453 19475 15487
rect 21373 15453 21407 15487
rect 7472 15385 7506 15419
rect 10894 15385 10928 15419
rect 11529 15385 11563 15419
rect 13194 15385 13228 15419
rect 15310 15385 15344 15419
rect 16098 15385 16132 15419
rect 21106 15385 21140 15419
rect 4629 15317 4663 15351
rect 5365 15317 5399 15351
rect 6101 15317 6135 15351
rect 6561 15317 6595 15351
rect 8585 15317 8619 15351
rect 14197 15317 14231 15351
rect 17233 15317 17267 15351
rect 19993 15317 20027 15351
rect 4905 15113 4939 15147
rect 6561 15113 6595 15147
rect 6837 15113 6871 15147
rect 8217 15113 8251 15147
rect 9045 15113 9079 15147
rect 9321 15113 9355 15147
rect 11069 15113 11103 15147
rect 11621 15113 11655 15147
rect 12081 15113 12115 15147
rect 12449 15113 12483 15147
rect 14933 15113 14967 15147
rect 16865 15113 16899 15147
rect 17325 15113 17359 15147
rect 17969 15113 18003 15147
rect 18705 15113 18739 15147
rect 4997 15045 5031 15079
rect 7297 15045 7331 15079
rect 8125 15045 8159 15079
rect 13277 15045 13311 15079
rect 13645 15045 13679 15079
rect 14289 15045 14323 15079
rect 14657 15045 14691 15079
rect 7205 14977 7239 15011
rect 9689 14977 9723 15011
rect 9945 14977 9979 15011
rect 16046 14977 16080 15011
rect 16313 14977 16347 15011
rect 17049 14977 17083 15011
rect 17509 14977 17543 15011
rect 17785 14977 17819 15011
rect 18429 14977 18463 15011
rect 18889 14977 18923 15011
rect 19165 14977 19199 15011
rect 19717 14977 19751 15011
rect 19973 14977 20007 15011
rect 4813 14909 4847 14943
rect 7481 14909 7515 14943
rect 8033 14909 8067 14943
rect 8585 14841 8619 14875
rect 18245 14841 18279 14875
rect 5365 14773 5399 14807
rect 5917 14773 5951 14807
rect 12817 14773 12851 14807
rect 19349 14773 19383 14807
rect 21097 14773 21131 14807
rect 6929 14569 6963 14603
rect 9229 14569 9263 14603
rect 10977 14569 11011 14603
rect 11529 14569 11563 14603
rect 11897 14569 11931 14603
rect 12265 14569 12299 14603
rect 12633 14569 12667 14603
rect 13737 14569 13771 14603
rect 14105 14569 14139 14603
rect 14473 14569 14507 14603
rect 13277 14501 13311 14535
rect 4169 14433 4203 14467
rect 5181 14433 5215 14467
rect 7481 14433 7515 14467
rect 10609 14433 10643 14467
rect 14841 14433 14875 14467
rect 16486 14433 16520 14467
rect 4261 14365 4295 14399
rect 4353 14365 4387 14399
rect 5365 14365 5399 14399
rect 7389 14365 7423 14399
rect 15097 14365 15131 14399
rect 18429 14365 18463 14399
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 21373 14365 21407 14399
rect 5273 14297 5307 14331
rect 10342 14297 10376 14331
rect 13001 14297 13035 14331
rect 16742 14297 16776 14331
rect 21128 14297 21162 14331
rect 4721 14229 4755 14263
rect 5733 14229 5767 14263
rect 7297 14229 7331 14263
rect 16221 14229 16255 14263
rect 17877 14229 17911 14263
rect 18245 14229 18279 14263
rect 18889 14229 18923 14263
rect 19625 14229 19659 14263
rect 19993 14229 20027 14263
rect 5181 14025 5215 14059
rect 9229 14025 9263 14059
rect 10977 14025 11011 14059
rect 11621 14025 11655 14059
rect 11989 14025 12023 14059
rect 16037 14025 16071 14059
rect 18061 14025 18095 14059
rect 4813 13957 4847 13991
rect 12878 13957 12912 13991
rect 16948 13957 16982 13991
rect 10342 13889 10376 13923
rect 10609 13889 10643 13923
rect 12265 13889 12299 13923
rect 12633 13889 12667 13923
rect 15413 13889 15447 13923
rect 15669 13889 15703 13923
rect 16681 13889 16715 13923
rect 19450 13889 19484 13923
rect 19717 13889 19751 13923
rect 21117 13889 21151 13923
rect 21373 13889 21407 13923
rect 14289 13753 14323 13787
rect 18337 13753 18371 13787
rect 7849 13685 7883 13719
rect 8217 13685 8251 13719
rect 8585 13685 8619 13719
rect 8953 13685 8987 13719
rect 14013 13685 14047 13719
rect 19993 13685 20027 13719
rect 10701 13481 10735 13515
rect 17601 13481 17635 13515
rect 18337 13481 18371 13515
rect 21281 13481 21315 13515
rect 10425 13413 10459 13447
rect 15853 13413 15887 13447
rect 18705 13413 18739 13447
rect 5089 13345 5123 13379
rect 5273 13345 5307 13379
rect 13737 13345 13771 13379
rect 15485 13345 15519 13379
rect 16221 13345 16255 13379
rect 20637 13345 20671 13379
rect 7205 13277 7239 13311
rect 9045 13277 9079 13311
rect 12081 13277 12115 13311
rect 18153 13277 18187 13311
rect 18889 13277 18923 13311
rect 21097 13277 21131 13311
rect 5365 13209 5399 13243
rect 7472 13209 7506 13243
rect 9312 13209 9346 13243
rect 11836 13209 11870 13243
rect 13481 13209 13515 13243
rect 15218 13209 15252 13243
rect 16488 13209 16522 13243
rect 20370 13209 20404 13243
rect 5733 13141 5767 13175
rect 6101 13141 6135 13175
rect 8585 13141 8619 13175
rect 12357 13141 12391 13175
rect 14105 13141 14139 13175
rect 19257 13141 19291 13175
rect 5273 12937 5307 12971
rect 7849 12937 7883 12971
rect 16221 12937 16255 12971
rect 5365 12869 5399 12903
rect 11621 12869 11655 12903
rect 12265 12869 12299 12903
rect 12633 12869 12667 12903
rect 17794 12869 17828 12903
rect 21106 12869 21140 12903
rect 6469 12801 6503 12835
rect 6725 12801 6759 12835
rect 8125 12801 8159 12835
rect 8392 12801 8426 12835
rect 9781 12801 9815 12835
rect 10048 12801 10082 12835
rect 14033 12801 14067 12835
rect 14289 12801 14323 12835
rect 15678 12801 15712 12835
rect 15945 12801 15979 12835
rect 18061 12801 18095 12835
rect 18337 12801 18371 12835
rect 18604 12801 18638 12835
rect 21373 12801 21407 12835
rect 5181 12733 5215 12767
rect 5733 12665 5767 12699
rect 9505 12665 9539 12699
rect 19717 12665 19751 12699
rect 11161 12597 11195 12631
rect 12909 12597 12943 12631
rect 14565 12597 14599 12631
rect 16681 12597 16715 12631
rect 19993 12597 20027 12631
rect 10517 12393 10551 12427
rect 13001 12393 13035 12427
rect 13369 12393 13403 12427
rect 13737 12393 13771 12427
rect 14105 12393 14139 12427
rect 19533 12393 19567 12427
rect 5549 12325 5583 12359
rect 8585 12325 8619 12359
rect 17417 12325 17451 12359
rect 6653 12257 6687 12291
rect 6837 12257 6871 12291
rect 15485 12257 15519 12291
rect 17141 12257 17175 12291
rect 18797 12257 18831 12291
rect 7205 12189 7239 12223
rect 9137 12189 9171 12223
rect 9393 12189 9427 12223
rect 10885 12189 10919 12223
rect 11253 12189 11287 12223
rect 11509 12189 11543 12223
rect 16874 12189 16908 12223
rect 19717 12189 19751 12223
rect 21373 12189 21407 12223
rect 5917 12121 5951 12155
rect 7472 12121 7506 12155
rect 15218 12121 15252 12155
rect 18530 12121 18564 12155
rect 21128 12121 21162 12155
rect 6193 12053 6227 12087
rect 6561 12053 6595 12087
rect 12633 12053 12667 12087
rect 15761 12053 15795 12087
rect 19993 12053 20027 12087
rect 7021 11849 7055 11883
rect 8125 11849 8159 11883
rect 11621 11849 11655 11883
rect 12909 11849 12943 11883
rect 14381 11849 14415 11883
rect 15577 11849 15611 11883
rect 17049 11849 17083 11883
rect 17693 11849 17727 11883
rect 5641 11781 5675 11815
rect 8493 11781 8527 11815
rect 10885 11781 10919 11815
rect 19625 11781 19659 11815
rect 20238 11781 20272 11815
rect 7389 11713 7423 11747
rect 10353 11713 10387 11747
rect 11897 11713 11931 11747
rect 12265 11713 12299 11747
rect 13277 11713 13311 11747
rect 14749 11713 14783 11747
rect 16313 11713 16347 11747
rect 17233 11713 17267 11747
rect 17509 11713 17543 11747
rect 17969 11713 18003 11747
rect 18236 11713 18270 11747
rect 19993 11713 20027 11747
rect 5457 11645 5491 11679
rect 5549 11645 5583 11679
rect 6745 11645 6779 11679
rect 7481 11645 7515 11679
rect 7665 11645 7699 11679
rect 8585 11645 8619 11679
rect 8769 11645 8803 11679
rect 10609 11645 10643 11679
rect 13369 11645 13403 11679
rect 13461 11645 13495 11679
rect 13921 11645 13955 11679
rect 14841 11645 14875 11679
rect 14933 11645 14967 11679
rect 16681 11577 16715 11611
rect 4905 11509 4939 11543
rect 6009 11509 6043 11543
rect 9229 11509 9263 11543
rect 16129 11509 16163 11543
rect 19349 11509 19383 11543
rect 21373 11509 21407 11543
rect 6561 11305 6595 11339
rect 7573 11305 7607 11339
rect 7849 11305 7883 11339
rect 14933 11305 14967 11339
rect 15209 11305 15243 11339
rect 16405 11305 16439 11339
rect 17049 11305 17083 11339
rect 18797 11305 18831 11339
rect 9505 11237 9539 11271
rect 12173 11237 12207 11271
rect 19257 11237 19291 11271
rect 5917 11169 5951 11203
rect 6101 11169 6135 11203
rect 7021 11169 7055 11203
rect 8401 11169 8435 11203
rect 11621 11169 11655 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 14381 11169 14415 11203
rect 15761 11169 15795 11203
rect 17877 11169 17911 11203
rect 19901 11169 19935 11203
rect 20821 11169 20855 11203
rect 21281 11169 21315 11203
rect 7205 11101 7239 11135
rect 10885 11101 10919 11135
rect 12817 11101 12851 11135
rect 14473 11101 14507 11135
rect 16865 11101 16899 11135
rect 5549 11033 5583 11067
rect 6193 11033 6227 11067
rect 7113 11033 7147 11067
rect 8217 11033 8251 11067
rect 8953 11033 8987 11067
rect 10640 11033 10674 11067
rect 15577 11033 15611 11067
rect 19625 11033 19659 11067
rect 19717 11033 19751 11067
rect 20729 11033 20763 11067
rect 8309 10965 8343 10999
rect 11713 10965 11747 10999
rect 11805 10965 11839 10999
rect 12449 10965 12483 10999
rect 13461 10965 13495 10999
rect 14565 10965 14599 10999
rect 15669 10965 15703 10999
rect 17325 10965 17359 10999
rect 17693 10965 17727 10999
rect 17785 10965 17819 10999
rect 18337 10965 18371 10999
rect 20269 10965 20303 10999
rect 20637 10965 20671 10999
rect 7389 10761 7423 10795
rect 8309 10761 8343 10795
rect 9413 10761 9447 10795
rect 11161 10761 11195 10795
rect 12357 10761 12391 10795
rect 12817 10761 12851 10795
rect 13737 10761 13771 10795
rect 14381 10761 14415 10795
rect 16865 10761 16899 10795
rect 17141 10761 17175 10795
rect 18337 10761 18371 10795
rect 18705 10761 18739 10795
rect 19533 10761 19567 10795
rect 20269 10761 20303 10795
rect 21373 10761 21407 10795
rect 9873 10693 9907 10727
rect 11989 10693 12023 10727
rect 12725 10693 12759 10727
rect 14749 10693 14783 10727
rect 15669 10693 15703 10727
rect 19625 10693 19659 10727
rect 6745 10625 6779 10659
rect 8677 10625 8711 10659
rect 9781 10625 9815 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 15945 10625 15979 10659
rect 16681 10625 16715 10659
rect 17509 10625 17543 10659
rect 20637 10625 20671 10659
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 8769 10557 8803 10591
rect 8953 10557 8987 10591
rect 10057 10557 10091 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 12909 10557 12943 10591
rect 13553 10557 13587 10591
rect 13645 10557 13679 10591
rect 14841 10557 14875 10591
rect 15025 10557 15059 10591
rect 18061 10557 18095 10591
rect 18245 10557 18279 10591
rect 19441 10557 19475 10591
rect 20729 10557 20763 10591
rect 20821 10557 20855 10591
rect 7113 10489 7147 10523
rect 16129 10489 16163 10523
rect 5917 10421 5951 10455
rect 8033 10421 8067 10455
rect 14105 10421 14139 10455
rect 17693 10421 17727 10455
rect 19993 10421 20027 10455
rect 13093 10217 13127 10251
rect 14197 10217 14231 10251
rect 14841 10217 14875 10251
rect 17693 10217 17727 10251
rect 20821 10217 20855 10251
rect 21281 10217 21315 10251
rect 6377 10149 6411 10183
rect 7389 10149 7423 10183
rect 10885 10149 10919 10183
rect 13737 10149 13771 10183
rect 17325 10149 17359 10183
rect 5457 10081 5491 10115
rect 6929 10081 6963 10115
rect 9229 10081 9263 10115
rect 10241 10081 10275 10115
rect 12541 10081 12575 10115
rect 15761 10081 15795 10115
rect 16405 10081 16439 10115
rect 18153 10081 18187 10115
rect 18337 10081 18371 10115
rect 20361 10081 20395 10115
rect 6745 10013 6779 10047
rect 6837 10013 6871 10047
rect 9505 10013 9539 10047
rect 11621 10013 11655 10047
rect 12725 10013 12759 10047
rect 15485 10013 15519 10047
rect 17141 10013 17175 10047
rect 18889 10013 18923 10047
rect 19257 10013 19291 10047
rect 19717 10013 19751 10047
rect 21005 10013 21039 10047
rect 7757 9945 7791 9979
rect 8585 9945 8619 9979
rect 10517 9945 10551 9979
rect 11161 9945 11195 9979
rect 18061 9945 18095 9979
rect 5641 9877 5675 9911
rect 5733 9877 5767 9911
rect 6101 9877 6135 9911
rect 8125 9877 8159 9911
rect 9413 9877 9447 9911
rect 9873 9877 9907 9911
rect 10425 9877 10459 9911
rect 12633 9877 12667 9911
rect 15117 9877 15151 9911
rect 15577 9877 15611 9911
rect 16865 9877 16899 9911
rect 18705 9877 18739 9911
rect 19441 9877 19475 9911
rect 19901 9877 19935 9911
rect 6745 9673 6779 9707
rect 7113 9673 7147 9707
rect 7665 9673 7699 9707
rect 10241 9673 10275 9707
rect 10885 9673 10919 9707
rect 14749 9673 14783 9707
rect 17049 9673 17083 9707
rect 18429 9673 18463 9707
rect 18705 9673 18739 9707
rect 19901 9673 19935 9707
rect 6653 9605 6687 9639
rect 8677 9605 8711 9639
rect 11621 9605 11655 9639
rect 13645 9605 13679 9639
rect 20637 9605 20671 9639
rect 4997 9537 5031 9571
rect 5641 9537 5675 9571
rect 7757 9537 7791 9571
rect 8769 9537 8803 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 15669 9537 15703 9571
rect 17969 9537 18003 9571
rect 18061 9537 18095 9571
rect 18889 9537 18923 9571
rect 19441 9537 19475 9571
rect 19717 9537 19751 9571
rect 20545 9537 20579 9571
rect 21373 9537 21407 9571
rect 5457 9469 5491 9503
rect 5549 9469 5583 9503
rect 6561 9469 6595 9503
rect 7573 9469 7607 9503
rect 8493 9469 8527 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 12633 9469 12667 9503
rect 12817 9469 12851 9503
rect 13829 9469 13863 9503
rect 14933 9469 14967 9503
rect 15393 9469 15427 9503
rect 15577 9469 15611 9503
rect 16865 9469 16899 9503
rect 16957 9469 16991 9503
rect 17785 9469 17819 9503
rect 20729 9469 20763 9503
rect 4629 9401 4663 9435
rect 8125 9401 8159 9435
rect 9137 9401 9171 9435
rect 12173 9401 12207 9435
rect 13185 9401 13219 9435
rect 16037 9401 16071 9435
rect 19257 9401 19291 9435
rect 21189 9401 21223 9435
rect 6009 9333 6043 9367
rect 9505 9333 9539 9367
rect 10609 9333 10643 9367
rect 14289 9333 14323 9367
rect 17417 9333 17451 9367
rect 20177 9333 20211 9367
rect 5917 9129 5951 9163
rect 9965 9129 9999 9163
rect 10701 9129 10735 9163
rect 11069 9129 11103 9163
rect 11621 9129 11655 9163
rect 14197 9129 14231 9163
rect 15117 9129 15151 9163
rect 18429 9129 18463 9163
rect 20453 9129 20487 9163
rect 20177 9061 20211 9095
rect 5365 8993 5399 9027
rect 6929 8993 6963 9027
rect 7113 8993 7147 9027
rect 7849 8993 7883 9027
rect 9413 8993 9447 9027
rect 12449 8993 12483 9027
rect 13277 8993 13311 9027
rect 15945 8993 15979 9027
rect 17877 8993 17911 9027
rect 19717 8993 19751 9027
rect 21005 8993 21039 9027
rect 5549 8925 5583 8959
rect 7205 8925 7239 8959
rect 12357 8925 12391 8959
rect 13645 8925 13679 8959
rect 16865 8925 16899 8959
rect 18705 8925 18739 8959
rect 19993 8925 20027 8959
rect 5457 8857 5491 8891
rect 9505 8857 9539 8891
rect 16037 8857 16071 8891
rect 20913 8857 20947 8891
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 9597 8789 9631 8823
rect 10333 8789 10367 8823
rect 11897 8789 11931 8823
rect 12265 8789 12299 8823
rect 14565 8789 14599 8823
rect 16129 8789 16163 8823
rect 16497 8789 16531 8823
rect 17049 8789 17083 8823
rect 17417 8789 17451 8823
rect 17969 8789 18003 8823
rect 18061 8789 18095 8823
rect 18889 8789 18923 8823
rect 20821 8789 20855 8823
rect 7297 8585 7331 8619
rect 10149 8585 10183 8619
rect 11621 8585 11655 8619
rect 12265 8585 12299 8619
rect 12725 8585 12759 8619
rect 16313 8585 16347 8619
rect 16957 8585 16991 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 18153 8585 18187 8619
rect 20637 8585 20671 8619
rect 10517 8517 10551 8551
rect 21097 8517 21131 8551
rect 9505 8449 9539 8483
rect 13093 8449 13127 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 15025 8449 15059 8483
rect 16129 8449 16163 8483
rect 17693 8449 17727 8483
rect 18521 8449 18555 8483
rect 18613 8449 18647 8483
rect 19165 8449 19199 8483
rect 19901 8449 19935 8483
rect 20361 8449 20395 8483
rect 21005 8449 21039 8483
rect 5273 8381 5307 8415
rect 6377 8381 6411 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10609 8381 10643 8415
rect 10701 8381 10735 8415
rect 13553 8381 13587 8415
rect 14473 8381 14507 8415
rect 15577 8381 15611 8415
rect 16865 8381 16899 8415
rect 18705 8381 18739 8415
rect 21281 8381 21315 8415
rect 6929 8313 6963 8347
rect 11989 8313 12023 8347
rect 19349 8313 19383 8347
rect 20177 8313 20211 8347
rect 8033 8245 8067 8279
rect 9137 8245 9171 8279
rect 14105 8245 14139 8279
rect 19717 8245 19751 8279
rect 6837 8041 6871 8075
rect 8953 8041 8987 8075
rect 10057 8041 10091 8075
rect 10885 8041 10919 8075
rect 12909 8041 12943 8075
rect 13277 8041 13311 8075
rect 15393 8041 15427 8075
rect 18061 8041 18095 8075
rect 19901 8041 19935 8075
rect 20361 8041 20395 8075
rect 21281 8041 21315 8075
rect 21005 7973 21039 8007
rect 5273 7905 5307 7939
rect 6193 7905 6227 7939
rect 6377 7905 6411 7939
rect 9413 7905 9447 7939
rect 9505 7905 9539 7939
rect 11345 7905 11379 7939
rect 11529 7905 11563 7939
rect 12357 7905 12391 7939
rect 14289 7905 14323 7939
rect 17233 7905 17267 7939
rect 18705 7905 18739 7939
rect 5457 7837 5491 7871
rect 8585 7837 8619 7871
rect 12541 7837 12575 7871
rect 17049 7837 17083 7871
rect 20085 7837 20119 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 9321 7769 9355 7803
rect 10609 7769 10643 7803
rect 16957 7769 16991 7803
rect 19257 7769 19291 7803
rect 4721 7701 4755 7735
rect 5365 7701 5399 7735
rect 5825 7701 5859 7735
rect 6469 7701 6503 7735
rect 7113 7701 7147 7735
rect 11253 7701 11287 7735
rect 12449 7701 12483 7735
rect 13645 7701 13679 7735
rect 14381 7701 14415 7735
rect 14473 7701 14507 7735
rect 14841 7701 14875 7735
rect 15669 7701 15703 7735
rect 16037 7701 16071 7735
rect 16589 7701 16623 7735
rect 17601 7701 17635 7735
rect 18429 7701 18463 7735
rect 18521 7701 18555 7735
rect 5273 7497 5307 7531
rect 5641 7497 5675 7531
rect 6745 7497 6779 7531
rect 8033 7497 8067 7531
rect 8401 7497 8435 7531
rect 9781 7497 9815 7531
rect 11529 7497 11563 7531
rect 11989 7497 12023 7531
rect 13921 7497 13955 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 15669 7497 15703 7531
rect 16313 7497 16347 7531
rect 17049 7497 17083 7531
rect 18245 7497 18279 7531
rect 18613 7497 18647 7531
rect 18889 7497 18923 7531
rect 19809 7497 19843 7531
rect 20269 7497 20303 7531
rect 20913 7497 20947 7531
rect 6009 7429 6043 7463
rect 6653 7429 6687 7463
rect 9321 7429 9355 7463
rect 14473 7429 14507 7463
rect 18153 7429 18187 7463
rect 9413 7361 9447 7395
rect 10057 7361 10091 7395
rect 11069 7361 11103 7395
rect 11897 7361 11931 7395
rect 13553 7361 13587 7395
rect 15577 7361 15611 7395
rect 19073 7361 19107 7395
rect 19349 7361 19383 7395
rect 19993 7361 20027 7395
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 21373 7361 21407 7395
rect 4997 7293 5031 7327
rect 5181 7293 5215 7327
rect 6561 7293 6595 7327
rect 9137 7293 9171 7327
rect 12081 7293 12115 7327
rect 13277 7293 13311 7327
rect 13461 7293 13495 7327
rect 14381 7293 14415 7327
rect 15853 7293 15887 7327
rect 16773 7293 16807 7327
rect 16957 7293 16991 7327
rect 18061 7293 18095 7327
rect 7113 7225 7147 7259
rect 8769 7225 8803 7259
rect 12541 7225 12575 7259
rect 17417 7225 17451 7259
rect 19533 7225 19567 7259
rect 4537 7157 4571 7191
rect 10701 7157 10735 7191
rect 15209 7157 15243 7191
rect 21189 7157 21223 7191
rect 11437 6953 11471 6987
rect 13645 6953 13679 6987
rect 15577 6953 15611 6987
rect 17325 6953 17359 6987
rect 18613 6953 18647 6987
rect 20453 6953 20487 6987
rect 10425 6885 10459 6919
rect 10701 6885 10735 6919
rect 20729 6885 20763 6919
rect 7849 6817 7883 6851
rect 8217 6817 8251 6851
rect 11989 6817 12023 6851
rect 14749 6817 14783 6851
rect 15209 6817 15243 6851
rect 16221 6817 16255 6851
rect 16773 6817 16807 6851
rect 18061 6817 18095 6851
rect 9137 6749 9171 6783
rect 9505 6749 9539 6783
rect 15945 6749 15979 6783
rect 16865 6749 16899 6783
rect 18245 6749 18279 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 20269 6749 20303 6783
rect 20913 6749 20947 6783
rect 21373 6749 21407 6783
rect 8585 6681 8619 6715
rect 11069 6681 11103 6715
rect 12081 6681 12115 6715
rect 14473 6681 14507 6715
rect 9781 6613 9815 6647
rect 12173 6613 12207 6647
rect 12541 6613 12575 6647
rect 13001 6613 13035 6647
rect 13369 6613 13403 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 16037 6613 16071 6647
rect 16957 6613 16991 6647
rect 18153 6613 18187 6647
rect 19349 6613 19383 6647
rect 19993 6613 20027 6647
rect 21189 6613 21223 6647
rect 8401 6409 8435 6443
rect 9505 6409 9539 6443
rect 10057 6409 10091 6443
rect 12173 6409 12207 6443
rect 14473 6409 14507 6443
rect 14565 6409 14599 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 18061 6409 18095 6443
rect 18153 6409 18187 6443
rect 19901 6409 19935 6443
rect 21005 6409 21039 6443
rect 21097 6409 21131 6443
rect 9045 6341 9079 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 9137 6273 9171 6307
rect 10149 6273 10183 6307
rect 11161 6273 11195 6307
rect 13185 6273 13219 6307
rect 15485 6273 15519 6307
rect 16313 6273 16347 6307
rect 18981 6273 19015 6307
rect 19441 6273 19475 6307
rect 19717 6273 19751 6307
rect 20361 6273 20395 6307
rect 8861 6205 8895 6239
rect 9965 6205 9999 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 13277 6205 13311 6239
rect 13369 6205 13403 6239
rect 14657 6205 14691 6239
rect 15209 6205 15243 6239
rect 15393 6205 15427 6239
rect 17141 6205 17175 6239
rect 17325 6205 17359 6239
rect 18245 6205 18279 6239
rect 21189 6205 21223 6239
rect 1593 6137 1627 6171
rect 8125 6137 8159 6171
rect 12541 6137 12575 6171
rect 12817 6137 12851 6171
rect 16129 6137 16163 6171
rect 20177 6137 20211 6171
rect 10517 6069 10551 6103
rect 14105 6069 14139 6103
rect 15853 6069 15887 6103
rect 17693 6069 17727 6103
rect 18797 6069 18831 6103
rect 19257 6069 19291 6103
rect 20637 6069 20671 6103
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 10057 5865 10091 5899
rect 10425 5865 10459 5899
rect 11897 5865 11931 5899
rect 15945 5865 15979 5899
rect 16957 5865 16991 5899
rect 12909 5797 12943 5831
rect 14197 5797 14231 5831
rect 9413 5729 9447 5763
rect 10793 5729 10827 5763
rect 12449 5729 12483 5763
rect 13461 5729 13495 5763
rect 15577 5729 15611 5763
rect 16405 5729 16439 5763
rect 16589 5729 16623 5763
rect 17601 5729 17635 5763
rect 18337 5729 18371 5763
rect 19717 5729 19751 5763
rect 21097 5729 21131 5763
rect 9597 5661 9631 5695
rect 11069 5661 11103 5695
rect 12265 5661 12299 5695
rect 13277 5661 13311 5695
rect 15301 5661 15335 5695
rect 16313 5661 16347 5695
rect 17325 5661 17359 5695
rect 19901 5661 19935 5695
rect 21005 5661 21039 5695
rect 10977 5593 11011 5627
rect 12357 5593 12391 5627
rect 14657 5593 14691 5627
rect 18429 5593 18463 5627
rect 18521 5593 18555 5627
rect 9689 5525 9723 5559
rect 11437 5525 11471 5559
rect 13369 5525 13403 5559
rect 14933 5525 14967 5559
rect 15393 5525 15427 5559
rect 17417 5525 17451 5559
rect 18889 5525 18923 5559
rect 19809 5525 19843 5559
rect 20269 5525 20303 5559
rect 20545 5525 20579 5559
rect 20913 5525 20947 5559
rect 8401 5321 8435 5355
rect 8769 5321 8803 5355
rect 9505 5321 9539 5355
rect 10609 5321 10643 5355
rect 11069 5321 11103 5355
rect 11713 5321 11747 5355
rect 13461 5321 13495 5355
rect 14841 5321 14875 5355
rect 14933 5321 14967 5355
rect 17785 5321 17819 5355
rect 18337 5321 18371 5355
rect 18705 5321 18739 5355
rect 19717 5321 19751 5355
rect 20729 5321 20763 5355
rect 8125 5253 8159 5287
rect 12081 5253 12115 5287
rect 20821 5253 20855 5287
rect 9873 5185 9907 5219
rect 13553 5185 13587 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16681 5185 16715 5219
rect 17693 5185 17727 5219
rect 9965 5117 9999 5151
rect 10149 5117 10183 5151
rect 12173 5117 12207 5151
rect 12357 5117 12391 5151
rect 12909 5117 12943 5151
rect 13277 5117 13311 5151
rect 14749 5117 14783 5151
rect 15761 5117 15795 5151
rect 17877 5117 17911 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 19809 5117 19843 5151
rect 19901 5117 19935 5151
rect 21005 5117 21039 5151
rect 9137 5049 9171 5083
rect 14197 5049 14231 5083
rect 16865 5049 16899 5083
rect 19349 5049 19383 5083
rect 13921 4981 13955 5015
rect 15301 4981 15335 5015
rect 16313 4981 16347 5015
rect 17325 4981 17359 5015
rect 20361 4981 20395 5015
rect 9505 4777 9539 4811
rect 10609 4777 10643 4811
rect 14105 4777 14139 4811
rect 17877 4777 17911 4811
rect 7849 4709 7883 4743
rect 19993 4709 20027 4743
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 11161 4641 11195 4675
rect 12173 4641 12207 4675
rect 13185 4641 13219 4675
rect 14657 4641 14691 4675
rect 15577 4641 15611 4675
rect 15761 4641 15795 4675
rect 18337 4641 18371 4675
rect 18521 4641 18555 4675
rect 19717 4641 19751 4675
rect 20821 4641 20855 4675
rect 8585 4573 8619 4607
rect 9045 4573 9079 4607
rect 9873 4573 9907 4607
rect 12081 4573 12115 4607
rect 13001 4573 13035 4607
rect 15485 4573 15519 4607
rect 16405 4573 16439 4607
rect 16865 4573 16899 4607
rect 17325 4573 17359 4607
rect 20545 4573 20579 4607
rect 8217 4505 8251 4539
rect 11069 4505 11103 4539
rect 11989 4505 12023 4539
rect 13093 4505 13127 4539
rect 20177 4505 20211 4539
rect 9229 4437 9263 4471
rect 10977 4437 11011 4471
rect 11621 4437 11655 4471
rect 12633 4437 12667 4471
rect 13737 4437 13771 4471
rect 14473 4437 14507 4471
rect 14565 4437 14599 4471
rect 15117 4437 15151 4471
rect 16589 4437 16623 4471
rect 17049 4437 17083 4471
rect 17509 4437 17543 4471
rect 18245 4437 18279 4471
rect 10425 4233 10459 4267
rect 11161 4233 11195 4267
rect 12265 4233 12299 4267
rect 13001 4233 13035 4267
rect 14197 4233 14231 4267
rect 15761 4233 15795 4267
rect 18245 4233 18279 4267
rect 18705 4233 18739 4267
rect 9689 4165 9723 4199
rect 11897 4165 11931 4199
rect 13369 4165 13403 4199
rect 15117 4165 15151 4199
rect 20177 4165 20211 4199
rect 8585 4097 8619 4131
rect 10701 4097 10735 4131
rect 11805 4097 11839 4131
rect 12725 4097 12759 4131
rect 14473 4097 14507 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17785 4097 17819 4131
rect 18889 4097 18923 4131
rect 19441 4097 19475 4131
rect 20545 4097 20579 4131
rect 20821 4097 20855 4131
rect 8861 4029 8895 4063
rect 10057 4029 10091 4063
rect 11713 4029 11747 4063
rect 13461 4029 13495 4063
rect 13553 4029 13587 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 7481 3961 7515 3995
rect 16865 3961 16899 3995
rect 19625 3961 19659 3995
rect 1409 3893 1443 3927
rect 7849 3893 7883 3927
rect 8125 3893 8159 3927
rect 9229 3893 9263 3927
rect 12541 3893 12575 3927
rect 14657 3893 14691 3927
rect 16129 3893 16163 3927
rect 17509 3893 17543 3927
rect 17969 3893 18003 3927
rect 20085 3893 20119 3927
rect 1593 3689 1627 3723
rect 7113 3689 7147 3723
rect 18245 3689 18279 3723
rect 7849 3621 7883 3655
rect 9873 3621 9907 3655
rect 10517 3621 10551 3655
rect 10977 3621 11011 3655
rect 19625 3621 19659 3655
rect 7481 3553 7515 3587
rect 14841 3553 14875 3587
rect 15761 3553 15795 3587
rect 16681 3553 16715 3587
rect 16773 3553 16807 3587
rect 19993 3553 20027 3587
rect 1409 3485 1443 3519
rect 1869 3485 1903 3519
rect 8493 3485 8527 3519
rect 9505 3485 9539 3519
rect 11345 3485 11379 3519
rect 11805 3485 11839 3519
rect 12265 3485 12299 3519
rect 12725 3485 12759 3519
rect 13185 3485 13219 3519
rect 16589 3485 16623 3519
rect 17601 3485 17635 3519
rect 18061 3485 18095 3519
rect 18521 3485 18555 3519
rect 19441 3485 19475 3519
rect 20545 3485 20579 3519
rect 20821 3485 20855 3519
rect 2237 3417 2271 3451
rect 6745 3417 6779 3451
rect 9137 3417 9171 3451
rect 13645 3417 13679 3451
rect 14565 3417 14599 3451
rect 20177 3417 20211 3451
rect 4261 3349 4295 3383
rect 4813 3349 4847 3383
rect 5365 3349 5399 3383
rect 6101 3349 6135 3383
rect 8217 3349 8251 3383
rect 10149 3349 10183 3383
rect 11529 3349 11563 3383
rect 11989 3349 12023 3383
rect 12449 3349 12483 3383
rect 12909 3349 12943 3383
rect 13369 3349 13403 3383
rect 14197 3349 14231 3383
rect 14657 3349 14691 3383
rect 15209 3349 15243 3383
rect 15577 3349 15611 3383
rect 15669 3349 15703 3383
rect 16221 3349 16255 3383
rect 17233 3349 17267 3383
rect 17785 3349 17819 3383
rect 18705 3349 18739 3383
rect 1777 3145 1811 3179
rect 9505 3145 9539 3179
rect 11805 3145 11839 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 14841 3145 14875 3179
rect 15301 3145 15335 3179
rect 18981 3145 19015 3179
rect 5549 3077 5583 3111
rect 5733 3077 5767 3111
rect 9045 3077 9079 3111
rect 15209 3077 15243 3111
rect 1593 3009 1627 3043
rect 4077 3009 4111 3043
rect 4905 3009 4939 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9321 3009 9355 3043
rect 9873 3009 9907 3043
rect 10977 3009 11011 3043
rect 11621 3009 11655 3043
rect 12081 3009 12115 3043
rect 12541 3009 12575 3043
rect 13001 3009 13035 3043
rect 13461 3009 13495 3043
rect 16037 3009 16071 3043
rect 16865 3009 16899 3043
rect 17141 3009 17175 3043
rect 17601 3009 17635 3043
rect 18153 3009 18187 3043
rect 19073 3009 19107 3043
rect 19441 3009 19475 3043
rect 19993 3009 20027 3043
rect 20545 3009 20579 3043
rect 20821 3009 20855 3043
rect 3525 2941 3559 2975
rect 3801 2941 3835 2975
rect 10241 2941 10275 2975
rect 10609 2941 10643 2975
rect 14289 2941 14323 2975
rect 14381 2941 14415 2975
rect 15485 2941 15519 2975
rect 5089 2873 5123 2907
rect 7205 2873 7239 2907
rect 8677 2873 8711 2907
rect 11161 2873 11195 2907
rect 17785 2873 17819 2907
rect 19625 2873 19659 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 3157 2805 3191 2839
rect 6469 2805 6503 2839
rect 6837 2805 6871 2839
rect 7941 2805 7975 2839
rect 12265 2805 12299 2839
rect 12725 2805 12759 2839
rect 13185 2805 13219 2839
rect 15853 2805 15887 2839
rect 16681 2805 16715 2839
rect 17325 2805 17359 2839
rect 18337 2805 18371 2839
rect 20177 2805 20211 2839
rect 6745 2601 6779 2635
rect 7849 2601 7883 2635
rect 8401 2601 8435 2635
rect 10609 2601 10643 2635
rect 11161 2601 11195 2635
rect 17969 2601 18003 2635
rect 3249 2533 3283 2567
rect 10149 2533 10183 2567
rect 11805 2533 11839 2567
rect 14749 2533 14783 2567
rect 15945 2533 15979 2567
rect 18521 2533 18555 2567
rect 19993 2533 20027 2567
rect 21097 2533 21131 2567
rect 4077 2465 4111 2499
rect 4629 2465 4663 2499
rect 5733 2465 5767 2499
rect 9229 2465 9263 2499
rect 9597 2465 9631 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 7113 2397 7147 2431
rect 9045 2397 9079 2431
rect 9965 2397 9999 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 11621 2397 11655 2431
rect 12081 2397 12115 2431
rect 12633 2397 12667 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 15209 2397 15243 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 19257 2397 19291 2431
rect 19809 2397 19843 2431
rect 20361 2397 20395 2431
rect 20913 2397 20947 2431
rect 2605 2329 2639 2363
rect 3893 2329 3927 2363
rect 5917 2329 5951 2363
rect 6653 2329 6687 2363
rect 7757 2329 7791 2363
rect 8309 2329 8343 2363
rect 2697 2261 2731 2295
rect 7297 2261 7331 2295
rect 12265 2261 12299 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 19441 2261 19475 2295
rect 20545 2261 20579 2295
<< metal1 >>
rect 14550 20816 14556 20868
rect 14608 20856 14614 20868
rect 17954 20856 17960 20868
rect 14608 20828 17960 20856
rect 14608 20816 14614 20828
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 2314 20748 2320 20800
rect 2372 20788 2378 20800
rect 20346 20788 20352 20800
rect 2372 20760 20352 20788
rect 2372 20748 2378 20760
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 9309 20587 9367 20593
rect 9309 20553 9321 20587
rect 9355 20584 9367 20587
rect 10965 20587 11023 20593
rect 10965 20584 10977 20587
rect 9355 20556 10977 20584
rect 9355 20553 9367 20556
rect 9309 20547 9367 20553
rect 10965 20553 10977 20556
rect 11011 20553 11023 20587
rect 10965 20547 11023 20553
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12805 20587 12863 20593
rect 12805 20584 12817 20587
rect 12584 20556 12817 20584
rect 12584 20544 12590 20556
rect 12805 20553 12817 20556
rect 12851 20553 12863 20587
rect 12805 20547 12863 20553
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 13136 20556 13369 20584
rect 13136 20544 13142 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 13357 20547 13415 20553
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13872 20556 14289 20584
rect 13872 20544 13878 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 14792 20556 15393 20584
rect 14792 20544 14798 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 15896 20556 16865 20584
rect 15896 20544 15902 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 18509 20587 18567 20593
rect 18509 20584 18521 20587
rect 17552 20556 18521 20584
rect 17552 20544 17558 20556
rect 18509 20553 18521 20556
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 18656 20556 19441 20584
rect 18656 20544 18662 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 10318 20516 10324 20528
rect 3936 20488 10324 20516
rect 3936 20476 3942 20488
rect 10318 20476 10324 20488
rect 10376 20516 10382 20528
rect 10505 20519 10563 20525
rect 10505 20516 10517 20519
rect 10376 20488 10517 20516
rect 10376 20476 10382 20488
rect 10505 20485 10517 20488
rect 10551 20485 10563 20519
rect 10505 20479 10563 20485
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20516 10747 20519
rect 11698 20516 11704 20528
rect 10735 20488 11704 20516
rect 10735 20485 10747 20488
rect 10689 20479 10747 20485
rect 11698 20476 11704 20488
rect 11756 20476 11762 20528
rect 11900 20488 12664 20516
rect 382 20408 388 20460
rect 440 20448 446 20460
rect 2222 20448 2228 20460
rect 440 20420 2228 20448
rect 440 20408 446 20420
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 3050 20408 3056 20460
rect 3108 20448 3114 20460
rect 3694 20448 3700 20460
rect 3108 20420 3700 20448
rect 3108 20408 3114 20420
rect 3694 20408 3700 20420
rect 3752 20448 3758 20460
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3752 20420 3801 20448
rect 3752 20408 3758 20420
rect 3789 20417 3801 20420
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 4982 20448 4988 20460
rect 4304 20420 4988 20448
rect 4304 20408 4310 20420
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 5074 20408 5080 20460
rect 5132 20448 5138 20460
rect 5350 20448 5356 20460
rect 5132 20420 5356 20448
rect 5132 20408 5138 20420
rect 5350 20408 5356 20420
rect 5408 20448 5414 20460
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 5408 20420 5549 20448
rect 5408 20408 5414 20420
rect 5537 20417 5549 20420
rect 5583 20417 5595 20451
rect 9950 20448 9956 20460
rect 9911 20420 9956 20448
rect 5537 20411 5595 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11256 20420 11805 20448
rect 1949 20383 2007 20389
rect 1949 20349 1961 20383
rect 1995 20380 2007 20383
rect 2130 20380 2136 20392
rect 1995 20352 2136 20380
rect 1995 20349 2007 20352
rect 1949 20343 2007 20349
rect 2130 20340 2136 20352
rect 2188 20340 2194 20392
rect 3145 20383 3203 20389
rect 3145 20349 3157 20383
rect 3191 20349 3203 20383
rect 3145 20343 3203 20349
rect 3160 20312 3188 20343
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3292 20352 3433 20380
rect 3292 20340 3298 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 4430 20380 4436 20392
rect 4111 20352 4436 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4430 20340 4436 20352
rect 4488 20340 4494 20392
rect 5994 20340 6000 20392
rect 6052 20380 6058 20392
rect 6546 20380 6552 20392
rect 6052 20352 6552 20380
rect 6052 20340 6058 20352
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6914 20380 6920 20392
rect 6871 20352 6920 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7650 20380 7656 20392
rect 7611 20352 7656 20380
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20380 7987 20383
rect 9306 20380 9312 20392
rect 7975 20352 9312 20380
rect 7975 20349 7987 20352
rect 7929 20343 7987 20349
rect 4706 20312 4712 20324
rect 3160 20284 4712 20312
rect 4706 20272 4712 20284
rect 4764 20272 4770 20324
rect 7944 20312 7972 20343
rect 9306 20340 9312 20352
rect 9364 20380 9370 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 9364 20352 9413 20380
rect 9364 20340 9370 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20380 9643 20383
rect 10318 20380 10324 20392
rect 9631 20352 10324 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11256 20380 11284 20420
rect 11793 20417 11805 20420
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 11514 20380 11520 20392
rect 11112 20352 11284 20380
rect 11475 20352 11520 20380
rect 11112 20340 11118 20352
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 11606 20340 11612 20392
rect 11664 20380 11670 20392
rect 11900 20380 11928 20488
rect 12636 20457 12664 20488
rect 15396 20488 19288 20516
rect 15396 20460 15424 20488
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 11664 20352 11928 20380
rect 11664 20340 11670 20352
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 13188 20380 13216 20411
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 13320 20420 14105 20448
rect 13320 20408 13326 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 14645 20451 14703 20457
rect 14645 20417 14657 20451
rect 14691 20417 14703 20451
rect 15194 20448 15200 20460
rect 15155 20420 15200 20448
rect 14645 20411 14703 20417
rect 12124 20352 13216 20380
rect 12124 20340 12130 20352
rect 13538 20340 13544 20392
rect 13596 20380 13602 20392
rect 14660 20380 14688 20411
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15746 20448 15752 20460
rect 15707 20420 15752 20448
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 17770 20448 17776 20460
rect 17731 20420 17776 20448
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20448 18383 20451
rect 18506 20448 18512 20460
rect 18371 20420 18512 20448
rect 18371 20417 18383 20420
rect 18325 20411 18383 20417
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 19260 20457 19288 20488
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 21094 20451 21152 20457
rect 21094 20448 21106 20451
rect 20128 20420 21106 20448
rect 20128 20408 20134 20420
rect 21094 20417 21106 20420
rect 21140 20417 21152 20451
rect 21094 20411 21152 20417
rect 13596 20352 14688 20380
rect 13596 20340 13602 20352
rect 16758 20340 16764 20392
rect 16816 20380 16822 20392
rect 20254 20380 20260 20392
rect 16816 20352 20260 20380
rect 16816 20340 16822 20352
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 4816 20284 7972 20312
rect 10137 20315 10195 20321
rect 3418 20204 3424 20256
rect 3476 20244 3482 20256
rect 4816 20244 4844 20284
rect 10137 20281 10149 20315
rect 10183 20312 10195 20315
rect 11882 20312 11888 20324
rect 10183 20284 11888 20312
rect 10183 20281 10195 20284
rect 10137 20275 10195 20281
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 12526 20312 12532 20324
rect 12406 20284 12532 20312
rect 3476 20216 4844 20244
rect 3476 20204 3482 20216
rect 4890 20204 4896 20256
rect 4948 20244 4954 20256
rect 5077 20247 5135 20253
rect 5077 20244 5089 20247
rect 4948 20216 5089 20244
rect 4948 20204 4954 20216
rect 5077 20213 5089 20216
rect 5123 20213 5135 20247
rect 5077 20207 5135 20213
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5629 20247 5687 20253
rect 5629 20244 5641 20247
rect 5592 20216 5641 20244
rect 5592 20204 5598 20216
rect 5629 20213 5641 20216
rect 5675 20213 5687 20247
rect 5629 20207 5687 20213
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8720 20216 8953 20244
rect 8720 20204 8726 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 10686 20204 10692 20256
rect 10744 20244 10750 20256
rect 12406 20244 12434 20284
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 14182 20272 14188 20324
rect 14240 20312 14246 20324
rect 14829 20315 14887 20321
rect 14829 20312 14841 20315
rect 14240 20284 14841 20312
rect 14240 20272 14246 20284
rect 14829 20281 14841 20284
rect 14875 20281 14887 20315
rect 14829 20275 14887 20281
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 15933 20315 15991 20321
rect 15933 20312 15945 20315
rect 15344 20284 15945 20312
rect 15344 20272 15350 20284
rect 15933 20281 15945 20284
rect 15979 20281 15991 20315
rect 15933 20275 15991 20281
rect 16390 20272 16396 20324
rect 16448 20312 16454 20324
rect 17405 20315 17463 20321
rect 17405 20312 17417 20315
rect 16448 20284 17417 20312
rect 16448 20272 16454 20284
rect 17405 20281 17417 20284
rect 17451 20281 17463 20315
rect 17405 20275 17463 20281
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 19150 20312 19156 20324
rect 18196 20284 19156 20312
rect 18196 20272 18202 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 10744 20216 12434 20244
rect 10744 20204 10750 20216
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17000 20216 17969 20244
rect 17000 20204 17006 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 17957 20207 18015 20213
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 18748 20216 19993 20244
rect 18748 20204 18754 20216
rect 19981 20213 19993 20216
rect 20027 20213 20039 20247
rect 19981 20207 20039 20213
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 21376 20244 21404 20343
rect 20772 20216 21404 20244
rect 20772 20204 20778 20216
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 3418 20040 3424 20052
rect 3379 20012 3424 20040
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 3878 20040 3884 20052
rect 3839 20012 3884 20040
rect 3878 20000 3884 20012
rect 3936 20000 3942 20052
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 10686 20040 10692 20052
rect 5307 20012 10692 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11606 20040 11612 20052
rect 10796 20012 11612 20040
rect 1765 19975 1823 19981
rect 1765 19941 1777 19975
rect 1811 19972 1823 19975
rect 3970 19972 3976 19984
rect 1811 19944 3976 19972
rect 1811 19941 1823 19944
rect 1765 19935 1823 19941
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 5718 19972 5724 19984
rect 5679 19944 5724 19972
rect 5718 19932 5724 19944
rect 5776 19932 5782 19984
rect 6546 19904 6552 19916
rect 4632 19876 6552 19904
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 1581 19839 1639 19845
rect 1581 19836 1593 19839
rect 1544 19808 1593 19836
rect 1544 19796 1550 19808
rect 1581 19805 1593 19808
rect 1627 19805 1639 19839
rect 1581 19799 1639 19805
rect 2038 19796 2044 19848
rect 2096 19836 2102 19848
rect 2225 19839 2283 19845
rect 2225 19836 2237 19839
rect 2096 19808 2237 19836
rect 2096 19796 2102 19808
rect 2225 19805 2237 19808
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 2685 19839 2743 19845
rect 2685 19836 2697 19839
rect 2648 19808 2697 19836
rect 2648 19796 2654 19808
rect 2685 19805 2697 19808
rect 2731 19805 2743 19839
rect 2685 19799 2743 19805
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4522 19836 4528 19848
rect 4203 19808 4528 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4632 19845 4660 19876
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7558 19904 7564 19916
rect 7340 19876 7564 19904
rect 7340 19864 7346 19876
rect 7558 19864 7564 19876
rect 7616 19904 7622 19916
rect 8110 19904 8116 19916
rect 7616 19876 8116 19904
rect 7616 19864 7622 19876
rect 8110 19864 8116 19876
rect 8168 19864 8174 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 9582 19904 9588 19916
rect 8444 19876 9588 19904
rect 8444 19864 8450 19876
rect 9582 19864 9588 19876
rect 9640 19864 9646 19916
rect 10796 19904 10824 20012
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12032 20012 12725 20040
rect 12032 20000 12038 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 12713 20003 12771 20009
rect 13633 20043 13691 20049
rect 13633 20009 13645 20043
rect 13679 20040 13691 20043
rect 17954 20040 17960 20052
rect 13679 20012 17960 20040
rect 13679 20009 13691 20012
rect 13633 20003 13691 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 18104 20012 18337 20040
rect 18104 20000 18110 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 18325 20003 18383 20009
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 14458 19972 14464 19984
rect 12216 19944 14464 19972
rect 12216 19932 12222 19944
rect 14458 19932 14464 19944
rect 14516 19932 14522 19984
rect 16025 19975 16083 19981
rect 16025 19941 16037 19975
rect 16071 19972 16083 19975
rect 17773 19975 17831 19981
rect 16071 19944 17724 19972
rect 16071 19941 16083 19944
rect 16025 19935 16083 19941
rect 10520 19876 10824 19904
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19836 5595 19839
rect 5626 19836 5632 19848
rect 5583 19808 5632 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 2409 19771 2467 19777
rect 2409 19737 2421 19771
rect 2455 19768 2467 19771
rect 2774 19768 2780 19780
rect 2455 19740 2780 19768
rect 2455 19737 2467 19740
rect 2409 19731 2467 19737
rect 2774 19728 2780 19740
rect 2832 19728 2838 19780
rect 4246 19768 4252 19780
rect 2884 19740 4252 19768
rect 2884 19709 2912 19740
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 5092 19768 5120 19799
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 5997 19839 6055 19845
rect 5997 19836 6009 19839
rect 5960 19808 6009 19836
rect 5960 19796 5966 19808
rect 5997 19805 6009 19808
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19836 6331 19839
rect 6638 19836 6644 19848
rect 6319 19808 6644 19836
rect 6319 19805 6331 19808
rect 6273 19799 6331 19805
rect 6638 19796 6644 19808
rect 6696 19796 6702 19848
rect 10520 19836 10548 19876
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 14366 19904 14372 19916
rect 11940 19876 14372 19904
rect 11940 19864 11946 19876
rect 14366 19864 14372 19876
rect 14424 19864 14430 19916
rect 17696 19904 17724 19944
rect 17773 19941 17785 19975
rect 17819 19972 17831 19975
rect 18138 19972 18144 19984
rect 17819 19944 18144 19972
rect 17819 19941 17831 19944
rect 17773 19935 17831 19941
rect 18138 19932 18144 19944
rect 18196 19932 18202 19984
rect 18046 19904 18052 19916
rect 16132 19876 17632 19904
rect 17696 19876 18052 19904
rect 7208 19808 10548 19836
rect 10597 19839 10655 19845
rect 6730 19768 6736 19780
rect 5092 19740 6736 19768
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19669 2927 19703
rect 4338 19700 4344 19712
rect 4299 19672 4344 19700
rect 2869 19663 2927 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 7208 19700 7236 19808
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10643 19808 10885 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10873 19805 10885 19808
rect 10919 19836 10931 19839
rect 10919 19808 12434 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 7340 19740 7385 19768
rect 7340 19728 7346 19740
rect 7466 19728 7472 19780
rect 7524 19768 7530 19780
rect 7837 19771 7895 19777
rect 7837 19768 7849 19771
rect 7524 19740 7849 19768
rect 7524 19728 7530 19740
rect 7837 19737 7849 19740
rect 7883 19768 7895 19771
rect 8202 19768 8208 19780
rect 7883 19740 8208 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 8202 19728 8208 19740
rect 8260 19728 8266 19780
rect 8386 19768 8392 19780
rect 8347 19740 8392 19768
rect 8386 19728 8392 19740
rect 8444 19728 8450 19780
rect 8573 19771 8631 19777
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 9398 19768 9404 19780
rect 8619 19740 9404 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 10318 19728 10324 19780
rect 10376 19777 10382 19780
rect 11146 19777 11152 19780
rect 10376 19768 10388 19777
rect 10376 19740 10421 19768
rect 10376 19731 10388 19740
rect 11140 19731 11152 19777
rect 11204 19768 11210 19780
rect 12406 19768 12434 19808
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 13446 19836 13452 19848
rect 12584 19808 12629 19836
rect 13407 19808 13452 19836
rect 12584 19796 12590 19808
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 15028 19832 15485 19836
rect 14936 19808 15485 19832
rect 14936 19804 15056 19808
rect 15473 19805 15485 19808
rect 15519 19836 15531 19839
rect 16022 19836 16028 19848
rect 15519 19808 16028 19836
rect 15519 19805 15531 19808
rect 13081 19771 13139 19777
rect 13081 19768 13093 19771
rect 11204 19740 11240 19768
rect 12406 19740 13093 19768
rect 10376 19728 10382 19731
rect 11146 19728 11152 19731
rect 11204 19728 11210 19740
rect 13081 19737 13093 19740
rect 13127 19768 13139 19771
rect 14936 19768 14964 19804
rect 15473 19799 15531 19805
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 13127 19740 14964 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 15206 19771 15264 19777
rect 15206 19768 15218 19771
rect 15160 19740 15218 19768
rect 15160 19728 15166 19740
rect 15206 19737 15218 19740
rect 15252 19737 15264 19771
rect 16132 19768 16160 19876
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 15206 19731 15264 19737
rect 15304 19740 16160 19768
rect 16224 19768 16252 19799
rect 16298 19796 16304 19848
rect 16356 19836 16362 19848
rect 17604 19845 17632 19876
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 16356 19808 16497 19836
rect 16356 19796 16362 19808
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 17589 19799 17647 19805
rect 17034 19768 17040 19780
rect 16224 19740 17040 19768
rect 7374 19700 7380 19712
rect 4847 19672 7236 19700
rect 7335 19672 7380 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 7926 19700 7932 19712
rect 7887 19672 7932 19700
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 8478 19660 8484 19712
rect 8536 19700 8542 19712
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 8536 19672 9229 19700
rect 8536 19660 8542 19672
rect 9217 19669 9229 19672
rect 9263 19700 9275 19703
rect 9490 19700 9496 19712
rect 9263 19672 9496 19700
rect 9263 19669 9275 19672
rect 9217 19663 9275 19669
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 9858 19660 9864 19712
rect 9916 19700 9922 19712
rect 10870 19700 10876 19712
rect 9916 19672 10876 19700
rect 9916 19660 9922 19672
rect 10870 19660 10876 19672
rect 10928 19700 10934 19712
rect 11514 19700 11520 19712
rect 10928 19672 11520 19700
rect 10928 19660 10934 19672
rect 11514 19660 11520 19672
rect 11572 19660 11578 19712
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 12618 19700 12624 19712
rect 12299 19672 12624 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 14093 19703 14151 19709
rect 14093 19669 14105 19703
rect 14139 19700 14151 19703
rect 14274 19700 14280 19712
rect 14139 19672 14280 19700
rect 14139 19669 14151 19672
rect 14093 19663 14151 19669
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 15304 19700 15332 19740
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 17328 19768 17356 19799
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18708 19836 18736 20003
rect 18874 19836 18880 19848
rect 18248 19808 18736 19836
rect 18835 19808 18880 19836
rect 18248 19768 18276 19808
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 20714 19836 20720 19848
rect 19567 19808 20720 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 21361 19839 21419 19845
rect 21361 19836 21373 19839
rect 20956 19808 21373 19836
rect 20956 19796 20962 19808
rect 21361 19805 21373 19808
rect 21407 19805 21419 19839
rect 21361 19799 21419 19805
rect 19794 19777 19800 19780
rect 19788 19768 19800 19777
rect 17328 19740 18276 19768
rect 18432 19740 18828 19768
rect 19755 19740 19800 19768
rect 14516 19672 15332 19700
rect 16669 19703 16727 19709
rect 14516 19660 14522 19672
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 16758 19700 16764 19712
rect 16715 19672 16764 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 16758 19660 16764 19672
rect 16816 19660 16822 19712
rect 17129 19703 17187 19709
rect 17129 19669 17141 19703
rect 17175 19700 17187 19703
rect 18432 19700 18460 19740
rect 17175 19672 18460 19700
rect 18800 19700 18828 19740
rect 19788 19731 19800 19740
rect 19794 19728 19800 19731
rect 19852 19728 19858 19780
rect 19978 19728 19984 19780
rect 20036 19768 20042 19780
rect 20036 19740 21220 19768
rect 20036 19728 20042 19740
rect 19702 19700 19708 19712
rect 18800 19672 19708 19700
rect 17175 19669 17187 19672
rect 17129 19663 17187 19669
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 20901 19703 20959 19709
rect 20901 19669 20913 19703
rect 20947 19700 20959 19703
rect 20990 19700 20996 19712
rect 20947 19672 20996 19700
rect 20947 19669 20959 19672
rect 20901 19663 20959 19669
rect 20990 19660 20996 19672
rect 21048 19660 21054 19712
rect 21192 19709 21220 19740
rect 21177 19703 21235 19709
rect 21177 19669 21189 19703
rect 21223 19669 21235 19703
rect 21177 19663 21235 19669
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 4062 19496 4068 19508
rect 1627 19468 4068 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 5721 19499 5779 19505
rect 5721 19496 5733 19499
rect 5031 19468 5733 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5721 19465 5733 19468
rect 5767 19465 5779 19499
rect 5721 19459 5779 19465
rect 5810 19456 5816 19508
rect 5868 19496 5874 19508
rect 6365 19499 6423 19505
rect 6365 19496 6377 19499
rect 5868 19468 6377 19496
rect 5868 19456 5874 19468
rect 6365 19465 6377 19468
rect 6411 19465 6423 19499
rect 6365 19459 6423 19465
rect 6638 19456 6644 19508
rect 6696 19496 6702 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6696 19468 6837 19496
rect 6696 19456 6702 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 7006 19496 7012 19508
rect 6825 19459 6883 19465
rect 6932 19468 7012 19496
rect 4154 19428 4160 19440
rect 4115 19400 4160 19428
rect 4154 19388 4160 19400
rect 4212 19388 4218 19440
rect 6932 19428 6960 19468
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7190 19456 7196 19508
rect 7248 19456 7254 19508
rect 8110 19496 8116 19508
rect 8023 19468 8116 19496
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 9306 19456 9312 19508
rect 9364 19496 9370 19508
rect 9490 19496 9496 19508
rect 9364 19468 9496 19496
rect 9364 19456 9370 19468
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 11149 19499 11207 19505
rect 11149 19465 11161 19499
rect 11195 19496 11207 19499
rect 11330 19496 11336 19508
rect 11195 19468 11336 19496
rect 11195 19465 11207 19468
rect 11149 19459 11207 19465
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 11701 19499 11759 19505
rect 11701 19465 11713 19499
rect 11747 19496 11759 19499
rect 11882 19496 11888 19508
rect 11747 19468 11888 19496
rect 11747 19465 11759 19468
rect 11701 19459 11759 19465
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12158 19496 12164 19508
rect 12119 19468 12164 19496
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12621 19499 12679 19505
rect 12621 19465 12633 19499
rect 12667 19496 12679 19499
rect 14550 19496 14556 19508
rect 12667 19468 14556 19496
rect 12667 19465 12679 19468
rect 12621 19459 12679 19465
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14642 19456 14648 19508
rect 14700 19496 14706 19508
rect 14700 19468 14745 19496
rect 14700 19456 14706 19468
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 16298 19496 16304 19508
rect 14884 19468 16304 19496
rect 14884 19456 14890 19468
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 18417 19499 18475 19505
rect 18417 19465 18429 19499
rect 18463 19465 18475 19499
rect 18417 19459 18475 19465
rect 18693 19499 18751 19505
rect 18693 19465 18705 19499
rect 18739 19496 18751 19499
rect 18782 19496 18788 19508
rect 18739 19468 18788 19496
rect 18739 19465 18751 19468
rect 18693 19459 18751 19465
rect 7098 19428 7104 19440
rect 6748 19400 6960 19428
rect 7024 19400 7104 19428
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 1320 19332 1409 19360
rect 934 19252 940 19304
rect 992 19292 998 19304
rect 1320 19292 1348 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 4798 19360 4804 19372
rect 4759 19332 4804 19360
rect 1397 19323 1455 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5592 19332 5641 19360
rect 5592 19320 5598 19332
rect 5629 19329 5641 19332
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5718 19320 5724 19372
rect 5776 19360 5782 19372
rect 6748 19369 6776 19400
rect 6733 19363 6791 19369
rect 5776 19332 5856 19360
rect 5776 19320 5782 19332
rect 2314 19292 2320 19304
rect 992 19264 1348 19292
rect 2275 19264 2320 19292
rect 992 19252 998 19264
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 5828 19301 5856 19332
rect 6733 19329 6745 19363
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 7024 19301 7052 19400
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 3789 19295 3847 19301
rect 2731 19264 3372 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 3053 19227 3111 19233
rect 3053 19193 3065 19227
rect 3099 19224 3111 19227
rect 3142 19224 3148 19236
rect 3099 19196 3148 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3344 19156 3372 19264
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 5813 19295 5871 19301
rect 3835 19264 5580 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 3421 19227 3479 19233
rect 3421 19193 3433 19227
rect 3467 19224 3479 19227
rect 4338 19224 4344 19236
rect 3467 19196 4344 19224
rect 3467 19193 3479 19196
rect 3421 19187 3479 19193
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 3878 19156 3884 19168
rect 3344 19128 3884 19156
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4212 19128 4445 19156
rect 4212 19116 4218 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5261 19159 5319 19165
rect 5261 19156 5273 19159
rect 5224 19128 5273 19156
rect 5224 19116 5230 19128
rect 5261 19125 5273 19128
rect 5307 19125 5319 19159
rect 5552 19156 5580 19264
rect 5813 19261 5825 19295
rect 5859 19261 5871 19295
rect 5813 19255 5871 19261
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19261 7067 19295
rect 7208 19292 7236 19456
rect 8128 19428 8156 19456
rect 10014 19431 10072 19437
rect 10014 19428 10026 19431
rect 8128 19400 10026 19428
rect 10014 19397 10026 19400
rect 10060 19397 10072 19431
rect 10014 19391 10072 19397
rect 10318 19388 10324 19440
rect 10376 19428 10382 19440
rect 12986 19428 12992 19440
rect 10376 19400 12992 19428
rect 10376 19388 10382 19400
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 15758 19431 15816 19437
rect 15758 19428 15770 19431
rect 13780 19400 15770 19428
rect 13780 19388 13786 19400
rect 15758 19397 15770 19400
rect 15804 19397 15816 19431
rect 18432 19428 18460 19459
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 20438 19496 20444 19508
rect 19628 19468 20444 19496
rect 19628 19428 19656 19468
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 18432 19400 19656 19428
rect 15758 19391 15816 19397
rect 19702 19388 19708 19440
rect 19760 19428 19766 19440
rect 19806 19431 19864 19437
rect 19806 19428 19818 19431
rect 19760 19400 19818 19428
rect 19760 19388 19766 19400
rect 19806 19397 19818 19400
rect 19852 19397 19864 19431
rect 19806 19391 19864 19397
rect 7653 19363 7711 19369
rect 7653 19329 7665 19363
rect 7699 19360 7711 19363
rect 7742 19360 7748 19372
rect 7699 19332 7748 19360
rect 7699 19329 7711 19332
rect 7653 19323 7711 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 9237 19363 9295 19369
rect 9237 19329 9249 19363
rect 9283 19360 9295 19363
rect 9582 19360 9588 19372
rect 9283 19332 9588 19360
rect 9283 19329 9295 19332
rect 9237 19323 9295 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 11514 19360 11520 19372
rect 11475 19332 11520 19360
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 11977 19323 12035 19329
rect 8386 19292 8392 19304
rect 7208 19264 8392 19292
rect 7009 19255 7067 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9769 19295 9827 19301
rect 9769 19292 9781 19295
rect 9539 19264 9781 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9769 19261 9781 19264
rect 9815 19261 9827 19295
rect 9769 19255 9827 19261
rect 7466 19156 7472 19168
rect 5552 19128 7472 19156
rect 5261 19119 5319 19125
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 7834 19156 7840 19168
rect 7795 19128 7840 19156
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 9508 19156 9536 19255
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11992 19292 12020 19323
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14102 19363 14160 19369
rect 14102 19360 14114 19363
rect 13872 19332 14114 19360
rect 13872 19320 13878 19332
rect 14102 19329 14114 19332
rect 14148 19329 14160 19363
rect 16022 19360 16028 19372
rect 15983 19332 16028 19360
rect 14102 19323 14160 19329
rect 16022 19320 16028 19332
rect 16080 19360 16086 19372
rect 16850 19360 16856 19372
rect 16080 19332 16856 19360
rect 16080 19320 16086 19332
rect 16850 19320 16856 19332
rect 16908 19360 16914 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16908 19332 17049 19360
rect 16908 19320 16914 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17304 19363 17362 19369
rect 17304 19329 17316 19363
rect 17350 19360 17362 19363
rect 20162 19360 20168 19372
rect 17350 19332 20168 19360
rect 17350 19329 17362 19332
rect 17304 19323 17362 19329
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 20346 19360 20352 19372
rect 20307 19332 20352 19360
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 14366 19292 14372 19304
rect 11020 19264 12020 19292
rect 14327 19264 14372 19292
rect 11020 19252 11026 19264
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19292 20131 19295
rect 20714 19292 20720 19304
rect 20119 19264 20720 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 13262 19224 13268 19236
rect 10836 19196 13268 19224
rect 10836 19184 10842 19196
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 16020 19196 16804 19224
rect 12986 19156 12992 19168
rect 8628 19128 9536 19156
rect 12947 19128 12992 19156
rect 8628 19116 8634 19128
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 16020 19156 16048 19196
rect 13780 19128 16048 19156
rect 13780 19116 13786 19128
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16632 19128 16681 19156
rect 16632 19116 16638 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16776 19156 16804 19196
rect 18230 19156 18236 19168
rect 16776 19128 18236 19156
rect 16669 19119 16727 19125
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 18598 19116 18604 19168
rect 18656 19156 18662 19168
rect 21542 19156 21548 19168
rect 18656 19128 21548 19156
rect 18656 19116 18662 19128
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 2038 18952 2044 18964
rect 1627 18924 2044 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4798 18952 4804 18964
rect 3467 18924 4804 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 8202 18952 8208 18964
rect 6503 18924 8208 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 9214 18912 9220 18964
rect 9272 18952 9278 18964
rect 9582 18952 9588 18964
rect 9272 18924 9588 18952
rect 9272 18912 9278 18924
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 11149 18955 11207 18961
rect 11149 18921 11161 18955
rect 11195 18952 11207 18955
rect 13446 18952 13452 18964
rect 11195 18924 13452 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 15194 18952 15200 18964
rect 13556 18924 15200 18952
rect 1949 18887 2007 18893
rect 1949 18853 1961 18887
rect 1995 18884 2007 18887
rect 2590 18884 2596 18896
rect 1995 18856 2596 18884
rect 1995 18853 2007 18856
rect 1949 18847 2007 18853
rect 2590 18844 2596 18856
rect 2648 18844 2654 18896
rect 3053 18887 3111 18893
rect 3053 18853 3065 18887
rect 3099 18884 3111 18887
rect 5074 18884 5080 18896
rect 3099 18856 5080 18884
rect 3099 18853 3111 18856
rect 3053 18847 3111 18853
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 6730 18884 6736 18896
rect 6691 18856 6736 18884
rect 6730 18844 6736 18856
rect 6788 18844 6794 18896
rect 6914 18844 6920 18896
rect 6972 18884 6978 18896
rect 7374 18884 7380 18896
rect 6972 18856 7380 18884
rect 6972 18844 6978 18856
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 8938 18884 8944 18896
rect 8899 18856 8944 18884
rect 8938 18844 8944 18856
rect 8996 18844 9002 18896
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 13556 18884 13584 18924
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 21358 18952 21364 18964
rect 18012 18924 21364 18952
rect 18012 18912 18018 18924
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 12860 18856 13584 18884
rect 12860 18844 12866 18856
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 4522 18816 4528 18828
rect 2363 18788 4528 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 4801 18819 4859 18825
rect 4801 18785 4813 18819
rect 4847 18816 4859 18819
rect 7282 18816 7288 18828
rect 4847 18788 7288 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 12728 18788 13032 18816
rect 4430 18748 4436 18760
rect 4391 18720 4436 18748
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18717 5871 18751
rect 5813 18711 5871 18717
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18748 6331 18751
rect 6638 18748 6644 18760
rect 6319 18720 6644 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 2685 18683 2743 18689
rect 2685 18649 2697 18683
rect 2731 18680 2743 18683
rect 3973 18683 4031 18689
rect 3973 18680 3985 18683
rect 2731 18652 3985 18680
rect 2731 18649 2743 18652
rect 2685 18643 2743 18649
rect 3973 18649 3985 18652
rect 4019 18680 4031 18683
rect 4154 18680 4160 18692
rect 4019 18652 4160 18680
rect 4019 18649 4031 18652
rect 3973 18643 4031 18649
rect 4154 18640 4160 18652
rect 4212 18680 4218 18692
rect 5077 18683 5135 18689
rect 5077 18680 5089 18683
rect 4212 18652 5089 18680
rect 4212 18640 4218 18652
rect 5077 18649 5089 18652
rect 5123 18680 5135 18683
rect 5258 18680 5264 18692
rect 5123 18652 5264 18680
rect 5123 18649 5135 18652
rect 5077 18643 5135 18649
rect 5258 18640 5264 18652
rect 5316 18680 5322 18692
rect 5445 18683 5503 18689
rect 5445 18680 5457 18683
rect 5316 18652 5457 18680
rect 5316 18640 5322 18652
rect 5445 18649 5457 18652
rect 5491 18649 5503 18683
rect 5828 18680 5856 18711
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 6914 18748 6920 18760
rect 6875 18720 6920 18748
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 8570 18748 8576 18760
rect 8531 18720 8576 18748
rect 8570 18708 8576 18720
rect 8628 18748 8634 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 8628 18720 10333 18748
rect 8628 18708 8634 18720
rect 10321 18717 10333 18720
rect 10367 18748 10379 18751
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10367 18720 10609 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10597 18717 10609 18720
rect 10643 18748 10655 18751
rect 10686 18748 10692 18760
rect 10643 18720 10692 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 12526 18748 12532 18760
rect 12584 18757 12590 18760
rect 11011 18720 12434 18748
rect 12496 18720 12532 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 7098 18680 7104 18692
rect 5828 18652 7104 18680
rect 5445 18643 5503 18649
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 8328 18683 8386 18689
rect 8328 18649 8340 18683
rect 8374 18680 8386 18683
rect 8938 18680 8944 18692
rect 8374 18652 8944 18680
rect 8374 18649 8386 18652
rect 8328 18643 8386 18649
rect 8938 18640 8944 18652
rect 8996 18640 9002 18692
rect 10054 18683 10112 18689
rect 10054 18680 10066 18683
rect 9048 18652 10066 18680
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 5626 18612 5632 18624
rect 3936 18584 5632 18612
rect 3936 18572 3942 18584
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 5997 18615 6055 18621
rect 5997 18581 6009 18615
rect 6043 18612 6055 18615
rect 6822 18612 6828 18624
rect 6043 18584 6828 18612
rect 6043 18581 6055 18584
rect 5997 18575 6055 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7193 18615 7251 18621
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 7282 18612 7288 18624
rect 7239 18584 7288 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 7650 18572 7656 18624
rect 7708 18612 7714 18624
rect 9048 18612 9076 18652
rect 10054 18649 10066 18652
rect 10100 18680 10112 18683
rect 12406 18680 12434 18720
rect 12526 18708 12532 18720
rect 12584 18711 12596 18757
rect 12584 18708 12590 18711
rect 12728 18680 12756 18788
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18717 12863 18751
rect 13004 18748 13032 18788
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 16850 18816 16856 18828
rect 13136 18788 14596 18816
rect 13136 18776 13142 18788
rect 13538 18748 13544 18760
rect 13004 18720 13544 18748
rect 12805 18711 12863 18717
rect 10100 18652 11468 18680
rect 12406 18652 12756 18680
rect 12820 18680 12848 18711
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13688 18720 13737 18748
rect 13688 18708 13694 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 14182 18748 14188 18760
rect 14095 18720 14188 18748
rect 13725 18711 13783 18717
rect 14182 18708 14188 18720
rect 14240 18748 14246 18760
rect 14366 18748 14372 18760
rect 14240 18720 14372 18748
rect 14240 18708 14246 18720
rect 14366 18708 14372 18720
rect 14424 18748 14430 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14424 18720 14473 18748
rect 14424 18708 14430 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14568 18748 14596 18788
rect 15488 18788 16528 18816
rect 16811 18788 16856 18816
rect 14717 18751 14775 18757
rect 14717 18748 14729 18751
rect 14568 18720 14729 18748
rect 14461 18711 14519 18717
rect 14717 18717 14729 18720
rect 14763 18717 14775 18751
rect 14717 18711 14775 18717
rect 12986 18680 12992 18692
rect 12820 18652 12992 18680
rect 10100 18649 10112 18652
rect 10054 18643 10112 18649
rect 11440 18621 11468 18652
rect 12986 18640 12992 18652
rect 13044 18640 13050 18692
rect 14476 18680 14504 18711
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15488 18748 15516 18788
rect 15160 18720 15516 18748
rect 15160 18708 15166 18720
rect 15746 18680 15752 18692
rect 14476 18652 15752 18680
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 16500 18680 16528 18788
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 20714 18816 20720 18828
rect 20671 18788 20720 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 20714 18776 20720 18788
rect 20772 18816 20778 18828
rect 21266 18816 21272 18828
rect 20772 18788 21272 18816
rect 20772 18776 20778 18788
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 18230 18748 18236 18760
rect 16623 18720 18236 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18690 18748 18696 18760
rect 18340 18720 18696 18748
rect 17120 18683 17178 18689
rect 17120 18680 17132 18683
rect 16500 18652 17132 18680
rect 17120 18649 17132 18652
rect 17166 18680 17178 18683
rect 18340 18680 18368 18720
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18748 18935 18751
rect 18923 18720 20852 18748
rect 18923 18717 18935 18720
rect 18877 18711 18935 18717
rect 19794 18680 19800 18692
rect 17166 18652 18368 18680
rect 18432 18652 19800 18680
rect 17166 18649 17178 18652
rect 17120 18643 17178 18649
rect 18432 18624 18460 18652
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 20438 18689 20444 18692
rect 20380 18683 20444 18689
rect 20380 18649 20392 18683
rect 20426 18649 20444 18683
rect 20380 18643 20444 18649
rect 20438 18640 20444 18643
rect 20496 18640 20502 18692
rect 20824 18680 20852 18720
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20956 18720 21097 18748
rect 20956 18708 20962 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 22554 18680 22560 18692
rect 20824 18652 22560 18680
rect 22554 18640 22560 18652
rect 22612 18640 22618 18692
rect 7708 18584 9076 18612
rect 11425 18615 11483 18621
rect 7708 18572 7714 18584
rect 11425 18581 11437 18615
rect 11471 18581 11483 18615
rect 11425 18575 11483 18581
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12308 18584 13093 18612
rect 12308 18572 12314 18584
rect 13081 18581 13093 18584
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 13541 18615 13599 18621
rect 13541 18581 13553 18615
rect 13587 18612 13599 18615
rect 13722 18612 13728 18624
rect 13587 18584 13728 18612
rect 13587 18581 13599 18584
rect 13541 18575 13599 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 15838 18612 15844 18624
rect 15799 18584 15844 18612
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16393 18615 16451 18621
rect 16393 18581 16405 18615
rect 16439 18612 16451 18615
rect 17954 18612 17960 18624
rect 16439 18584 17960 18612
rect 16439 18581 16451 18584
rect 16393 18575 16451 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 18414 18612 18420 18624
rect 18279 18584 18420 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18690 18612 18696 18624
rect 18651 18584 18696 18612
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18612 19303 18615
rect 19702 18612 19708 18624
rect 19291 18584 19708 18612
rect 19291 18581 19303 18584
rect 19245 18575 19303 18581
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 21269 18615 21327 18621
rect 21269 18581 21281 18615
rect 21315 18612 21327 18615
rect 21450 18612 21456 18624
rect 21315 18584 21456 18612
rect 21315 18581 21327 18584
rect 21269 18575 21327 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 934 18368 940 18420
rect 992 18408 998 18420
rect 1397 18411 1455 18417
rect 1397 18408 1409 18411
rect 992 18380 1409 18408
rect 992 18368 998 18380
rect 1397 18377 1409 18380
rect 1443 18377 1455 18411
rect 1397 18371 1455 18377
rect 1486 18368 1492 18420
rect 1544 18408 1550 18420
rect 1765 18411 1823 18417
rect 1765 18408 1777 18411
rect 1544 18380 1777 18408
rect 1544 18368 1550 18380
rect 1765 18377 1777 18380
rect 1811 18377 1823 18411
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 1765 18371 1823 18377
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 4154 18408 4160 18420
rect 3835 18380 4160 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 5258 18408 5264 18420
rect 5219 18380 5264 18408
rect 5258 18368 5264 18380
rect 5316 18408 5322 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5316 18380 5917 18408
rect 5316 18368 5322 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 5905 18371 5963 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7006 18408 7012 18420
rect 6967 18380 7012 18408
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8757 18411 8815 18417
rect 8757 18377 8769 18411
rect 8803 18408 8815 18411
rect 10778 18408 10784 18420
rect 8803 18380 10784 18408
rect 8803 18377 8815 18380
rect 8757 18371 8815 18377
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12434 18408 12440 18420
rect 12299 18380 12440 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12618 18368 12624 18420
rect 12676 18408 12682 18420
rect 13354 18408 13360 18420
rect 12676 18380 13360 18408
rect 12676 18368 12682 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 13538 18368 13544 18420
rect 13596 18408 13602 18420
rect 15562 18408 15568 18420
rect 13596 18380 15568 18408
rect 13596 18368 13602 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 15657 18411 15715 18417
rect 15657 18377 15669 18411
rect 15703 18408 15715 18411
rect 16850 18408 16856 18420
rect 15703 18380 16856 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 16942 18368 16948 18420
rect 17000 18368 17006 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 22186 18408 22192 18420
rect 17184 18380 22192 18408
rect 17184 18368 17190 18380
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 2685 18343 2743 18349
rect 2685 18309 2697 18343
rect 2731 18340 2743 18343
rect 3234 18340 3240 18352
rect 2731 18312 3240 18340
rect 2731 18309 2743 18312
rect 2685 18303 2743 18309
rect 3234 18300 3240 18312
rect 3292 18300 3298 18352
rect 3421 18343 3479 18349
rect 3421 18309 3433 18343
rect 3467 18340 3479 18343
rect 4982 18340 4988 18352
rect 3467 18312 4988 18340
rect 3467 18309 3479 18312
rect 3421 18303 3479 18309
rect 4982 18300 4988 18312
rect 5040 18300 5046 18352
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 5675 18312 7236 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 7208 18284 7236 18312
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 12710 18340 12716 18352
rect 9272 18312 11284 18340
rect 9272 18300 9278 18312
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 5902 18272 5908 18284
rect 4203 18244 5908 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 6730 18272 6736 18284
rect 6691 18244 6736 18272
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7190 18272 7196 18284
rect 7151 18244 7196 18272
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 7432 18244 7941 18272
rect 7432 18232 7438 18244
rect 7929 18241 7941 18244
rect 7975 18241 7987 18275
rect 7929 18235 7987 18241
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8076 18244 8585 18272
rect 8076 18232 8082 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 9766 18232 9772 18284
rect 9824 18272 9830 18284
rect 10146 18275 10204 18281
rect 10146 18272 10158 18275
rect 9824 18244 10158 18272
rect 9824 18232 9830 18244
rect 10146 18241 10158 18244
rect 10192 18241 10204 18275
rect 10146 18235 10204 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18272 10471 18275
rect 10686 18272 10692 18284
rect 10459 18244 10692 18272
rect 10459 18241 10471 18244
rect 10413 18235 10471 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 7558 18204 7564 18216
rect 4939 18176 7564 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 8113 18207 8171 18213
rect 8113 18173 8125 18207
rect 8159 18204 8171 18207
rect 8938 18204 8944 18216
rect 8159 18176 8944 18204
rect 8159 18173 8171 18176
rect 8113 18167 8171 18173
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 4525 18139 4583 18145
rect 4525 18105 4537 18139
rect 4571 18136 4583 18139
rect 5534 18136 5540 18148
rect 4571 18108 5540 18136
rect 4571 18105 4583 18108
rect 4525 18099 4583 18105
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 5718 18096 5724 18148
rect 5776 18136 5782 18148
rect 11146 18136 11152 18148
rect 5776 18108 9076 18136
rect 5776 18096 5782 18108
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 9048 18077 9076 18108
rect 10428 18108 11152 18136
rect 7469 18071 7527 18077
rect 7469 18068 7481 18071
rect 7064 18040 7481 18068
rect 7064 18028 7070 18040
rect 7469 18037 7481 18040
rect 7515 18037 7527 18071
rect 7469 18031 7527 18037
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 10428 18068 10456 18108
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 9079 18040 10456 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 10962 18068 10968 18080
rect 10652 18040 10968 18068
rect 10652 18028 10658 18040
rect 10962 18028 10968 18040
rect 11020 18068 11026 18080
rect 11057 18071 11115 18077
rect 11057 18068 11069 18071
rect 11020 18040 11069 18068
rect 11020 18028 11026 18040
rect 11057 18037 11069 18040
rect 11103 18037 11115 18071
rect 11256 18068 11284 18312
rect 11624 18312 12716 18340
rect 11624 18281 11652 18312
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 16960 18340 16988 18368
rect 17862 18340 17868 18352
rect 12912 18312 16068 18340
rect 11609 18275 11667 18281
rect 11609 18241 11621 18275
rect 11655 18241 11667 18275
rect 11609 18235 11667 18241
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12250 18272 12256 18284
rect 12115 18244 12256 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 11793 18139 11851 18145
rect 11793 18105 11805 18139
rect 11839 18136 11851 18139
rect 12912 18136 12940 18312
rect 13354 18232 13360 18284
rect 13412 18272 13418 18284
rect 13642 18275 13700 18281
rect 13642 18272 13654 18275
rect 13412 18244 13654 18272
rect 13412 18232 13418 18244
rect 13642 18241 13654 18244
rect 13688 18241 13700 18275
rect 13642 18235 13700 18241
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14182 18272 14188 18284
rect 13955 18244 14188 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14182 18232 14188 18244
rect 14240 18272 14246 18284
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14240 18244 14289 18272
rect 14240 18232 14246 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 16040 18281 16068 18312
rect 16684 18312 17868 18340
rect 16684 18281 16712 18312
rect 17862 18300 17868 18312
rect 17920 18340 17926 18352
rect 17920 18312 18368 18340
rect 17920 18300 17926 18312
rect 18340 18281 18368 18312
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 21116 18343 21174 18349
rect 21116 18340 21128 18343
rect 21048 18312 21128 18340
rect 21048 18300 21054 18312
rect 21116 18309 21128 18312
rect 21162 18340 21174 18343
rect 21542 18340 21548 18352
rect 21162 18312 21548 18340
rect 21162 18309 21174 18312
rect 21116 18303 21174 18309
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 14533 18275 14591 18281
rect 14533 18272 14545 18275
rect 14424 18244 14545 18272
rect 14424 18232 14430 18244
rect 14533 18241 14545 18244
rect 14579 18241 14591 18275
rect 14533 18235 14591 18241
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 16925 18275 16983 18281
rect 16925 18272 16937 18275
rect 16669 18235 16727 18241
rect 16776 18244 16937 18272
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16776 18204 16804 18244
rect 16925 18241 16937 18244
rect 16971 18241 16983 18275
rect 16925 18235 16983 18241
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 18581 18275 18639 18281
rect 18581 18241 18593 18275
rect 18627 18272 18639 18275
rect 18966 18272 18972 18284
rect 18627 18244 18972 18272
rect 18627 18241 18639 18244
rect 18581 18235 18639 18241
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 21266 18232 21272 18284
rect 21324 18272 21330 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 21324 18244 21373 18272
rect 21324 18232 21330 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 15896 18176 16804 18204
rect 15896 18164 15902 18176
rect 11839 18108 12940 18136
rect 11839 18105 11851 18108
rect 11793 18099 11851 18105
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 16298 18136 16304 18148
rect 15620 18108 16304 18136
rect 15620 18096 15626 18108
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 18322 18136 18328 18148
rect 17972 18108 18328 18136
rect 12529 18071 12587 18077
rect 12529 18068 12541 18071
rect 11256 18040 12541 18068
rect 11057 18031 11115 18037
rect 12529 18037 12541 18040
rect 12575 18037 12587 18071
rect 12529 18031 12587 18037
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 17972 18068 18000 18108
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 19705 18139 19763 18145
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 19751 18108 20484 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 16255 18040 18000 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 18104 18040 18149 18068
rect 18104 18028 18110 18040
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 18966 18068 18972 18080
rect 18748 18040 18972 18068
rect 18748 18028 18754 18040
rect 18966 18028 18972 18040
rect 19024 18068 19030 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19024 18040 19993 18068
rect 19024 18028 19030 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 20456 18068 20484 18108
rect 21082 18068 21088 18080
rect 20456 18040 21088 18068
rect 19981 18031 20039 18037
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 4154 17864 4160 17876
rect 4115 17836 4160 17864
rect 4154 17824 4160 17836
rect 4212 17864 4218 17876
rect 4433 17867 4491 17873
rect 4433 17864 4445 17867
rect 4212 17836 4445 17864
rect 4212 17824 4218 17836
rect 4433 17833 4445 17836
rect 4479 17864 4491 17867
rect 5350 17864 5356 17876
rect 4479 17836 5356 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 5350 17824 5356 17836
rect 5408 17864 5414 17876
rect 5537 17867 5595 17873
rect 5537 17864 5549 17867
rect 5408 17836 5549 17864
rect 5408 17824 5414 17836
rect 5537 17833 5549 17836
rect 5583 17864 5595 17867
rect 5905 17867 5963 17873
rect 5905 17864 5917 17867
rect 5583 17836 5917 17864
rect 5583 17833 5595 17836
rect 5537 17827 5595 17833
rect 5905 17833 5917 17836
rect 5951 17833 5963 17867
rect 5905 17827 5963 17833
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7098 17864 7104 17876
rect 7055 17836 7104 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 12158 17864 12164 17876
rect 7975 17836 12164 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13814 17864 13820 17876
rect 12492 17836 13820 17864
rect 12492 17824 12498 17836
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 14826 17864 14832 17876
rect 14200 17836 14688 17864
rect 14787 17836 14832 17864
rect 4893 17799 4951 17805
rect 4893 17765 4905 17799
rect 4939 17796 4951 17799
rect 5994 17796 6000 17808
rect 4939 17768 6000 17796
rect 4939 17765 4951 17768
rect 4893 17759 4951 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 6733 17799 6791 17805
rect 6733 17765 6745 17799
rect 6779 17796 6791 17799
rect 7834 17796 7840 17808
rect 6779 17768 7840 17796
rect 6779 17765 6791 17768
rect 6733 17759 6791 17765
rect 7834 17756 7840 17768
rect 7892 17796 7898 17808
rect 8018 17796 8024 17808
rect 7892 17768 8024 17796
rect 7892 17756 7898 17768
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 8389 17799 8447 17805
rect 8389 17765 8401 17799
rect 8435 17796 8447 17799
rect 9490 17796 9496 17808
rect 8435 17768 9496 17796
rect 8435 17765 8447 17768
rect 8389 17759 8447 17765
rect 9490 17756 9496 17768
rect 9548 17756 9554 17808
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11790 17796 11796 17808
rect 10928 17768 11796 17796
rect 10928 17756 10934 17768
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 13725 17799 13783 17805
rect 13725 17765 13737 17799
rect 13771 17796 13783 17799
rect 14200 17796 14228 17836
rect 13771 17768 14228 17796
rect 14277 17799 14335 17805
rect 13771 17765 13783 17768
rect 13725 17759 13783 17765
rect 14277 17765 14289 17799
rect 14323 17796 14335 17799
rect 14660 17796 14688 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 17218 17864 17224 17876
rect 15120 17836 17224 17864
rect 15120 17796 15148 17836
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 17402 17824 17408 17876
rect 17460 17864 17466 17876
rect 22462 17864 22468 17876
rect 17460 17836 22468 17864
rect 17460 17824 17466 17836
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 14323 17768 14596 17796
rect 14660 17768 15148 17796
rect 17129 17799 17187 17805
rect 14323 17765 14335 17768
rect 14277 17759 14335 17765
rect 2038 17728 2044 17740
rect 1999 17700 2044 17728
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 7374 17728 7380 17740
rect 6288 17700 7380 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 2056 17660 2084 17688
rect 1719 17632 2084 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 5169 17527 5227 17533
rect 5169 17524 5181 17527
rect 4212 17496 5181 17524
rect 4212 17484 4218 17496
rect 5169 17493 5181 17496
rect 5215 17524 5227 17527
rect 5442 17524 5448 17536
rect 5215 17496 5448 17524
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 6288 17533 6316 17700
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 14568 17728 14596 17768
rect 17129 17765 17141 17799
rect 17175 17765 17187 17799
rect 17129 17759 17187 17765
rect 15010 17728 15016 17740
rect 14568 17700 15016 17728
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 7190 17660 7196 17672
rect 7151 17632 7196 17660
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 7742 17660 7748 17672
rect 7703 17632 7748 17660
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8202 17660 8208 17672
rect 8163 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9364 17632 9781 17660
rect 9364 17620 9370 17632
rect 9769 17629 9781 17632
rect 9815 17660 9827 17663
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 9815 17632 11529 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 11517 17629 11529 17632
rect 11563 17660 11575 17663
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11563 17632 11805 17660
rect 11563 17629 11575 17632
rect 11517 17623 11575 17629
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 11940 17632 13553 17660
rect 11940 17620 11946 17632
rect 13541 17629 13553 17632
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14458 17660 14464 17672
rect 14139 17632 14464 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17660 14703 17663
rect 14734 17660 14740 17672
rect 14691 17632 14740 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15102 17660 15108 17672
rect 15063 17632 15108 17660
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 17144 17660 17172 17759
rect 15212 17632 17172 17660
rect 15212 17604 15240 17632
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 17920 17632 18521 17660
rect 17920 17620 17926 17632
rect 18509 17629 18521 17632
rect 18555 17660 18567 17663
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18555 17632 18797 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 18785 17629 18797 17632
rect 18831 17660 18843 17663
rect 18874 17660 18880 17672
rect 18831 17632 18880 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19659 17632 21036 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 21008 17604 21036 17632
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21324 17632 21373 17660
rect 21324 17620 21330 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 10014 17595 10072 17601
rect 10014 17592 10026 17595
rect 7340 17564 10026 17592
rect 7340 17552 7346 17564
rect 10014 17561 10026 17564
rect 10060 17561 10072 17595
rect 10014 17555 10072 17561
rect 10778 17552 10784 17604
rect 10836 17592 10842 17604
rect 12038 17595 12096 17601
rect 12038 17592 12050 17595
rect 10836 17564 12050 17592
rect 10836 17552 10842 17564
rect 12038 17561 12050 17564
rect 12084 17561 12096 17595
rect 12038 17555 12096 17561
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 15194 17592 15200 17604
rect 12216 17564 15200 17592
rect 12216 17552 12222 17564
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 15361 17595 15419 17601
rect 15361 17592 15373 17595
rect 15304 17564 15373 17592
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 5960 17496 6285 17524
rect 5960 17484 5966 17496
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6273 17487 6331 17493
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8628 17496 9045 17524
rect 8628 17484 8634 17496
rect 9033 17493 9045 17496
rect 9079 17524 9091 17527
rect 9306 17524 9312 17536
rect 9079 17496 9312 17524
rect 9079 17493 9091 17496
rect 9033 17487 9091 17493
rect 9306 17484 9312 17496
rect 9364 17524 9370 17536
rect 9401 17527 9459 17533
rect 9401 17524 9413 17527
rect 9364 17496 9413 17524
rect 9364 17484 9370 17496
rect 9401 17493 9413 17496
rect 9447 17493 9459 17527
rect 9401 17487 9459 17493
rect 9490 17484 9496 17536
rect 9548 17524 9554 17536
rect 10870 17524 10876 17536
rect 9548 17496 10876 17524
rect 9548 17484 9554 17496
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 11020 17496 11161 17524
rect 11020 17484 11026 17496
rect 11149 17493 11161 17496
rect 11195 17524 11207 17527
rect 12434 17524 12440 17536
rect 11195 17496 12440 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13173 17527 13231 17533
rect 13173 17524 13185 17527
rect 12584 17496 13185 17524
rect 12584 17484 12590 17496
rect 13173 17493 13185 17496
rect 13219 17524 13231 17527
rect 15304 17524 15332 17564
rect 15361 17561 15373 17564
rect 15407 17561 15419 17595
rect 15361 17555 15419 17561
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 16390 17592 16396 17604
rect 15620 17564 16396 17592
rect 15620 17552 15626 17564
rect 16390 17552 16396 17564
rect 16448 17552 16454 17604
rect 17126 17552 17132 17604
rect 17184 17592 17190 17604
rect 18046 17592 18052 17604
rect 17184 17564 18052 17592
rect 17184 17552 17190 17564
rect 18046 17552 18052 17564
rect 18104 17592 18110 17604
rect 18242 17595 18300 17601
rect 18242 17592 18254 17595
rect 18104 17564 18254 17592
rect 18104 17552 18110 17564
rect 18242 17561 18254 17564
rect 18288 17561 18300 17595
rect 18242 17555 18300 17561
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 21082 17552 21088 17604
rect 21140 17601 21146 17604
rect 21140 17595 21174 17601
rect 21162 17592 21174 17595
rect 22094 17592 22100 17604
rect 21162 17564 22100 17592
rect 21162 17561 21174 17564
rect 21140 17555 21174 17561
rect 21140 17552 21146 17555
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 13219 17496 15332 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 15470 17484 15476 17536
rect 15528 17524 15534 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 15528 17496 16497 17524
rect 15528 17484 15534 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16853 17527 16911 17533
rect 16853 17493 16865 17527
rect 16899 17524 16911 17527
rect 17218 17524 17224 17536
rect 16899 17496 17224 17524
rect 16899 17493 16911 17496
rect 16853 17487 16911 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17310 17484 17316 17536
rect 17368 17524 17374 17536
rect 18598 17524 18604 17536
rect 17368 17496 18604 17524
rect 17368 17484 17374 17496
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 19242 17484 19248 17536
rect 19300 17524 19306 17536
rect 19429 17527 19487 17533
rect 19429 17524 19441 17527
rect 19300 17496 19441 17524
rect 19300 17484 19306 17496
rect 19429 17493 19441 17496
rect 19475 17493 19487 17527
rect 19429 17487 19487 17493
rect 19518 17484 19524 17536
rect 19576 17524 19582 17536
rect 19981 17527 20039 17533
rect 19981 17524 19993 17527
rect 19576 17496 19993 17524
rect 19576 17484 19582 17496
rect 19981 17493 19993 17496
rect 20027 17493 20039 17527
rect 19981 17487 20039 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 5537 17323 5595 17329
rect 5537 17320 5549 17323
rect 4304 17292 5549 17320
rect 4304 17280 4310 17292
rect 5537 17289 5549 17292
rect 5583 17289 5595 17323
rect 5537 17283 5595 17289
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7742 17320 7748 17332
rect 6963 17292 7748 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 12158 17320 12164 17332
rect 8260 17292 12164 17320
rect 8260 17280 8266 17292
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13449 17323 13507 17329
rect 13449 17289 13461 17323
rect 13495 17320 13507 17323
rect 16209 17323 16267 17329
rect 13495 17292 16068 17320
rect 13495 17289 13507 17292
rect 13449 17283 13507 17289
rect 8570 17212 8576 17264
rect 8628 17252 8634 17264
rect 14734 17252 14740 17264
rect 8628 17224 10456 17252
rect 8628 17212 8634 17224
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4948 17156 4997 17184
rect 4948 17144 4954 17156
rect 4985 17153 4997 17156
rect 5031 17184 5043 17187
rect 5626 17184 5632 17196
rect 5031 17156 5632 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 9858 17184 9864 17196
rect 8067 17156 9864 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10134 17144 10140 17196
rect 10192 17193 10198 17196
rect 10428 17193 10456 17224
rect 12820 17224 14740 17252
rect 12820 17193 12848 17224
rect 14734 17212 14740 17224
rect 14792 17212 14798 17264
rect 15746 17252 15752 17264
rect 15120 17224 15752 17252
rect 15120 17196 15148 17224
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 10192 17184 10204 17193
rect 10413 17187 10471 17193
rect 10192 17156 10237 17184
rect 10192 17147 10204 17156
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10459 17156 10701 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 10689 17153 10701 17156
rect 10735 17184 10747 17187
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10735 17156 11069 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 11057 17153 11069 17156
rect 11103 17184 11115 17187
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11103 17156 11713 17184
rect 11103 17153 11115 17156
rect 11057 17147 11115 17153
rect 11701 17153 11713 17156
rect 11747 17184 11759 17187
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11747 17156 12081 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 12069 17153 12081 17156
rect 12115 17184 12127 17187
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12115 17156 12449 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17153 12863 17187
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 12805 17147 12863 17153
rect 10192 17144 10198 17147
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 14838 17188 14896 17193
rect 14838 17187 14964 17188
rect 14838 17153 14850 17187
rect 14884 17184 14964 17187
rect 14884 17160 15056 17184
rect 14884 17153 14896 17160
rect 14936 17156 15056 17160
rect 14838 17147 14896 17153
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5534 17116 5540 17128
rect 5491 17088 5540 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 9306 17116 9312 17128
rect 7699 17088 9312 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 15028 17116 15056 17156
rect 15102 17144 15108 17196
rect 15160 17184 15166 17196
rect 15562 17184 15568 17196
rect 15160 17156 15253 17184
rect 15523 17156 15568 17184
rect 15160 17144 15166 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 16040 17193 16068 17292
rect 16209 17289 16221 17323
rect 16255 17289 16267 17323
rect 16209 17283 16267 17289
rect 16853 17323 16911 17329
rect 16853 17289 16865 17323
rect 16899 17320 16911 17323
rect 17310 17320 17316 17332
rect 16899 17292 17316 17320
rect 16899 17289 16911 17292
rect 16853 17283 16911 17289
rect 16224 17252 16252 17283
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 17957 17323 18015 17329
rect 17957 17289 17969 17323
rect 18003 17289 18015 17323
rect 18414 17320 18420 17332
rect 18375 17292 18420 17320
rect 17957 17283 18015 17289
rect 17402 17252 17408 17264
rect 16224 17224 17408 17252
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 17972 17252 18000 17283
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 20806 17252 20812 17264
rect 17972 17224 20812 17252
rect 20806 17212 20812 17224
rect 20864 17212 20870 17264
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 16025 17147 16083 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17218 17184 17224 17196
rect 17179 17156 17224 17184
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17368 17156 17785 17184
rect 17368 17144 17374 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 18598 17184 18604 17196
rect 18559 17156 18604 17184
rect 17773 17147 17831 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 20001 17187 20059 17193
rect 20001 17153 20013 17187
rect 20047 17184 20059 17187
rect 20346 17184 20352 17196
rect 20047 17156 20352 17184
rect 20047 17153 20059 17156
rect 20001 17147 20059 17153
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17184 21143 17187
rect 21634 17184 21640 17196
rect 21131 17156 21640 17184
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 15286 17116 15292 17128
rect 15028 17088 15292 17116
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 18506 17116 18512 17128
rect 17052 17088 18512 17116
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 6457 17051 6515 17057
rect 6457 17048 6469 17051
rect 5408 17020 6469 17048
rect 5408 17008 5414 17020
rect 6457 17017 6469 17020
rect 6503 17048 6515 17051
rect 7193 17051 7251 17057
rect 7193 17048 7205 17051
rect 6503 17020 7205 17048
rect 6503 17017 6515 17020
rect 6457 17011 6515 17017
rect 7193 17017 7205 17020
rect 7239 17048 7251 17051
rect 8297 17051 8355 17057
rect 8297 17048 8309 17051
rect 7239 17020 8309 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 8297 17017 8309 17020
rect 8343 17048 8355 17051
rect 8570 17048 8576 17060
rect 8343 17020 8576 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 8570 17008 8576 17020
rect 8628 17048 8634 17060
rect 8665 17051 8723 17057
rect 8665 17048 8677 17051
rect 8628 17020 8677 17048
rect 8628 17008 8634 17020
rect 8665 17017 8677 17020
rect 8711 17017 8723 17051
rect 8665 17011 8723 17017
rect 12989 17051 13047 17057
rect 12989 17017 13001 17051
rect 13035 17048 13047 17051
rect 15749 17051 15807 17057
rect 13035 17020 14228 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 5994 16980 6000 16992
rect 5955 16952 6000 16980
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 9033 16983 9091 16989
rect 9033 16949 9045 16983
rect 9079 16980 9091 16983
rect 10226 16980 10232 16992
rect 9079 16952 10232 16980
rect 9079 16949 9091 16952
rect 9033 16943 9091 16949
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 12492 16952 13737 16980
rect 12492 16940 12498 16952
rect 13725 16949 13737 16952
rect 13771 16949 13783 16983
rect 14200 16980 14228 17020
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 17052 17048 17080 17088
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 20257 17119 20315 17125
rect 20257 17085 20269 17119
rect 20303 17116 20315 17119
rect 21266 17116 21272 17128
rect 20303 17088 21272 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 19058 17048 19064 17060
rect 15795 17020 17080 17048
rect 17328 17020 19064 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 17328 16980 17356 17020
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 14200 16952 17356 16980
rect 17405 16983 17463 16989
rect 13725 16943 13783 16949
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 17954 16980 17960 16992
rect 17451 16952 17960 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 18877 16983 18935 16989
rect 18877 16980 18889 16983
rect 18564 16952 18889 16980
rect 18564 16940 18570 16952
rect 18877 16949 18889 16952
rect 18923 16949 18935 16983
rect 18877 16943 18935 16949
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20680 16952 20729 16980
rect 20680 16940 20686 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 5350 16776 5356 16788
rect 5311 16748 5356 16776
rect 5350 16736 5356 16748
rect 5408 16776 5414 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5408 16748 6009 16776
rect 5408 16736 5414 16748
rect 5997 16745 6009 16748
rect 6043 16776 6055 16779
rect 6825 16779 6883 16785
rect 6825 16776 6837 16779
rect 6043 16748 6837 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6825 16745 6837 16748
rect 6871 16745 6883 16779
rect 6825 16739 6883 16745
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7248 16748 7665 16776
rect 7248 16736 7254 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 13538 16776 13544 16788
rect 7653 16739 7711 16745
rect 8128 16748 13544 16776
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 4948 16612 5641 16640
rect 4948 16600 4954 16612
rect 5629 16609 5641 16612
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 8128 16649 8156 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 13725 16779 13783 16785
rect 13725 16745 13737 16779
rect 13771 16776 13783 16779
rect 16666 16776 16672 16788
rect 13771 16748 16672 16776
rect 13771 16745 13783 16748
rect 13725 16739 13783 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 19518 16776 19524 16788
rect 16776 16748 19524 16776
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15473 16711 15531 16717
rect 15473 16708 15485 16711
rect 15344 16680 15485 16708
rect 15344 16668 15350 16680
rect 15473 16677 15485 16680
rect 15519 16677 15531 16711
rect 15473 16671 15531 16677
rect 7193 16643 7251 16649
rect 7193 16640 7205 16643
rect 6880 16612 7205 16640
rect 6880 16600 6886 16612
rect 7193 16609 7205 16612
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8260 16612 8305 16640
rect 8260 16600 8266 16612
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8628 16612 8953 16640
rect 8628 16600 8634 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 12342 16640 12348 16652
rect 8941 16603 8999 16609
rect 11992 16612 12348 16640
rect 8956 16572 8984 16603
rect 10686 16572 10692 16584
rect 8956 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 10956 16575 11014 16581
rect 10956 16541 10968 16575
rect 11002 16572 11014 16575
rect 11992 16572 12020 16612
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12483 16612 13277 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 13265 16609 13277 16612
rect 13311 16640 13323 16643
rect 13446 16640 13452 16652
rect 13311 16612 13452 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13446 16600 13452 16612
rect 13504 16640 13510 16652
rect 15746 16640 15752 16652
rect 13504 16612 14136 16640
rect 13504 16600 13510 16612
rect 13078 16572 13084 16584
rect 11002 16544 12020 16572
rect 12084 16544 13084 16572
rect 11002 16541 11014 16544
rect 10956 16535 11014 16541
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 5592 16476 8156 16504
rect 5592 16464 5598 16476
rect 8128 16448 8156 16476
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 9186 16507 9244 16513
rect 9186 16504 9198 16507
rect 8996 16476 9198 16504
rect 8996 16464 9002 16476
rect 9186 16473 9198 16476
rect 9232 16473 9244 16507
rect 9186 16467 9244 16473
rect 12084 16448 12112 16544
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 14108 16581 14136 16612
rect 15100 16612 15752 16640
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13280 16544 13553 16572
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4212 16408 4537 16436
rect 4212 16396 4218 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 5718 16396 5724 16448
rect 5776 16436 5782 16448
rect 6365 16439 6423 16445
rect 6365 16436 6377 16439
rect 5776 16408 6377 16436
rect 5776 16396 5782 16408
rect 6365 16405 6377 16408
rect 6411 16405 6423 16439
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 6365 16399 6423 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 8168 16408 10333 16436
rect 8168 16396 8174 16408
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 10321 16399 10379 16405
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12802 16436 12808 16448
rect 12763 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16436 12866 16448
rect 13280 16436 13308 16544
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 15100 16572 15128 16612
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 14139 16544 15128 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 16005 16575 16063 16581
rect 16005 16572 16017 16575
rect 15252 16544 16017 16572
rect 15252 16532 15258 16544
rect 16005 16541 16017 16544
rect 16051 16541 16063 16575
rect 16005 16535 16063 16541
rect 13354 16464 13360 16516
rect 13412 16504 13418 16516
rect 14338 16507 14396 16513
rect 14338 16504 14350 16507
rect 13412 16476 14350 16504
rect 13412 16464 13418 16476
rect 14338 16473 14350 16476
rect 14384 16473 14396 16507
rect 14338 16467 14396 16473
rect 16206 16464 16212 16516
rect 16264 16504 16270 16516
rect 16776 16504 16804 16748
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 17129 16711 17187 16717
rect 17129 16677 17141 16711
rect 17175 16677 17187 16711
rect 17129 16671 17187 16677
rect 17144 16572 17172 16671
rect 18874 16640 18880 16652
rect 18835 16612 18880 16640
rect 18874 16600 18880 16612
rect 18932 16640 18938 16652
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 18932 16612 19257 16640
rect 18932 16600 18938 16612
rect 19245 16609 19257 16612
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 17586 16572 17592 16584
rect 17144 16544 17592 16572
rect 17586 16532 17592 16544
rect 17644 16572 17650 16584
rect 19501 16575 19559 16581
rect 19501 16572 19513 16575
rect 17644 16544 19513 16572
rect 17644 16532 17650 16544
rect 19501 16541 19513 16544
rect 19547 16541 19559 16575
rect 19501 16535 19559 16541
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 16264 16476 16804 16504
rect 16264 16464 16270 16476
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 18610 16507 18668 16513
rect 18610 16504 18622 16507
rect 18564 16476 18622 16504
rect 18564 16464 18570 16476
rect 18610 16473 18622 16476
rect 18656 16473 18668 16507
rect 18610 16467 18668 16473
rect 12860 16408 13308 16436
rect 12860 16396 12866 16408
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 15988 16408 17509 16436
rect 15988 16396 15994 16408
rect 17497 16405 17509 16408
rect 17543 16436 17555 16439
rect 17678 16436 17684 16448
rect 17543 16408 17684 16436
rect 17543 16405 17555 16408
rect 17497 16399 17555 16405
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 20346 16396 20352 16448
rect 20404 16436 20410 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20404 16408 20637 16436
rect 20404 16396 20410 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16436 21327 16439
rect 21450 16436 21456 16448
rect 21315 16408 21456 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5810 16232 5816 16244
rect 5307 16204 5816 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 7006 16232 7012 16244
rect 6687 16204 7012 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 9122 16232 9128 16244
rect 7484 16204 9128 16232
rect 7484 16164 7512 16204
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 14921 16235 14979 16241
rect 14921 16201 14933 16235
rect 14967 16232 14979 16235
rect 15654 16232 15660 16244
rect 14967 16204 15660 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16201 16175 16235
rect 16117 16195 16175 16201
rect 8570 16164 8576 16176
rect 5736 16136 7512 16164
rect 7576 16136 8576 16164
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4948 16068 5181 16096
rect 4948 16056 4954 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 16028 4123 16031
rect 4614 16028 4620 16040
rect 4111 16000 4620 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 3988 15960 4016 15991
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 16028 5503 16031
rect 5736 16028 5764 16136
rect 5810 16056 5816 16108
rect 5868 16096 5874 16108
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 5868 16068 6745 16096
rect 5868 16056 5874 16068
rect 6733 16065 6745 16068
rect 6779 16096 6791 16099
rect 6822 16096 6828 16108
rect 6779 16068 6828 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7576 16105 7604 16136
rect 8570 16124 8576 16136
rect 8628 16124 8634 16176
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 10330 16167 10388 16173
rect 10330 16164 10342 16167
rect 10284 16136 10342 16164
rect 10284 16124 10290 16136
rect 10330 16133 10342 16136
rect 10376 16133 10388 16167
rect 10330 16127 10388 16133
rect 13630 16124 13636 16176
rect 13688 16164 13694 16176
rect 16132 16164 16160 16195
rect 16850 16192 16856 16244
rect 16908 16232 16914 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 16908 16204 18061 16232
rect 16908 16192 16914 16204
rect 18049 16201 18061 16204
rect 18095 16232 18107 16235
rect 18095 16204 18644 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 17862 16164 17868 16176
rect 13688 16136 16160 16164
rect 16684 16136 17868 16164
rect 13688 16124 13694 16136
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7817 16099 7875 16105
rect 7817 16096 7829 16099
rect 7561 16059 7619 16065
rect 7668 16068 7829 16096
rect 5491 16000 5764 16028
rect 6549 16031 6607 16037
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 6549 15997 6561 16031
rect 6595 16028 6607 16031
rect 7006 16028 7012 16040
rect 6595 16000 7012 16028
rect 6595 15997 6607 16000
rect 6549 15991 6607 15997
rect 5460 15960 5488 15991
rect 7006 15988 7012 16000
rect 7064 16028 7070 16040
rect 7282 16028 7288 16040
rect 7064 16000 7288 16028
rect 7064 15988 7070 16000
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 7668 16028 7696 16068
rect 7817 16065 7829 16068
rect 7863 16096 7875 16099
rect 10597 16099 10655 16105
rect 7863 16068 10548 16096
rect 7863 16065 7875 16068
rect 7817 16059 7875 16065
rect 7576 16000 7696 16028
rect 10520 16028 10548 16068
rect 10597 16065 10609 16099
rect 10643 16096 10655 16099
rect 10686 16096 10692 16108
rect 10643 16068 10692 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 12998 16099 13056 16105
rect 12998 16096 13010 16099
rect 12768 16068 13010 16096
rect 12768 16056 12774 16068
rect 12998 16065 13010 16068
rect 13044 16065 13056 16099
rect 12998 16059 13056 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13446 16096 13452 16108
rect 13311 16068 13452 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13446 16056 13452 16068
rect 13504 16096 13510 16108
rect 13814 16105 13820 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13504 16068 13553 16096
rect 13504 16056 13510 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13808 16096 13820 16105
rect 13775 16068 13820 16096
rect 13541 16059 13599 16065
rect 13808 16059 13820 16068
rect 13814 16056 13820 16059
rect 13872 16056 13878 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15841 16099 15899 16105
rect 15243 16068 15700 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 10520 16000 11928 16028
rect 3988 15932 5488 15960
rect 7190 15920 7196 15972
rect 7248 15960 7254 15972
rect 7576 15960 7604 16000
rect 11900 15969 11928 16000
rect 15672 15969 15700 16068
rect 15841 16065 15853 16099
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16482 16096 16488 16108
rect 16347 16068 16488 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 15856 16028 15884 16059
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 16684 16105 16712 16136
rect 17862 16124 17868 16136
rect 17920 16164 17926 16176
rect 18616 16164 18644 16204
rect 18754 16167 18812 16173
rect 18754 16164 18766 16167
rect 17920 16136 18552 16164
rect 18616 16136 18766 16164
rect 17920 16124 17926 16136
rect 16942 16105 16948 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16936 16096 16948 16105
rect 16903 16068 16948 16096
rect 16669 16059 16727 16065
rect 16936 16059 16948 16068
rect 16574 16028 16580 16040
rect 15856 16000 16580 16028
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 7248 15932 7604 15960
rect 11885 15963 11943 15969
rect 7248 15920 7254 15932
rect 11885 15929 11897 15963
rect 11931 15929 11943 15963
rect 11885 15923 11943 15929
rect 15381 15963 15439 15969
rect 15381 15929 15393 15963
rect 15427 15960 15439 15963
rect 15657 15963 15715 15969
rect 15427 15932 15608 15960
rect 15427 15929 15439 15932
rect 15381 15923 15439 15929
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5997 15895 6055 15901
rect 5997 15861 6009 15895
rect 6043 15892 6055 15895
rect 6362 15892 6368 15904
rect 6043 15864 6368 15892
rect 6043 15861 6055 15864
rect 5997 15855 6055 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7926 15892 7932 15904
rect 7147 15864 7932 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8938 15892 8944 15904
rect 8352 15864 8944 15892
rect 8352 15852 8358 15864
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 9950 15892 9956 15904
rect 9263 15864 9956 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10744 15864 10977 15892
rect 10744 15852 10750 15864
rect 10965 15861 10977 15864
rect 11011 15892 11023 15895
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11011 15864 11621 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11609 15861 11621 15864
rect 11655 15892 11667 15895
rect 11698 15892 11704 15904
rect 11655 15864 11704 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12618 15892 12624 15904
rect 12032 15864 12624 15892
rect 12032 15852 12038 15864
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 15580 15892 15608 15932
rect 15657 15929 15669 15963
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 15746 15920 15752 15972
rect 15804 15960 15810 15972
rect 16684 15960 16712 16059
rect 16942 16056 16948 16059
rect 17000 16056 17006 16108
rect 18524 16105 18552 16136
rect 18754 16133 18766 16136
rect 18800 16133 18812 16167
rect 20070 16164 20076 16176
rect 18754 16127 18812 16133
rect 18892 16136 20076 16164
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16065 18567 16099
rect 18892 16096 18920 16136
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 18509 16059 18567 16065
rect 18616 16068 18920 16096
rect 17678 15988 17684 16040
rect 17736 16028 17742 16040
rect 18616 16028 18644 16068
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 19944 16068 20545 16096
rect 19944 16056 19950 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16096 21143 16099
rect 21174 16096 21180 16108
rect 21131 16068 21180 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 17736 16000 18644 16028
rect 17736 15988 17742 16000
rect 15804 15932 16712 15960
rect 15804 15920 15810 15932
rect 19518 15920 19524 15972
rect 19576 15960 19582 15972
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 19576 15932 20177 15960
rect 19576 15920 19582 15932
rect 20165 15929 20177 15932
rect 20211 15929 20223 15963
rect 20165 15923 20223 15929
rect 17310 15892 17316 15904
rect 15580 15864 17316 15892
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 19794 15852 19800 15904
rect 19852 15892 19858 15904
rect 19889 15895 19947 15901
rect 19889 15892 19901 15895
rect 19852 15864 19901 15892
rect 19852 15852 19858 15864
rect 19889 15861 19901 15864
rect 19935 15861 19947 15895
rect 20714 15892 20720 15904
rect 20675 15864 20720 15892
rect 19889 15855 19947 15861
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 7006 15688 7012 15700
rect 5276 15660 7012 15688
rect 5276 15561 5304 15660
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 8570 15688 8576 15700
rect 7208 15660 8576 15688
rect 5813 15623 5871 15629
rect 5813 15589 5825 15623
rect 5859 15620 5871 15623
rect 7098 15620 7104 15632
rect 5859 15592 7104 15620
rect 5859 15589 5871 15592
rect 5813 15583 5871 15589
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 7208 15561 7236 15660
rect 8570 15648 8576 15660
rect 8628 15688 8634 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8628 15660 8953 15688
rect 8628 15648 8634 15660
rect 8941 15657 8953 15660
rect 8987 15688 8999 15691
rect 9030 15688 9036 15700
rect 8987 15660 9036 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9030 15648 9036 15660
rect 9088 15688 9094 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 9088 15660 9321 15688
rect 9088 15648 9094 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10100 15660 11192 15688
rect 10100 15648 10106 15660
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 9766 15620 9772 15632
rect 8260 15592 9772 15620
rect 8260 15580 8266 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 11164 15620 11192 15660
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 14366 15688 14372 15700
rect 13596 15660 14372 15688
rect 13596 15648 13602 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 17681 15691 17739 15697
rect 16540 15660 16804 15688
rect 16540 15648 16546 15660
rect 12069 15623 12127 15629
rect 12069 15620 12081 15623
rect 11164 15592 12081 15620
rect 12069 15589 12081 15592
rect 12115 15589 12127 15623
rect 16776 15620 16804 15660
rect 17681 15657 17693 15691
rect 17727 15688 17739 15691
rect 17770 15688 17776 15700
rect 17727 15660 17776 15688
rect 17727 15657 17739 15660
rect 17681 15651 17739 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 18230 15688 18236 15700
rect 18191 15660 18236 15688
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18656 15660 18705 15688
rect 18656 15648 18662 15660
rect 18693 15657 18705 15660
rect 18739 15657 18751 15691
rect 19610 15688 19616 15700
rect 19571 15660 19616 15688
rect 18693 15651 18751 15657
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 19978 15620 19984 15632
rect 16776 15592 19984 15620
rect 12069 15583 12127 15589
rect 19978 15580 19984 15592
rect 20036 15580 20042 15632
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15521 7251 15555
rect 7193 15515 7251 15521
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15552 11207 15555
rect 11698 15552 11704 15564
rect 11195 15524 11704 15552
rect 11195 15521 11207 15524
rect 11149 15515 11207 15521
rect 5445 15487 5503 15493
rect 5445 15453 5457 15487
rect 5491 15484 5503 15487
rect 5718 15484 5724 15496
rect 5491 15456 5724 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 6546 15484 6552 15496
rect 6503 15456 6552 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 6748 15484 6776 15515
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 13446 15552 13452 15564
rect 13407 15524 13452 15552
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 15746 15552 15752 15564
rect 15611 15524 15752 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 15746 15512 15752 15524
rect 15804 15552 15810 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 15804 15524 15853 15552
rect 15804 15512 15810 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 11974 15484 11980 15496
rect 6748 15456 11980 15484
rect 5074 15376 5080 15428
rect 5132 15416 5138 15428
rect 6748 15416 6776 15456
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 13280 15456 17509 15484
rect 5132 15388 6776 15416
rect 5132 15376 5138 15388
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 7460 15419 7518 15425
rect 7460 15416 7472 15419
rect 6880 15388 7472 15416
rect 6880 15376 6886 15388
rect 7460 15385 7472 15388
rect 7506 15416 7518 15419
rect 8110 15416 8116 15428
rect 7506 15388 8116 15416
rect 7506 15385 7518 15388
rect 7460 15379 7518 15385
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 9214 15416 9220 15428
rect 8588 15388 9220 15416
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15348 5411 15351
rect 5442 15348 5448 15360
rect 5399 15320 5448 15348
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5592 15320 6101 15348
rect 5592 15308 5598 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 8588 15357 8616 15388
rect 9214 15376 9220 15388
rect 9272 15416 9278 15428
rect 10882 15419 10940 15425
rect 10882 15416 10894 15419
rect 9272 15388 10894 15416
rect 9272 15376 9278 15388
rect 10882 15385 10894 15388
rect 10928 15385 10940 15419
rect 10882 15379 10940 15385
rect 11517 15419 11575 15425
rect 11517 15385 11529 15419
rect 11563 15416 11575 15419
rect 11698 15416 11704 15428
rect 11563 15388 11704 15416
rect 11563 15385 11575 15388
rect 11517 15379 11575 15385
rect 11698 15376 11704 15388
rect 11756 15376 11762 15428
rect 13182 15419 13240 15425
rect 13182 15416 13194 15419
rect 12406 15388 13194 15416
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 6420 15320 6561 15348
rect 6420 15308 6426 15320
rect 6549 15317 6561 15320
rect 6595 15317 6607 15351
rect 6549 15311 6607 15317
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15317 8631 15351
rect 8573 15311 8631 15317
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 12406 15348 12434 15388
rect 13182 15385 13194 15388
rect 13228 15385 13240 15419
rect 13182 15379 13240 15385
rect 13280 15360 13308 15456
rect 17497 15453 17509 15456
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 18598 15484 18604 15496
rect 18463 15456 18604 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 18874 15484 18880 15496
rect 18835 15456 18880 15484
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 19058 15444 19064 15496
rect 19116 15484 19122 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19116 15456 19441 15484
rect 19116 15444 19122 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 21324 15456 21373 15484
rect 21324 15444 21330 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 15298 15419 15356 15425
rect 15298 15416 15310 15419
rect 14976 15388 15310 15416
rect 14976 15376 14982 15388
rect 15298 15385 15310 15388
rect 15344 15385 15356 15419
rect 15298 15379 15356 15385
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 16086 15419 16144 15425
rect 16086 15416 16098 15419
rect 15712 15388 16098 15416
rect 15712 15376 15718 15388
rect 16086 15385 16098 15388
rect 16132 15385 16144 15419
rect 16086 15379 16144 15385
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 17770 15416 17776 15428
rect 16632 15388 17776 15416
rect 16632 15376 16638 15388
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 19904 15388 21036 15416
rect 10468 15320 12434 15348
rect 10468 15308 10474 15320
rect 13262 15308 13268 15360
rect 13320 15308 13326 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14182 15348 14188 15360
rect 13872 15320 14188 15348
rect 13872 15308 13878 15320
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 16390 15348 16396 15360
rect 14792 15320 16396 15348
rect 14792 15308 14798 15320
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 19904 15348 19932 15388
rect 17267 15320 19932 15348
rect 19981 15351 20039 15357
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 19981 15317 19993 15351
rect 20027 15348 20039 15351
rect 20162 15348 20168 15360
rect 20027 15320 20168 15348
rect 20027 15317 20039 15320
rect 19981 15311 20039 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 21008 15348 21036 15388
rect 21082 15376 21088 15428
rect 21140 15425 21146 15428
rect 21140 15416 21152 15425
rect 21140 15388 21185 15416
rect 21140 15379 21152 15388
rect 21140 15376 21146 15379
rect 22370 15348 22376 15360
rect 21008 15320 22376 15348
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 4856 15116 4905 15144
rect 4856 15104 4862 15116
rect 4893 15113 4905 15116
rect 4939 15113 4951 15147
rect 6546 15144 6552 15156
rect 6507 15116 6552 15144
rect 4893 15107 4951 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6696 15116 6837 15144
rect 6696 15104 6702 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7156 15116 8217 15144
rect 7156 15104 7162 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 9030 15144 9036 15156
rect 8991 15116 9036 15144
rect 8205 15107 8263 15113
rect 9030 15104 9036 15116
rect 9088 15144 9094 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9088 15116 9321 15144
rect 9088 15104 9094 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 4522 15036 4528 15088
rect 4580 15076 4586 15088
rect 4985 15079 5043 15085
rect 4985 15076 4997 15079
rect 4580 15048 4997 15076
rect 4580 15036 4586 15048
rect 4985 15045 4997 15048
rect 5031 15045 5043 15079
rect 4985 15039 5043 15045
rect 7285 15079 7343 15085
rect 7285 15045 7297 15079
rect 7331 15076 7343 15079
rect 7331 15048 7880 15076
rect 7331 15045 7343 15048
rect 7285 15039 7343 15045
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7558 15008 7564 15020
rect 7239 14980 7564 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7852 15008 7880 15048
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 8113 15079 8171 15085
rect 8113 15076 8125 15079
rect 7984 15048 8125 15076
rect 7984 15036 7990 15048
rect 8113 15045 8125 15048
rect 8159 15045 8171 15079
rect 8113 15039 8171 15045
rect 9324 15008 9352 15107
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 9640 15116 11069 15144
rect 9640 15104 9646 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11057 15107 11115 15113
rect 11609 15147 11667 15153
rect 11609 15113 11621 15147
rect 11655 15144 11667 15147
rect 11698 15144 11704 15156
rect 11655 15116 11704 15144
rect 11655 15113 11667 15116
rect 11609 15107 11667 15113
rect 10962 15076 10968 15088
rect 9784 15048 10968 15076
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 7852 14980 9260 15008
rect 9324 14980 9689 15008
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 7374 14940 7380 14952
rect 4847 14912 7380 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 9232 14940 9260 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9490 14940 9496 14952
rect 8067 14912 9168 14940
rect 9232 14912 9496 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5905 14807 5963 14813
rect 5905 14804 5917 14807
rect 5500 14776 5917 14804
rect 5500 14764 5506 14776
rect 5905 14773 5917 14776
rect 5951 14773 5963 14807
rect 7484 14804 7512 14903
rect 8570 14872 8576 14884
rect 8531 14844 8576 14872
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 9140 14872 9168 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9784 14940 9812 15048
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11072 15076 11100 15107
rect 11698 15104 11704 15116
rect 11756 15144 11762 15156
rect 11974 15144 11980 15156
rect 11756 15116 11980 15144
rect 11756 15104 11762 15116
rect 11974 15104 11980 15116
rect 12032 15144 12038 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 12032 15116 12081 15144
rect 12032 15104 12038 15116
rect 12069 15113 12081 15116
rect 12115 15144 12127 15147
rect 12437 15147 12495 15153
rect 12437 15144 12449 15147
rect 12115 15116 12449 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12437 15113 12449 15116
rect 12483 15113 12495 15147
rect 12437 15107 12495 15113
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 14918 15144 14924 15156
rect 14792 15116 14924 15144
rect 14792 15104 14798 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 16448 15116 16865 15144
rect 16448 15104 16454 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 16853 15107 16911 15113
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 17276 15116 17325 15144
rect 17276 15104 17282 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 18138 15144 18144 15156
rect 18003 15116 18144 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 18230 15104 18236 15156
rect 18288 15144 18294 15156
rect 18693 15147 18751 15153
rect 18693 15144 18705 15147
rect 18288 15116 18705 15144
rect 18288 15104 18294 15116
rect 18693 15113 18705 15116
rect 18739 15113 18751 15147
rect 18693 15107 18751 15113
rect 19978 15104 19984 15156
rect 20036 15104 20042 15156
rect 12158 15076 12164 15088
rect 11072 15048 12164 15076
rect 12158 15036 12164 15048
rect 12216 15036 12222 15088
rect 13265 15079 13323 15085
rect 13265 15045 13277 15079
rect 13311 15076 13323 15079
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 13311 15048 13645 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 13633 15045 13645 15048
rect 13679 15076 13691 15079
rect 13722 15076 13728 15088
rect 13679 15048 13728 15076
rect 13679 15045 13691 15048
rect 13633 15039 13691 15045
rect 13722 15036 13728 15048
rect 13780 15076 13786 15088
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 13780 15048 14289 15076
rect 13780 15036 13786 15048
rect 14277 15045 14289 15048
rect 14323 15076 14335 15079
rect 14645 15079 14703 15085
rect 14645 15076 14657 15079
rect 14323 15048 14657 15076
rect 14323 15045 14335 15048
rect 14277 15039 14335 15045
rect 14645 15045 14657 15048
rect 14691 15076 14703 15079
rect 15746 15076 15752 15088
rect 14691 15048 15752 15076
rect 14691 15045 14703 15048
rect 14645 15039 14703 15045
rect 15746 15036 15752 15048
rect 15804 15076 15810 15088
rect 16114 15076 16120 15088
rect 15804 15048 16120 15076
rect 15804 15036 15810 15048
rect 16114 15036 16120 15048
rect 16172 15076 16178 15088
rect 18322 15076 18328 15088
rect 16172 15048 16344 15076
rect 16172 15036 16178 15048
rect 9950 15017 9956 15020
rect 9933 15011 9956 15017
rect 9933 14977 9945 15011
rect 9933 14971 9956 14977
rect 9950 14968 9956 14971
rect 10008 14968 10014 15020
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 13354 15008 13360 15020
rect 10376 14980 13360 15008
rect 10376 14968 10382 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 16316 15017 16344 15048
rect 17512 15048 18328 15076
rect 16034 15011 16092 15017
rect 16034 15008 16046 15011
rect 13596 14980 16046 15008
rect 13596 14968 13602 14980
rect 16034 14977 16046 14980
rect 16080 14977 16092 15011
rect 16034 14971 16092 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16390 14968 16396 15020
rect 16448 15008 16454 15020
rect 17512 15017 17540 15048
rect 18322 15036 18328 15048
rect 18380 15076 18386 15088
rect 19518 15076 19524 15088
rect 18380 15048 19524 15076
rect 18380 15036 18386 15048
rect 19518 15036 19524 15048
rect 19576 15036 19582 15088
rect 19996 15076 20024 15104
rect 19720 15048 20024 15076
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16448 14980 17049 15008
rect 16448 14968 16454 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17678 14968 17684 15020
rect 17736 15008 17742 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17736 14980 17785 15008
rect 17736 14968 17742 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18196 14980 18429 15008
rect 18196 14968 18202 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 9646 14912 9812 14940
rect 9646 14872 9674 14912
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 14734 14940 14740 14952
rect 11940 14912 14740 14940
rect 11940 14900 11946 14912
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 18892 14940 18920 14971
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19720 15017 19748 15048
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 19116 14980 19165 15008
rect 19116 14968 19122 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 19961 15011 20019 15017
rect 19961 15008 19973 15011
rect 19852 14980 19973 15008
rect 19852 14968 19858 14980
rect 19961 14977 19973 14980
rect 20007 14977 20019 15011
rect 19961 14971 20019 14977
rect 19812 14940 19840 14968
rect 16316 14912 18920 14940
rect 19720 14912 19840 14940
rect 12066 14872 12072 14884
rect 9140 14844 9674 14872
rect 10980 14844 12072 14872
rect 10980 14804 11008 14844
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 12710 14872 12716 14884
rect 12216 14844 12716 14872
rect 12216 14832 12222 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 13872 14844 14596 14872
rect 13872 14832 13878 14844
rect 7484 14776 11008 14804
rect 5905 14767 5963 14773
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 12805 14807 12863 14813
rect 12805 14804 12817 14807
rect 11756 14776 12817 14804
rect 11756 14764 11762 14776
rect 12805 14773 12817 14776
rect 12851 14804 12863 14807
rect 14458 14804 14464 14816
rect 12851 14776 14464 14804
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14568 14804 14596 14844
rect 16316 14804 16344 14912
rect 17034 14832 17040 14884
rect 17092 14872 17098 14884
rect 18233 14875 18291 14881
rect 18233 14872 18245 14875
rect 17092 14844 18245 14872
rect 17092 14832 17098 14844
rect 18233 14841 18245 14844
rect 18279 14841 18291 14875
rect 19720 14872 19748 14912
rect 18233 14835 18291 14841
rect 18616 14844 19748 14872
rect 14568 14776 16344 14804
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 18616 14804 18644 14844
rect 17276 14776 18644 14804
rect 19337 14807 19395 14813
rect 17276 14764 17282 14776
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19518 14804 19524 14816
rect 19383 14776 19524 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 21082 14804 21088 14816
rect 20995 14776 21088 14804
rect 21082 14764 21088 14776
rect 21140 14804 21146 14816
rect 22462 14804 22468 14816
rect 21140 14776 22468 14804
rect 21140 14764 21146 14776
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 6914 14600 6920 14612
rect 6875 14572 6920 14600
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 8628 14572 9229 14600
rect 8628 14560 8634 14572
rect 9217 14569 9229 14572
rect 9263 14600 9275 14603
rect 10318 14600 10324 14612
rect 9263 14572 10324 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10965 14603 11023 14609
rect 10965 14569 10977 14603
rect 11011 14600 11023 14603
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11011 14572 11529 14600
rect 11011 14569 11023 14572
rect 10965 14563 11023 14569
rect 11517 14569 11529 14572
rect 11563 14600 11575 14603
rect 11885 14603 11943 14609
rect 11885 14600 11897 14603
rect 11563 14572 11897 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11885 14569 11897 14572
rect 11931 14600 11943 14603
rect 11974 14600 11980 14612
rect 11931 14572 11980 14600
rect 11931 14569 11943 14572
rect 11885 14563 11943 14569
rect 9582 14532 9588 14544
rect 4908 14504 9588 14532
rect 4908 14476 4936 14504
rect 9582 14492 9588 14504
rect 9640 14492 9646 14544
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4890 14464 4896 14476
rect 4203 14436 4896 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14464 5227 14467
rect 5258 14464 5264 14476
rect 5215 14436 5264 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 7469 14467 7527 14473
rect 7469 14464 7481 14467
rect 7300 14436 7481 14464
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4028 14368 4261 14396
rect 4028 14356 4034 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4396 14368 4441 14396
rect 4396 14356 4402 14368
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 5353 14399 5411 14405
rect 5353 14396 5365 14399
rect 4764 14368 5365 14396
rect 4764 14356 4770 14368
rect 5353 14365 5365 14368
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4120 14300 5273 14328
rect 4120 14288 4126 14300
rect 5261 14297 5273 14300
rect 5307 14297 5319 14331
rect 7300 14328 7328 14436
rect 7469 14433 7481 14436
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10980 14464 11008 14563
rect 11974 14560 11980 14572
rect 12032 14600 12038 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 12032 14572 12265 14600
rect 12032 14560 12038 14572
rect 12253 14569 12265 14572
rect 12299 14600 12311 14603
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 12299 14572 12633 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12621 14569 12633 14572
rect 12667 14600 12679 14603
rect 13722 14600 13728 14612
rect 12667 14572 13728 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 13722 14560 13728 14572
rect 13780 14600 13786 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13780 14572 14105 14600
rect 13780 14560 13786 14572
rect 14093 14569 14105 14572
rect 14139 14600 14151 14603
rect 14461 14603 14519 14609
rect 14461 14600 14473 14603
rect 14139 14572 14473 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14461 14569 14473 14572
rect 14507 14569 14519 14603
rect 14461 14563 14519 14569
rect 13262 14532 13268 14544
rect 13223 14504 13268 14532
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 10643 14436 11008 14464
rect 14476 14464 14504 14563
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 17954 14600 17960 14612
rect 14884 14572 17960 14600
rect 14884 14560 14890 14572
rect 17954 14560 17960 14572
rect 18012 14600 18018 14612
rect 18012 14572 18460 14600
rect 18012 14560 18018 14572
rect 14829 14467 14887 14473
rect 14829 14464 14841 14467
rect 14476 14436 14841 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 14829 14433 14841 14436
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 16474 14467 16532 14473
rect 16474 14464 16486 14467
rect 16172 14436 16486 14464
rect 16172 14424 16178 14436
rect 16474 14433 16486 14436
rect 16520 14433 16532 14467
rect 16474 14427 16532 14433
rect 18432 14405 18460 14572
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 15085 14399 15143 14405
rect 7423 14368 12296 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 7300 14300 7420 14328
rect 5261 14291 5319 14297
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5721 14263 5779 14269
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 7006 14260 7012 14272
rect 5767 14232 7012 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7282 14260 7288 14272
rect 7243 14232 7288 14260
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 7392 14260 7420 14300
rect 9950 14288 9956 14340
rect 10008 14328 10014 14340
rect 10330 14331 10388 14337
rect 10330 14328 10342 14331
rect 10008 14300 10342 14328
rect 10008 14288 10014 14300
rect 10330 14297 10342 14300
rect 10376 14297 10388 14331
rect 12268 14328 12296 14368
rect 15085 14365 15097 14399
rect 15131 14396 15143 14399
rect 18417 14399 18475 14405
rect 15131 14368 15240 14396
rect 15131 14365 15148 14368
rect 15085 14364 15148 14365
rect 15085 14359 15143 14364
rect 12342 14328 12348 14340
rect 12268 14300 12348 14328
rect 10330 14291 10388 14297
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 12989 14331 13047 14337
rect 12989 14297 13001 14331
rect 13035 14328 13047 14331
rect 14826 14328 14832 14340
rect 13035 14300 14832 14328
rect 13035 14297 13047 14300
rect 12989 14291 13047 14297
rect 14826 14288 14832 14300
rect 14884 14288 14890 14340
rect 12526 14260 12532 14272
rect 7392 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12894 14260 12900 14272
rect 12676 14232 12900 14260
rect 12676 14220 12682 14232
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15212 14260 15240 14368
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 19518 14396 19524 14408
rect 19475 14368 19524 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 16730 14331 16788 14337
rect 16730 14328 16742 14331
rect 16224 14300 16742 14328
rect 15160 14232 15240 14260
rect 15160 14220 15166 14232
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 16224 14269 16252 14300
rect 16730 14297 16742 14300
rect 16776 14297 16788 14331
rect 16730 14291 16788 14297
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 18708 14328 18736 14359
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 19978 14356 19984 14408
rect 20036 14396 20042 14408
rect 21266 14396 21272 14408
rect 20036 14368 21272 14396
rect 20036 14356 20042 14368
rect 21266 14356 21272 14368
rect 21324 14396 21330 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 21324 14368 21373 14396
rect 21324 14356 21330 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 20990 14328 20996 14340
rect 17000 14300 18736 14328
rect 18892 14300 20996 14328
rect 17000 14288 17006 14300
rect 16209 14263 16267 14269
rect 16209 14260 16221 14263
rect 15988 14232 16221 14260
rect 15988 14220 15994 14232
rect 16209 14229 16221 14232
rect 16255 14229 16267 14263
rect 17862 14260 17868 14272
rect 17823 14232 17868 14260
rect 16209 14223 16267 14229
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18230 14260 18236 14272
rect 18191 14232 18236 14260
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18892 14269 18920 14300
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 21116 14331 21174 14337
rect 21116 14297 21128 14331
rect 21162 14328 21174 14331
rect 21542 14328 21548 14340
rect 21162 14300 21548 14328
rect 21162 14297 21174 14300
rect 21116 14291 21174 14297
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 18877 14263 18935 14269
rect 18877 14229 18889 14263
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19300 14232 19625 14260
rect 19300 14220 19306 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19852 14232 19993 14260
rect 19852 14220 19858 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 4338 14016 4344 14068
rect 4396 14056 4402 14068
rect 4982 14056 4988 14068
rect 4396 14028 4988 14056
rect 4396 14016 4402 14028
rect 4982 14016 4988 14028
rect 5040 14056 5046 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 5040 14028 5181 14056
rect 5040 14016 5046 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 5169 14019 5227 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10962 14056 10968 14068
rect 10875 14028 10968 14056
rect 10962 14016 10968 14028
rect 11020 14056 11026 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11020 14028 11621 14056
rect 11020 14016 11026 14028
rect 11609 14025 11621 14028
rect 11655 14056 11667 14059
rect 11974 14056 11980 14068
rect 11655 14028 11980 14056
rect 11655 14025 11667 14028
rect 11609 14019 11667 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 13630 14016 13636 14068
rect 13688 14056 13694 14068
rect 15930 14056 15936 14068
rect 13688 14028 15936 14056
rect 13688 14016 13694 14028
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16114 14056 16120 14068
rect 16071 14028 16120 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18322 14056 18328 14068
rect 18095 14028 18328 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 20622 14056 20628 14068
rect 19628 14028 20628 14056
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 4801 13991 4859 13997
rect 4801 13988 4813 13991
rect 4672 13960 4813 13988
rect 4672 13948 4678 13960
rect 4801 13957 4813 13960
rect 4847 13957 4859 13991
rect 4801 13951 4859 13957
rect 5442 13948 5448 14000
rect 5500 13988 5506 14000
rect 11698 13988 11704 14000
rect 5500 13960 11704 13988
rect 5500 13948 5506 13960
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 12526 13948 12532 14000
rect 12584 13988 12590 14000
rect 12866 13991 12924 13997
rect 12866 13988 12878 13991
rect 12584 13960 12878 13988
rect 12584 13948 12590 13960
rect 12866 13957 12878 13960
rect 12912 13957 12924 13991
rect 12866 13951 12924 13957
rect 12986 13948 12992 14000
rect 13044 13988 13050 14000
rect 13538 13988 13544 14000
rect 13044 13960 13544 13988
rect 13044 13948 13050 13960
rect 13538 13948 13544 13960
rect 13596 13988 13602 14000
rect 16936 13991 16994 13997
rect 13596 13960 14228 13988
rect 13596 13948 13602 13960
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 10042 13920 10048 13932
rect 5316 13892 10048 13920
rect 5316 13880 5322 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10318 13920 10324 13932
rect 10376 13929 10382 13932
rect 10288 13892 10324 13920
rect 10318 13880 10324 13892
rect 10376 13883 10388 13929
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10962 13920 10968 13932
rect 10643 13892 10968 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10376 13880 10382 13883
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12253 13923 12311 13929
rect 12253 13920 12265 13923
rect 12032 13892 12265 13920
rect 12032 13880 12038 13892
rect 12253 13889 12265 13892
rect 12299 13920 12311 13923
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12299 13892 12633 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 13814 13920 13820 13932
rect 12621 13883 12679 13889
rect 12728 13892 13820 13920
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 6546 13852 6552 13864
rect 4120 13824 6552 13852
rect 4120 13812 4126 13824
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 12728 13852 12756 13892
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 11296 13824 12756 13852
rect 14200 13852 14228 13960
rect 16936 13957 16948 13991
rect 16982 13988 16994 13991
rect 17402 13988 17408 14000
rect 16982 13960 17408 13988
rect 16982 13957 16994 13960
rect 16936 13951 16994 13957
rect 17402 13948 17408 13960
rect 17460 13988 17466 14000
rect 17862 13988 17868 14000
rect 17460 13960 17868 13988
rect 17460 13948 17466 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 19628 13988 19656 14028
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 21082 14056 21088 14068
rect 20864 14028 21088 14056
rect 20864 14016 20870 14028
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 18340 13960 19656 13988
rect 15401 13923 15459 13929
rect 15401 13889 15413 13923
rect 15447 13920 15459 13923
rect 15562 13920 15568 13932
rect 15447 13892 15568 13920
rect 15447 13889 15459 13892
rect 15401 13883 15459 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 16114 13920 16120 13932
rect 15703 13892 16120 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 16114 13880 16120 13892
rect 16172 13920 16178 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16172 13892 16681 13920
rect 16172 13880 16178 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 14200 13824 14320 13852
rect 11296 13812 11302 13824
rect 9306 13784 9312 13796
rect 5460 13756 9312 13784
rect 5460 13728 5488 13756
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 14292 13793 14320 13824
rect 18340 13793 18368 13960
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 19438 13923 19496 13929
rect 19438 13920 19450 13923
rect 19024 13892 19450 13920
rect 19024 13880 19030 13892
rect 19438 13889 19450 13892
rect 19484 13889 19496 13923
rect 19438 13883 19496 13889
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13920 19763 13923
rect 19978 13920 19984 13932
rect 19751 13892 19984 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 21105 13923 21163 13929
rect 21105 13889 21117 13923
rect 21151 13920 21163 13923
rect 21151 13892 21312 13920
rect 21151 13889 21163 13892
rect 21105 13883 21163 13889
rect 21284 13852 21312 13892
rect 21358 13880 21364 13932
rect 21416 13920 21422 13932
rect 21416 13892 21461 13920
rect 21416 13880 21422 13892
rect 22094 13852 22100 13864
rect 21284 13824 22100 13852
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 14277 13787 14335 13793
rect 14277 13753 14289 13787
rect 14323 13753 14335 13787
rect 14277 13747 14335 13753
rect 18325 13787 18383 13793
rect 18325 13753 18337 13787
rect 18371 13753 18383 13787
rect 18325 13747 18383 13753
rect 5442 13676 5448 13728
rect 5500 13676 5506 13728
rect 7837 13719 7895 13725
rect 7837 13685 7849 13719
rect 7883 13716 7895 13719
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7883 13688 8217 13716
rect 7883 13685 7895 13688
rect 7837 13679 7895 13685
rect 8205 13685 8217 13688
rect 8251 13716 8263 13719
rect 8573 13719 8631 13725
rect 8573 13716 8585 13719
rect 8251 13688 8585 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8573 13685 8585 13688
rect 8619 13716 8631 13719
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8619 13688 8953 13716
rect 8619 13685 8631 13688
rect 8573 13679 8631 13685
rect 8941 13685 8953 13688
rect 8987 13716 8999 13719
rect 9122 13716 9128 13728
rect 8987 13688 9128 13716
rect 8987 13685 8999 13688
rect 8941 13679 8999 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 10410 13716 10416 13728
rect 9916 13688 10416 13716
rect 9916 13676 9922 13688
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13688 13688 14013 13716
rect 13688 13676 13694 13688
rect 14001 13685 14013 13688
rect 14047 13716 14059 13719
rect 14734 13716 14740 13728
rect 14047 13688 14740 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 16206 13716 16212 13728
rect 15344 13688 16212 13716
rect 15344 13676 15350 13688
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 19978 13716 19984 13728
rect 19939 13688 19984 13716
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 21082 13676 21088 13728
rect 21140 13716 21146 13728
rect 22002 13716 22008 13728
rect 21140 13688 22008 13716
rect 21140 13676 21146 13688
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 10689 13515 10747 13521
rect 6880 13484 10456 13512
rect 6880 13472 6886 13484
rect 10428 13453 10456 13484
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 10778 13512 10784 13524
rect 10735 13484 10784 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 15286 13512 15292 13524
rect 11756 13484 15292 13512
rect 11756 13472 11762 13484
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 17589 13515 17647 13521
rect 17589 13512 17601 13515
rect 16080 13484 17601 13512
rect 16080 13472 16086 13484
rect 17589 13481 17601 13484
rect 17635 13481 17647 13515
rect 17589 13475 17647 13481
rect 18325 13515 18383 13521
rect 18325 13481 18337 13515
rect 18371 13512 18383 13515
rect 19058 13512 19064 13524
rect 18371 13484 19064 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 10413 13447 10471 13453
rect 10413 13413 10425 13447
rect 10459 13444 10471 13447
rect 15841 13447 15899 13453
rect 10459 13416 11100 13444
rect 10459 13413 10471 13416
rect 10413 13407 10471 13413
rect 5074 13376 5080 13388
rect 5035 13348 5080 13376
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 5224 13348 5273 13376
rect 5224 13336 5230 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 5261 13339 5319 13345
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 9030 13308 9036 13320
rect 7239 13280 9036 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 11072 13308 11100 13416
rect 15841 13413 15853 13447
rect 15887 13444 15899 13447
rect 16114 13444 16120 13456
rect 15887 13416 16120 13444
rect 15887 13413 15899 13416
rect 15841 13407 15899 13413
rect 13722 13376 13728 13388
rect 13683 13348 13728 13376
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13376 15531 13379
rect 15856 13376 15884 13407
rect 16114 13404 16120 13416
rect 16172 13444 16178 13456
rect 16172 13416 16252 13444
rect 16172 13404 16178 13416
rect 16224 13385 16252 13416
rect 15519 13348 15884 13376
rect 16209 13379 16267 13385
rect 15519 13345 15531 13348
rect 15473 13339 15531 13345
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 17604 13376 17632 13475
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 20254 13512 20260 13524
rect 19306 13484 20260 13512
rect 18414 13404 18420 13456
rect 18472 13444 18478 13456
rect 18693 13447 18751 13453
rect 18693 13444 18705 13447
rect 18472 13416 18705 13444
rect 18472 13404 18478 13416
rect 18693 13413 18705 13416
rect 18739 13413 18751 13447
rect 18693 13407 18751 13413
rect 19306 13376 19334 13484
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 21269 13515 21327 13521
rect 21269 13481 21281 13515
rect 21315 13512 21327 13515
rect 21358 13512 21364 13524
rect 21315 13484 21364 13512
rect 21315 13481 21327 13484
rect 21269 13475 21327 13481
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 17604 13348 19334 13376
rect 20625 13379 20683 13385
rect 16209 13339 16267 13345
rect 20625 13345 20637 13379
rect 20671 13376 20683 13379
rect 21266 13376 21272 13388
rect 20671 13348 21272 13376
rect 20671 13345 20683 13348
rect 20625 13339 20683 13345
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 11072 13280 11845 13308
rect 5353 13243 5411 13249
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 7460 13243 7518 13249
rect 5399 13212 6132 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 5718 13172 5724 13184
rect 5679 13144 5724 13172
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 6104 13181 6132 13212
rect 7460 13209 7472 13243
rect 7506 13240 7518 13243
rect 7650 13240 7656 13252
rect 7506 13212 7656 13240
rect 7506 13209 7518 13212
rect 7460 13203 7518 13209
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 9306 13249 9312 13252
rect 9300 13203 9312 13249
rect 9364 13240 9370 13252
rect 11817 13249 11845 13280
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 12032 13280 12081 13308
rect 12032 13268 12038 13280
rect 12069 13277 12081 13280
rect 12115 13277 12127 13311
rect 16758 13308 16764 13320
rect 12069 13271 12127 13277
rect 13832 13280 16764 13308
rect 11817 13243 11882 13249
rect 9364 13212 9400 13240
rect 11817 13212 11836 13243
rect 9306 13200 9312 13203
rect 9364 13200 9370 13212
rect 11824 13209 11836 13212
rect 11870 13240 11882 13243
rect 12618 13240 12624 13252
rect 11870 13212 12624 13240
rect 11870 13209 11882 13212
rect 11824 13203 11882 13209
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 13469 13243 13527 13249
rect 13469 13209 13481 13243
rect 13515 13240 13527 13243
rect 13515 13212 13584 13240
rect 13515 13209 13527 13212
rect 13469 13203 13527 13209
rect 6089 13175 6147 13181
rect 6089 13141 6101 13175
rect 6135 13172 6147 13175
rect 7374 13172 7380 13184
rect 6135 13144 7380 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 9858 13172 9864 13184
rect 8619 13144 9864 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 11974 13172 11980 13184
rect 10008 13144 11980 13172
rect 10008 13132 10014 13144
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12345 13175 12403 13181
rect 12345 13172 12357 13175
rect 12216 13144 12357 13172
rect 12216 13132 12222 13144
rect 12345 13141 12357 13144
rect 12391 13141 12403 13175
rect 13556 13172 13584 13212
rect 13832 13172 13860 13280
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17736 13280 18153 13308
rect 17736 13268 17742 13280
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 20530 13308 20536 13320
rect 18923 13280 20536 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 21048 13280 21097 13308
rect 21048 13268 21054 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 15206 13243 15264 13249
rect 15206 13240 15218 13243
rect 14792 13212 15218 13240
rect 14792 13200 14798 13212
rect 15206 13209 15218 13212
rect 15252 13209 15264 13243
rect 15206 13203 15264 13209
rect 16476 13243 16534 13249
rect 16476 13209 16488 13243
rect 16522 13240 16534 13243
rect 17862 13240 17868 13252
rect 16522 13212 17868 13240
rect 16522 13209 16534 13212
rect 16476 13203 16534 13209
rect 17862 13200 17868 13212
rect 17920 13240 17926 13252
rect 19978 13240 19984 13252
rect 17920 13212 19984 13240
rect 17920 13200 17926 13212
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20254 13200 20260 13252
rect 20312 13240 20318 13252
rect 20358 13243 20416 13249
rect 20358 13240 20370 13243
rect 20312 13212 20370 13240
rect 20312 13200 20318 13212
rect 20358 13209 20370 13212
rect 20404 13209 20416 13243
rect 20358 13203 20416 13209
rect 13556 13144 13860 13172
rect 14093 13175 14151 13181
rect 12345 13135 12403 13141
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14458 13172 14464 13184
rect 14139 13144 14464 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 15620 13144 19257 13172
rect 15620 13132 15626 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 5261 12971 5319 12977
rect 5261 12937 5273 12971
rect 5307 12968 5319 12971
rect 5718 12968 5724 12980
rect 5307 12940 5724 12968
rect 5307 12937 5319 12940
rect 5261 12931 5319 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 10134 12968 10140 12980
rect 7883 12940 10140 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10560 12940 14596 12968
rect 10560 12928 10566 12940
rect 5353 12903 5411 12909
rect 5353 12869 5365 12903
rect 5399 12900 5411 12903
rect 5534 12900 5540 12912
rect 5399 12872 5540 12900
rect 5399 12869 5411 12872
rect 5353 12863 5411 12869
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 9030 12900 9036 12912
rect 6472 12872 9036 12900
rect 6472 12841 6500 12872
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 8128 12841 8156 12872
rect 9030 12860 9036 12872
rect 9088 12900 9094 12912
rect 11606 12900 11612 12912
rect 9088 12872 11612 12900
rect 9088 12860 9094 12872
rect 6713 12835 6771 12841
rect 6713 12832 6725 12835
rect 6604 12804 6725 12832
rect 6604 12792 6610 12804
rect 6713 12801 6725 12804
rect 6759 12801 6771 12835
rect 6713 12795 6771 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8380 12835 8438 12841
rect 8380 12801 8392 12835
rect 8426 12832 8438 12835
rect 9214 12832 9220 12844
rect 8426 12804 9220 12832
rect 8426 12801 8438 12804
rect 8380 12795 8438 12801
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9784 12841 9812 12872
rect 11606 12860 11612 12872
rect 11664 12900 11670 12912
rect 12253 12903 12311 12909
rect 12253 12900 12265 12903
rect 11664 12872 12265 12900
rect 11664 12860 11670 12872
rect 12253 12869 12265 12872
rect 12299 12900 12311 12903
rect 12621 12903 12679 12909
rect 12621 12900 12633 12903
rect 12299 12872 12633 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 12621 12869 12633 12872
rect 12667 12900 12679 12903
rect 13722 12900 13728 12912
rect 12667 12872 13728 12900
rect 12667 12869 12679 12872
rect 12621 12863 12679 12869
rect 13722 12860 13728 12872
rect 13780 12900 13786 12912
rect 13780 12872 14320 12900
rect 13780 12860 13786 12872
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 10036 12835 10094 12841
rect 10036 12832 10048 12835
rect 9769 12795 9827 12801
rect 9876 12804 10048 12832
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5442 12764 5448 12776
rect 5215 12736 5448 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 9876 12764 9904 12804
rect 10036 12801 10048 12804
rect 10082 12832 10094 12835
rect 12066 12832 12072 12844
rect 10082 12804 12072 12832
rect 10082 12801 10094 12804
rect 10036 12795 10094 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 14292 12841 14320 12872
rect 14021 12835 14079 12841
rect 12406 12804 13124 12832
rect 9508 12736 9904 12764
rect 5718 12696 5724 12708
rect 5679 12668 5724 12696
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 9508 12705 9536 12736
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12406 12764 12434 12804
rect 12032 12736 12434 12764
rect 12032 12724 12038 12736
rect 9493 12699 9551 12705
rect 9493 12665 9505 12699
rect 9539 12665 9551 12699
rect 9493 12659 9551 12665
rect 10704 12668 12572 12696
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9950 12628 9956 12640
rect 8536 12600 9956 12628
rect 8536 12588 8542 12600
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10704 12628 10732 12668
rect 11146 12628 11152 12640
rect 10100 12600 10732 12628
rect 11107 12600 11152 12628
rect 10100 12588 10106 12600
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 12544 12628 12572 12668
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12544 12600 12909 12628
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 13096 12628 13124 12804
rect 14021 12801 14033 12835
rect 14067 12832 14079 12835
rect 14277 12835 14335 12841
rect 14067 12804 14228 12832
rect 14067 12801 14079 12804
rect 14021 12795 14079 12801
rect 14200 12764 14228 12804
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14458 12764 14464 12776
rect 14200 12736 14464 12764
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 14568 12696 14596 12940
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16172 12940 16221 12968
rect 16172 12928 16178 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 17782 12903 17840 12909
rect 17782 12900 17794 12903
rect 14792 12872 17794 12900
rect 14792 12860 14798 12872
rect 17782 12869 17794 12872
rect 17828 12869 17840 12903
rect 17782 12863 17840 12869
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 19058 12900 19064 12912
rect 18196 12872 19064 12900
rect 18196 12860 18202 12872
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 21094 12903 21152 12909
rect 21094 12900 21106 12903
rect 20680 12872 21106 12900
rect 20680 12860 20686 12872
rect 21094 12869 21106 12872
rect 21140 12900 21152 12903
rect 22922 12900 22928 12912
rect 21140 12872 22928 12900
rect 21140 12869 21152 12872
rect 21094 12863 21152 12869
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15666 12835 15724 12841
rect 15666 12832 15678 12835
rect 15436 12804 15678 12832
rect 15436 12792 15442 12804
rect 15666 12801 15678 12804
rect 15712 12801 15724 12835
rect 15666 12795 15724 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16114 12832 16120 12844
rect 15979 12804 16120 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16114 12792 16120 12804
rect 16172 12832 16178 12844
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 16172 12804 18061 12832
rect 16172 12792 16178 12804
rect 18049 12801 18061 12804
rect 18095 12832 18107 12835
rect 18230 12832 18236 12844
rect 18095 12804 18236 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18230 12792 18236 12804
rect 18288 12832 18294 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18288 12804 18337 12832
rect 18288 12792 18294 12804
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 18414 12832 18420 12844
rect 18371 12804 18420 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18592 12835 18650 12841
rect 18592 12801 18604 12835
rect 18638 12832 18650 12835
rect 19794 12832 19800 12844
rect 18638 12804 19800 12832
rect 18638 12801 18650 12804
rect 18592 12795 18650 12801
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 21324 12804 21373 12832
rect 21324 12792 21330 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 19705 12699 19763 12705
rect 14568 12668 14688 12696
rect 14553 12631 14611 12637
rect 14553 12628 14565 12631
rect 13096 12600 14565 12628
rect 12897 12591 12955 12597
rect 14553 12597 14565 12600
rect 14599 12597 14611 12631
rect 14660 12628 14688 12668
rect 19705 12665 19717 12699
rect 19751 12696 19763 12699
rect 20162 12696 20168 12708
rect 19751 12668 20168 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 20162 12656 20168 12668
rect 20220 12656 20226 12708
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 14660 12600 16681 12628
rect 14553 12591 14611 12597
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 19978 12628 19984 12640
rect 19939 12600 19984 12628
rect 16669 12591 16727 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 7834 12424 7840 12436
rect 6656 12396 7840 12424
rect 5537 12359 5595 12365
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 6546 12356 6552 12368
rect 5583 12328 6552 12356
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 6546 12316 6552 12328
rect 6604 12356 6610 12368
rect 6656 12356 6684 12396
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8294 12424 8300 12436
rect 7984 12396 8300 12424
rect 7984 12384 7990 12396
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 10505 12427 10563 12433
rect 10505 12424 10517 12427
rect 10376 12396 10517 12424
rect 10376 12384 10382 12396
rect 10505 12393 10517 12396
rect 10551 12424 10563 12427
rect 12989 12427 13047 12433
rect 10551 12396 12434 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 6604 12328 6684 12356
rect 6604 12316 6610 12328
rect 6656 12297 6684 12328
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 8478 12356 8484 12368
rect 8260 12328 8484 12356
rect 8260 12316 8266 12328
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12325 8631 12359
rect 12406 12356 12434 12396
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 13035 12396 13369 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13357 12393 13369 12396
rect 13403 12424 13415 12427
rect 13722 12424 13728 12436
rect 13403 12396 13728 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14734 12424 14740 12436
rect 14139 12396 14740 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 13262 12356 13268 12368
rect 12406 12328 13268 12356
rect 8573 12319 8631 12325
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6822 12288 6828 12300
rect 6783 12260 6828 12288
rect 6641 12251 6699 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 8588 12288 8616 12319
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 13538 12316 13544 12368
rect 13596 12356 13602 12368
rect 14108 12356 14136 12387
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 16172 12396 17172 12424
rect 16172 12384 16178 12396
rect 13596 12328 14136 12356
rect 13596 12316 13602 12328
rect 8588 12260 9260 12288
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 9122 12220 9128 12232
rect 7239 12192 9128 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9232 12220 9260 12260
rect 10502 12248 10508 12300
rect 10560 12288 10566 12300
rect 11146 12288 11152 12300
rect 10560 12260 11152 12288
rect 10560 12248 10566 12260
rect 11146 12248 11152 12260
rect 11204 12288 11210 12300
rect 15473 12291 15531 12297
rect 11204 12260 11376 12288
rect 11204 12248 11210 12260
rect 9381 12223 9439 12229
rect 9381 12220 9393 12223
rect 9232 12192 9393 12220
rect 9381 12189 9393 12192
rect 9427 12220 9439 12223
rect 10594 12220 10600 12232
rect 9427 12192 10600 12220
rect 9427 12189 9439 12192
rect 9381 12183 9439 12189
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 10919 12192 11253 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11348 12220 11376 12260
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15562 12288 15568 12300
rect 15519 12260 15568 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 16114 12288 16120 12300
rect 15620 12260 16120 12288
rect 15620 12248 15626 12260
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 17144 12297 17172 12396
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 19518 12424 19524 12436
rect 18472 12396 18828 12424
rect 19479 12396 19524 12424
rect 18472 12384 18478 12396
rect 17405 12359 17463 12365
rect 17405 12356 17417 12359
rect 17236 12328 17417 12356
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 11497 12223 11555 12229
rect 11497 12220 11509 12223
rect 11348 12192 11509 12220
rect 11241 12183 11299 12189
rect 11497 12189 11509 12192
rect 11543 12189 11555 12223
rect 16850 12220 16856 12232
rect 16908 12229 16914 12232
rect 16820 12192 16856 12220
rect 11497 12183 11555 12189
rect 5905 12155 5963 12161
rect 5905 12121 5917 12155
rect 5951 12152 5963 12155
rect 7460 12155 7518 12161
rect 5951 12124 6592 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6564 12093 6592 12124
rect 7460 12121 7472 12155
rect 7506 12152 7518 12155
rect 7506 12124 9352 12152
rect 7506 12121 7518 12124
rect 7460 12115 7518 12121
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 6052 12056 6193 12084
rect 6052 12044 6058 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 7374 12084 7380 12096
rect 6595 12056 7380 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 9324 12084 9352 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10778 12152 10784 12164
rect 9916 12124 10784 12152
rect 9916 12112 9922 12124
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 11256 12152 11284 12183
rect 16850 12180 16856 12192
rect 16908 12183 16920 12229
rect 16908 12180 16914 12183
rect 11606 12152 11612 12164
rect 11072 12124 11612 12152
rect 11072 12096 11100 12124
rect 11606 12112 11612 12124
rect 11664 12152 11670 12164
rect 12158 12152 12164 12164
rect 11664 12124 12164 12152
rect 11664 12112 11670 12124
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 13170 12112 13176 12164
rect 13228 12152 13234 12164
rect 15206 12155 15264 12161
rect 15206 12152 15218 12155
rect 13228 12124 15218 12152
rect 13228 12112 13234 12124
rect 15206 12121 15218 12124
rect 15252 12152 15264 12155
rect 17236 12152 17264 12328
rect 17405 12325 17417 12328
rect 17451 12325 17463 12359
rect 17405 12319 17463 12325
rect 18800 12297 18828 12396
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 18785 12291 18843 12297
rect 18785 12257 18797 12291
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 15252 12124 17264 12152
rect 17328 12192 19717 12220
rect 15252 12121 15264 12124
rect 15206 12115 15264 12121
rect 10042 12084 10048 12096
rect 9324 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 11054 12044 11060 12096
rect 11112 12044 11118 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11974 12084 11980 12096
rect 11204 12056 11980 12084
rect 11204 12044 11210 12056
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12621 12087 12679 12093
rect 12621 12084 12633 12087
rect 12584 12056 12633 12084
rect 12584 12044 12590 12056
rect 12621 12053 12633 12056
rect 12667 12053 12679 12087
rect 12621 12047 12679 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15102 12084 15108 12096
rect 14792 12056 15108 12084
rect 14792 12044 14798 12056
rect 15102 12044 15108 12056
rect 15160 12084 15166 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15160 12056 15761 12084
rect 15160 12044 15166 12056
rect 15749 12053 15761 12056
rect 15795 12053 15807 12087
rect 15749 12047 15807 12053
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 17328 12084 17356 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21324 12192 21373 12220
rect 21324 12180 21330 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 18414 12112 18420 12164
rect 18472 12152 18478 12164
rect 18518 12155 18576 12161
rect 18518 12152 18530 12155
rect 18472 12124 18530 12152
rect 18472 12112 18478 12124
rect 18518 12121 18530 12124
rect 18564 12121 18576 12155
rect 18518 12115 18576 12121
rect 21116 12155 21174 12161
rect 21116 12121 21128 12155
rect 21162 12152 21174 12155
rect 22370 12152 22376 12164
rect 21162 12124 22376 12152
rect 21162 12121 21174 12124
rect 21116 12115 21174 12121
rect 22370 12112 22376 12124
rect 22428 12112 22434 12164
rect 16172 12056 17356 12084
rect 16172 12044 16178 12056
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18322 12084 18328 12096
rect 18012 12056 18328 12084
rect 18012 12044 18018 12056
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19024 12056 19993 12084
rect 19024 12044 19030 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6788 11852 7021 11880
rect 6788 11840 6794 11852
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 7009 11843 7067 11849
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 7742 11880 7748 11892
rect 7524 11852 7748 11880
rect 7524 11840 7530 11852
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 8076 11852 8125 11880
rect 8076 11840 8082 11852
rect 8113 11849 8125 11852
rect 8159 11849 8171 11883
rect 11514 11880 11520 11892
rect 8113 11843 8171 11849
rect 8404 11852 11520 11880
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 5629 11815 5687 11821
rect 5629 11812 5641 11815
rect 5592 11784 5641 11812
rect 5592 11772 5598 11784
rect 5629 11781 5641 11784
rect 5675 11781 5687 11815
rect 8404 11812 8432 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11609 11883 11667 11889
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 12158 11880 12164 11892
rect 11655 11852 12164 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12894 11880 12900 11892
rect 12855 11852 12900 11880
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 14366 11880 14372 11892
rect 14327 11852 14372 11880
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 15286 11880 15292 11892
rect 14700 11852 15292 11880
rect 14700 11840 14706 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 15896 11852 17049 11880
rect 15896 11840 15902 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 17678 11880 17684 11892
rect 17639 11852 17684 11880
rect 17037 11843 17095 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18046 11880 18052 11892
rect 17788 11852 18052 11880
rect 5629 11775 5687 11781
rect 7300 11784 8432 11812
rect 8481 11815 8539 11821
rect 7300 11744 7328 11784
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 10873 11815 10931 11821
rect 10873 11812 10885 11815
rect 8527 11784 10885 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 10873 11781 10885 11784
rect 10919 11781 10931 11815
rect 17788 11812 17816 11852
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18230 11840 18236 11892
rect 18288 11840 18294 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 21358 11880 21364 11892
rect 19392 11852 21364 11880
rect 19392 11840 19398 11852
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 18248 11812 18276 11840
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 10873 11775 10931 11781
rect 16316 11784 17816 11812
rect 17972 11784 19625 11812
rect 5460 11716 7328 11744
rect 7377 11747 7435 11753
rect 5460 11685 5488 11716
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7834 11744 7840 11756
rect 7423 11716 7840 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8018 11704 8024 11756
rect 8076 11744 8082 11756
rect 9858 11744 9864 11756
rect 8076 11716 9864 11744
rect 8076 11704 8082 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10318 11744 10324 11756
rect 10376 11753 10382 11756
rect 10376 11747 10399 11753
rect 10251 11716 10324 11744
rect 10318 11704 10324 11716
rect 10387 11744 10399 11747
rect 10778 11744 10784 11756
rect 10387 11716 10784 11744
rect 10387 11713 10399 11716
rect 10376 11707 10399 11713
rect 10376 11704 10382 11707
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11054 11744 11060 11756
rect 10888 11716 11060 11744
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 6733 11679 6791 11685
rect 6733 11645 6745 11679
rect 6779 11676 6791 11679
rect 7190 11676 7196 11688
rect 6779 11648 7196 11676
rect 6779 11645 6791 11648
rect 6733 11639 6791 11645
rect 4522 11568 4528 11620
rect 4580 11608 4586 11620
rect 5552 11608 5580 11639
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7466 11676 7472 11688
rect 7427 11648 7472 11676
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8386 11676 8392 11688
rect 7699 11648 8392 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 10597 11679 10655 11685
rect 8803 11648 9628 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 4580 11580 5580 11608
rect 4580 11568 4586 11580
rect 4908 11552 4936 11580
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6914 11540 6920 11552
rect 6043 11512 6920 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 9217 11543 9275 11549
rect 9217 11509 9229 11543
rect 9263 11540 9275 11543
rect 9306 11540 9312 11552
rect 9263 11512 9312 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9600 11540 9628 11648
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 10888 11676 10916 11716
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11480 11716 11897 11744
rect 11480 11704 11486 11716
rect 11885 11713 11897 11716
rect 11931 11744 11943 11747
rect 11974 11744 11980 11756
rect 11931 11716 11980 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 11974 11704 11980 11716
rect 12032 11744 12038 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12032 11716 12265 11744
rect 12032 11704 12038 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 14366 11744 14372 11756
rect 13311 11716 14372 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 15194 11744 15200 11756
rect 14783 11716 15200 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 16316 11753 16344 11784
rect 17972 11756 18000 11784
rect 19613 11781 19625 11784
rect 19659 11781 19671 11815
rect 19613 11775 19671 11781
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16390 11744 16396 11756
rect 16347 11716 16396 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 17126 11704 17132 11756
rect 17184 11704 17190 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11713 17279 11747
rect 17494 11744 17500 11756
rect 17455 11716 17500 11744
rect 17221 11707 17279 11713
rect 10643 11648 10916 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 12216 11648 13369 11676
rect 12216 11636 12222 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 11054 11568 11060 11620
rect 11112 11568 11118 11620
rect 13464 11608 13492 11639
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13780 11648 13921 11676
rect 13780 11636 13786 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 13909 11639 13967 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 17144 11676 17172 11704
rect 14967 11648 17172 11676
rect 17236 11676 17264 11707
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18230 11753 18236 11756
rect 18224 11744 18236 11753
rect 18012 11716 18105 11744
rect 18191 11716 18236 11744
rect 18012 11704 18018 11716
rect 18224 11707 18236 11716
rect 18230 11704 18236 11707
rect 18288 11704 18294 11756
rect 19628 11744 19656 11775
rect 20162 11772 20168 11824
rect 20220 11821 20226 11824
rect 20220 11815 20284 11821
rect 20220 11781 20238 11815
rect 20272 11781 20284 11815
rect 20220 11775 20284 11781
rect 20220 11772 20226 11775
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19628 11716 19993 11744
rect 19981 11713 19993 11716
rect 20027 11744 20039 11747
rect 21266 11744 21272 11756
rect 20027 11716 21272 11744
rect 20027 11713 20039 11716
rect 19981 11707 20039 11713
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 17770 11676 17776 11688
rect 17236 11648 17776 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 13372 11580 13492 11608
rect 9674 11540 9680 11552
rect 9600 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11072 11540 11100 11568
rect 10928 11512 11100 11540
rect 10928 11500 10934 11512
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 12434 11540 12440 11552
rect 11664 11512 12440 11540
rect 11664 11500 11670 11512
rect 12434 11500 12440 11512
rect 12492 11540 12498 11552
rect 13372 11540 13400 11580
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14936 11608 14964 11639
rect 14240 11580 14964 11608
rect 14240 11568 14246 11580
rect 15378 11568 15384 11620
rect 15436 11608 15442 11620
rect 15562 11608 15568 11620
rect 15436 11580 15568 11608
rect 15436 11568 15442 11580
rect 15562 11568 15568 11580
rect 15620 11608 15626 11620
rect 16669 11611 16727 11617
rect 16669 11608 16681 11611
rect 15620 11580 16681 11608
rect 15620 11568 15626 11580
rect 16669 11577 16681 11580
rect 16715 11608 16727 11611
rect 17126 11608 17132 11620
rect 16715 11580 17132 11608
rect 16715 11577 16727 11580
rect 16669 11571 16727 11577
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 12492 11512 13400 11540
rect 12492 11500 12498 11512
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 15010 11540 15016 11552
rect 13504 11512 15016 11540
rect 13504 11500 13510 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 15344 11512 16129 11540
rect 15344 11500 15350 11512
rect 16117 11509 16129 11512
rect 16163 11509 16175 11543
rect 16117 11503 16175 11509
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 17236 11540 17264 11648
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 19978 11608 19984 11620
rect 19260 11580 19984 11608
rect 16264 11512 17264 11540
rect 16264 11500 16270 11512
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18230 11540 18236 11552
rect 17828 11512 18236 11540
rect 17828 11500 17834 11512
rect 18230 11500 18236 11512
rect 18288 11540 18294 11552
rect 19260 11540 19288 11580
rect 19978 11568 19984 11580
rect 20036 11568 20042 11620
rect 22738 11608 22744 11620
rect 20916 11580 22744 11608
rect 18288 11512 19288 11540
rect 19337 11543 19395 11549
rect 18288 11500 18294 11512
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 19794 11540 19800 11552
rect 19383 11512 19800 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 19794 11500 19800 11512
rect 19852 11540 19858 11552
rect 20916 11540 20944 11580
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 19852 11512 20944 11540
rect 21361 11543 21419 11549
rect 19852 11500 19858 11512
rect 21361 11509 21373 11543
rect 21407 11540 21419 11543
rect 21542 11540 21548 11552
rect 21407 11512 21548 11540
rect 21407 11509 21419 11512
rect 21361 11503 21419 11509
rect 21542 11500 21548 11512
rect 21600 11500 21606 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 7282 11336 7288 11348
rect 6595 11308 7288 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7558 11336 7564 11348
rect 7519 11308 7564 11336
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 11606 11336 11612 11348
rect 8128 11308 11612 11336
rect 8018 11268 8024 11280
rect 5920 11240 8024 11268
rect 5920 11209 5948 11240
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 6052 11172 6101 11200
rect 6052 11160 6058 11172
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 8128 11200 8156 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 13446 11336 13452 11348
rect 11900 11308 13452 11336
rect 9493 11271 9551 11277
rect 9493 11268 9505 11271
rect 8864 11240 9505 11268
rect 7055 11172 8156 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8260 11172 8401 11200
rect 8260 11160 8266 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7558 11132 7564 11144
rect 7432 11104 7564 11132
rect 7432 11092 7438 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 8864 11132 8892 11240
rect 9493 11237 9505 11240
rect 9539 11237 9551 11271
rect 9493 11231 9551 11237
rect 10796 11172 11376 11200
rect 7708 11104 8892 11132
rect 7708 11092 7714 11104
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 10796 11132 10824 11172
rect 9088 11104 10824 11132
rect 9088 11092 9094 11104
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11348 11132 11376 11172
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11572 11172 11621 11200
rect 11572 11160 11578 11172
rect 11609 11169 11621 11172
rect 11655 11200 11667 11203
rect 11900 11200 11928 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14884 11308 14933 11336
rect 14884 11296 14890 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 15194 11336 15200 11348
rect 15155 11308 15200 11336
rect 14921 11299 14979 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 17037 11339 17095 11345
rect 17037 11305 17049 11339
rect 17083 11336 17095 11339
rect 17083 11308 17816 11336
rect 17083 11305 17095 11308
rect 17037 11299 17095 11305
rect 11974 11228 11980 11280
rect 12032 11268 12038 11280
rect 12032 11240 12112 11268
rect 12032 11228 12038 11240
rect 11655 11172 11928 11200
rect 12084 11200 12112 11240
rect 12158 11228 12164 11280
rect 12216 11268 12222 11280
rect 12216 11240 12261 11268
rect 12216 11228 12222 11240
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 17788 11268 17816 11308
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 18012 11308 18797 11336
rect 18012 11296 18018 11308
rect 18785 11305 18797 11308
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 12676 11240 15884 11268
rect 17788 11240 18000 11268
rect 12676 11228 12682 11240
rect 13004 11209 13032 11240
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 12084 11172 12909 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 15746 11200 15752 11212
rect 14415 11172 14596 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 10928 11104 10973 11132
rect 11348 11128 11845 11132
rect 11348 11104 12081 11128
rect 10928 11092 10934 11104
rect 11817 11100 12081 11104
rect 5534 11064 5540 11076
rect 5495 11036 5540 11064
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 6181 11067 6239 11073
rect 6181 11033 6193 11067
rect 6227 11064 6239 11067
rect 6227 11036 6868 11064
rect 6227 11033 6239 11036
rect 6181 11027 6239 11033
rect 6840 10996 6868 11036
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 6972 11036 7113 11064
rect 6972 11024 6978 11036
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 7101 11027 7159 11033
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8251 11036 8953 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 10628 11067 10686 11073
rect 10628 11033 10640 11067
rect 10674 11064 10686 11067
rect 10674 11036 11376 11064
rect 10674 11033 10686 11036
rect 10628 11027 10686 11033
rect 7374 10996 7380 11008
rect 6840 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 8076 10968 8309 10996
rect 8076 10956 8082 10968
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 8297 10959 8355 10965
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9398 10996 9404 11008
rect 9180 10968 9404 10996
rect 9180 10956 9186 10968
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 11348 10996 11376 11036
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 12053 11064 12081 11100
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12676 11104 12817 11132
rect 12676 11092 12682 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12912 11132 12940 11163
rect 14458 11132 14464 11144
rect 12912 11104 14464 11132
rect 12805 11095 12863 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14568 11132 14596 11172
rect 15100 11172 15752 11200
rect 15100 11132 15128 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 15856 11200 15884 11240
rect 17865 11203 17923 11209
rect 17865 11200 17877 11203
rect 15856 11172 17877 11200
rect 17865 11169 17877 11172
rect 17911 11169 17923 11203
rect 17972 11200 18000 11240
rect 18322 11228 18328 11280
rect 18380 11268 18386 11280
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 18380 11240 19257 11268
rect 18380 11228 18386 11240
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 21082 11268 21088 11280
rect 19245 11231 19303 11237
rect 19904 11240 21088 11268
rect 19904 11209 19932 11240
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 19889 11203 19947 11209
rect 17972 11172 19840 11200
rect 17865 11163 17923 11169
rect 14568 11104 15128 11132
rect 16853 11135 16911 11141
rect 14568 11064 14596 11104
rect 16853 11101 16865 11135
rect 16899 11132 16911 11135
rect 17954 11132 17960 11144
rect 16899 11104 17960 11132
rect 16899 11101 16911 11104
rect 16853 11095 16911 11101
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 19518 11132 19524 11144
rect 18064 11104 19524 11132
rect 11480 11036 11744 11064
rect 12053 11036 14596 11064
rect 15565 11067 15623 11073
rect 11480 11024 11486 11036
rect 11514 10996 11520 11008
rect 11348 10968 11520 10996
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11716 11005 11744 11036
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 15838 11064 15844 11076
rect 15611 11036 15844 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 12158 10996 12164 11008
rect 11839 10968 12164 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 13446 10996 13452 11008
rect 12492 10968 12537 10996
rect 13407 10968 13452 10996
rect 12492 10956 12498 10968
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 14826 10996 14832 11008
rect 14599 10968 14832 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 15657 10999 15715 11005
rect 15657 10965 15669 10999
rect 15703 10996 15715 10999
rect 15746 10996 15752 11008
rect 15703 10968 15752 10996
rect 15703 10965 15715 10968
rect 15657 10959 15715 10965
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 17313 10999 17371 11005
rect 17313 10996 17325 10999
rect 16356 10968 17325 10996
rect 16356 10956 16362 10968
rect 17313 10965 17325 10968
rect 17359 10965 17371 10999
rect 17678 10996 17684 11008
rect 17639 10968 17684 10996
rect 17313 10959 17371 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17773 10999 17831 11005
rect 17773 10965 17785 10999
rect 17819 10996 17831 10999
rect 18064 10996 18092 11104
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 19812 11132 19840 11172
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20496 11172 20821 11200
rect 20496 11160 20502 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 21266 11200 21272 11212
rect 21227 11172 21272 11200
rect 20809 11163 20867 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 20990 11132 20996 11144
rect 19812 11104 20996 11132
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19613 11067 19671 11073
rect 19613 11064 19625 11067
rect 18748 11036 19625 11064
rect 18748 11024 18754 11036
rect 19613 11033 19625 11036
rect 19659 11033 19671 11067
rect 19613 11027 19671 11033
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20346 11064 20352 11076
rect 19751 11036 20352 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 20717 11067 20775 11073
rect 20717 11033 20729 11067
rect 20763 11064 20775 11067
rect 21358 11064 21364 11076
rect 20763 11036 21364 11064
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 21358 11024 21364 11036
rect 21416 11064 21422 11076
rect 22554 11064 22560 11076
rect 21416 11036 22560 11064
rect 21416 11024 21422 11036
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 18322 10996 18328 11008
rect 17819 10968 18092 10996
rect 18283 10968 18328 10996
rect 17819 10965 17831 10968
rect 17773 10959 17831 10965
rect 18322 10956 18328 10968
rect 18380 10956 18386 11008
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 20257 10999 20315 11005
rect 20257 10996 20269 10999
rect 20036 10968 20269 10996
rect 20036 10956 20042 10968
rect 20257 10965 20269 10968
rect 20303 10965 20315 10999
rect 20622 10996 20628 11008
rect 20583 10968 20628 10996
rect 20257 10959 20315 10965
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6454 10792 6460 10804
rect 5776 10764 6460 10792
rect 5776 10752 5782 10764
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 7374 10792 7380 10804
rect 7335 10764 7380 10792
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 8570 10792 8576 10804
rect 8343 10764 8576 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10686 10792 10692 10804
rect 10192 10764 10692 10792
rect 10192 10752 10198 10764
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 11238 10792 11244 10804
rect 11195 10764 11244 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 12342 10792 12348 10804
rect 12303 10764 12348 10792
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12492 10764 12817 10792
rect 12492 10752 12498 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 12805 10755 12863 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 16853 10795 16911 10801
rect 14476 10764 16344 10792
rect 7926 10724 7932 10736
rect 6472 10696 7932 10724
rect 6472 10597 6500 10696
rect 7926 10684 7932 10696
rect 7984 10684 7990 10736
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 10318 10724 10324 10736
rect 9907 10696 10324 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 11974 10724 11980 10736
rect 10928 10696 11980 10724
rect 10928 10684 10934 10696
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 12713 10727 12771 10733
rect 12713 10693 12725 10727
rect 12759 10724 12771 10727
rect 13078 10724 13084 10736
rect 12759 10696 13084 10724
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 9674 10656 9680 10668
rect 8711 10628 9680 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10656 9827 10659
rect 10410 10656 10416 10668
rect 9815 10628 10416 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 10827 10628 11529 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 12342 10616 12348 10668
rect 12400 10656 12406 10668
rect 14476 10656 14504 10764
rect 14737 10727 14795 10733
rect 14737 10693 14749 10727
rect 14783 10724 14795 10727
rect 15286 10724 15292 10736
rect 14783 10696 15292 10724
rect 14783 10693 14795 10696
rect 14737 10687 14795 10693
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 15657 10727 15715 10733
rect 15657 10693 15669 10727
rect 15703 10724 15715 10727
rect 16206 10724 16212 10736
rect 15703 10696 16212 10724
rect 15703 10693 15715 10696
rect 15657 10687 15715 10693
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 16316 10724 16344 10764
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 16942 10792 16948 10804
rect 16899 10764 16948 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17126 10792 17132 10804
rect 17087 10764 17132 10792
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 18322 10792 18328 10804
rect 18283 10764 18328 10792
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 18690 10792 18696 10804
rect 18651 10764 18696 10792
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 19567 10764 20269 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21361 10795 21419 10801
rect 21361 10792 21373 10795
rect 21140 10764 21373 10792
rect 21140 10752 21146 10764
rect 21361 10761 21373 10764
rect 21407 10792 21419 10795
rect 22094 10792 22100 10804
rect 21407 10764 22100 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 19613 10727 19671 10733
rect 16316 10696 19334 10724
rect 12400 10628 14504 10656
rect 15933 10659 15991 10665
rect 12400 10616 12406 10628
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 16666 10656 16672 10668
rect 16627 10628 16672 10656
rect 15933 10619 15991 10625
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10557 6515 10591
rect 6638 10588 6644 10600
rect 6599 10560 6644 10588
rect 6457 10551 6515 10557
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 7800 10560 8769 10588
rect 7800 10548 7806 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9030 10588 9036 10600
rect 8987 10560 9036 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 10042 10588 10048 10600
rect 10003 10560 10048 10588
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 12897 10591 12955 10597
rect 11020 10560 12664 10588
rect 11020 10548 11026 10560
rect 7101 10523 7159 10529
rect 7101 10489 7113 10523
rect 7147 10520 7159 10523
rect 12636 10520 12664 10560
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 13538 10588 13544 10600
rect 13499 10560 13544 10588
rect 12897 10551 12955 10557
rect 12912 10520 12940 10551
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 13814 10588 13820 10600
rect 13679 10560 13820 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14424 10560 14841 10588
rect 14424 10548 14430 10560
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 15010 10588 15016 10600
rect 14971 10560 15016 10588
rect 14829 10551 14887 10557
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15948 10520 15976 10619
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17494 10656 17500 10668
rect 17000 10628 17500 10656
rect 17000 10616 17006 10628
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 18690 10656 18696 10668
rect 17972 10628 18696 10656
rect 17972 10588 18000 10628
rect 18690 10616 18696 10628
rect 18748 10656 18754 10668
rect 18966 10656 18972 10668
rect 18748 10628 18972 10656
rect 18748 10616 18754 10628
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 19306 10656 19334 10696
rect 19613 10693 19625 10727
rect 19659 10724 19671 10727
rect 19978 10724 19984 10736
rect 19659 10696 19984 10724
rect 19659 10693 19671 10696
rect 19613 10687 19671 10693
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 19794 10656 19800 10668
rect 19306 10628 19800 10656
rect 19794 10616 19800 10628
rect 19852 10656 19858 10668
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 19852 10628 20637 10656
rect 19852 10616 19858 10628
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 17512 10560 18000 10588
rect 18049 10591 18107 10597
rect 16114 10520 16120 10532
rect 7147 10492 9674 10520
rect 12636 10492 12940 10520
rect 13004 10492 15976 10520
rect 16075 10492 16120 10520
rect 7147 10489 7159 10492
rect 7101 10483 7159 10489
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5776 10424 5917 10452
rect 5776 10412 5782 10424
rect 5905 10421 5917 10424
rect 5951 10421 5963 10455
rect 8018 10452 8024 10464
rect 7979 10424 8024 10452
rect 5905 10415 5963 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 9646 10452 9674 10492
rect 13004 10452 13032 10492
rect 16114 10480 16120 10492
rect 16172 10480 16178 10532
rect 9646 10424 13032 10452
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 13596 10424 14105 10452
rect 13596 10412 13602 10424
rect 14093 10421 14105 10424
rect 14139 10421 14151 10455
rect 14093 10415 14151 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 17512 10452 17540 10560
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18230 10588 18236 10600
rect 18191 10560 18236 10588
rect 18049 10551 18107 10557
rect 18064 10520 18092 10551
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 19429 10591 19487 10597
rect 19429 10557 19441 10591
rect 19475 10588 19487 10591
rect 19702 10588 19708 10600
rect 19475 10560 19708 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20128 10560 20729 10588
rect 20128 10548 20134 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10557 20867 10591
rect 20809 10551 20867 10557
rect 18782 10520 18788 10532
rect 18064 10492 18788 10520
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 20438 10480 20444 10532
rect 20496 10520 20502 10532
rect 20824 10520 20852 10551
rect 20496 10492 20852 10520
rect 20496 10480 20502 10492
rect 17678 10452 17684 10464
rect 15252 10424 17540 10452
rect 17591 10424 17684 10452
rect 15252 10412 15258 10424
rect 17678 10412 17684 10424
rect 17736 10452 17742 10464
rect 18322 10452 18328 10464
rect 17736 10424 18328 10452
rect 17736 10412 17742 10424
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 19981 10455 20039 10461
rect 19981 10421 19993 10455
rect 20027 10452 20039 10455
rect 20070 10452 20076 10464
rect 20027 10424 20076 10452
rect 20027 10421 20039 10424
rect 19981 10415 20039 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 6822 10248 6828 10260
rect 5460 10220 6828 10248
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5460 10121 5488 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 10042 10248 10048 10260
rect 7392 10220 10048 10248
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6365 10183 6423 10189
rect 6365 10180 6377 10183
rect 5592 10152 6377 10180
rect 5592 10140 5598 10152
rect 6365 10149 6377 10152
rect 6411 10149 6423 10183
rect 6365 10143 6423 10149
rect 6454 10140 6460 10192
rect 6512 10180 6518 10192
rect 7392 10189 7420 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13354 10248 13360 10260
rect 13127 10220 13360 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13998 10248 14004 10260
rect 13657 10220 14004 10248
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 6512 10152 7389 10180
rect 6512 10140 6518 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 10134 10180 10140 10192
rect 9732 10152 10140 10180
rect 9732 10140 9738 10152
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 10873 10183 10931 10189
rect 10873 10149 10885 10183
rect 10919 10180 10931 10183
rect 13657 10180 13685 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14185 10251 14243 10257
rect 14185 10217 14197 10251
rect 14231 10248 14243 10251
rect 14458 10248 14464 10260
rect 14231 10220 14464 10248
rect 14231 10217 14243 10220
rect 14185 10211 14243 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 14918 10248 14924 10260
rect 14875 10220 14924 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 16666 10248 16672 10260
rect 15068 10220 16672 10248
rect 15068 10208 15074 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17644 10220 17693 10248
rect 17644 10208 17650 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 20806 10248 20812 10260
rect 20767 10220 20812 10248
rect 17681 10211 17739 10217
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 10919 10152 13685 10180
rect 13725 10183 13783 10189
rect 10919 10149 10931 10152
rect 10873 10143 10931 10149
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 16942 10180 16948 10192
rect 13771 10152 16948 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 17313 10183 17371 10189
rect 17313 10149 17325 10183
rect 17359 10180 17371 10183
rect 21358 10180 21364 10192
rect 17359 10152 21364 10180
rect 17359 10149 17371 10152
rect 17313 10143 17371 10149
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5408 10084 5457 10112
rect 5408 10072 5414 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 5445 10075 5503 10081
rect 6104 10084 6929 10112
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 6104 10044 6132 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 8352 10084 9229 10112
rect 8352 10072 8358 10084
rect 9217 10081 9229 10084
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 9364 10084 10241 10112
rect 9364 10072 9370 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 12529 10115 12587 10121
rect 10560 10084 11744 10112
rect 10560 10072 10566 10084
rect 5040 10016 6132 10044
rect 5040 10004 5046 10016
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6512 10016 6745 10044
rect 6512 10004 6518 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7834 10044 7840 10056
rect 6871 10016 7840 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 9539 10016 11621 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 5166 9976 5172 9988
rect 3936 9948 5172 9976
rect 3936 9936 3942 9948
rect 5166 9936 5172 9948
rect 5224 9976 5230 9988
rect 7742 9976 7748 9988
rect 5224 9948 7748 9976
rect 5224 9936 5230 9948
rect 7742 9936 7748 9948
rect 7800 9936 7806 9988
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 9766 9976 9772 9988
rect 8619 9948 9772 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10505 9979 10563 9985
rect 10505 9945 10517 9979
rect 10551 9976 10563 9979
rect 11149 9979 11207 9985
rect 11149 9976 11161 9979
rect 10551 9948 11161 9976
rect 10551 9945 10563 9948
rect 10505 9939 10563 9945
rect 11149 9945 11161 9948
rect 11195 9945 11207 9979
rect 11716 9976 11744 10084
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 13630 10112 13636 10124
rect 12575 10084 13636 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 14366 10072 14372 10124
rect 14424 10112 14430 10124
rect 15194 10112 15200 10124
rect 14424 10084 15200 10112
rect 14424 10072 14430 10084
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 15746 10112 15752 10124
rect 15707 10084 15752 10112
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 17954 10112 17960 10124
rect 16439 10084 17960 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18141 10115 18199 10121
rect 18141 10112 18153 10115
rect 18104 10084 18153 10112
rect 18104 10072 18110 10084
rect 18141 10081 18153 10084
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18506 10112 18512 10124
rect 18371 10084 18512 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 20349 10115 20407 10121
rect 18607 10084 19840 10112
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 13446 10044 13452 10056
rect 12759 10016 13452 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 15102 10044 15108 10056
rect 13780 10016 15108 10044
rect 13780 10004 13786 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 16206 10044 16212 10056
rect 15519 10016 16212 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 18607 10044 18635 10084
rect 17236 10016 18635 10044
rect 15010 9976 15016 9988
rect 11716 9948 15016 9976
rect 11149 9939 11207 9945
rect 15010 9936 15016 9948
rect 15068 9936 15074 9988
rect 17236 9976 17264 10016
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 18748 10016 18889 10044
rect 18748 10004 18754 10016
rect 18877 10013 18889 10016
rect 18923 10013 18935 10047
rect 19242 10044 19248 10056
rect 19203 10016 19248 10044
rect 18877 10007 18935 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19610 10004 19616 10056
rect 19668 10044 19674 10056
rect 19705 10047 19763 10053
rect 19705 10044 19717 10047
rect 19668 10016 19717 10044
rect 19668 10004 19674 10016
rect 19705 10013 19717 10016
rect 19751 10013 19763 10047
rect 19812 10044 19840 10084
rect 20349 10081 20361 10115
rect 20395 10112 20407 10115
rect 20622 10112 20628 10124
rect 20395 10084 20628 10112
rect 20395 10081 20407 10084
rect 20349 10075 20407 10081
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 19812 10016 21005 10044
rect 19705 10007 19763 10013
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 16776 9948 17264 9976
rect 18049 9979 18107 9985
rect 5258 9868 5264 9920
rect 5316 9908 5322 9920
rect 5629 9911 5687 9917
rect 5629 9908 5641 9911
rect 5316 9880 5641 9908
rect 5316 9868 5322 9880
rect 5629 9877 5641 9880
rect 5675 9877 5687 9911
rect 5629 9871 5687 9877
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5776 9880 5821 9908
rect 5776 9868 5782 9880
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 6052 9880 6101 9908
rect 6052 9868 6058 9880
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7616 9880 8125 9908
rect 7616 9868 7622 9880
rect 8113 9877 8125 9880
rect 8159 9908 8171 9911
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8159 9880 9413 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 9401 9877 9413 9880
rect 9447 9908 9459 9911
rect 9674 9908 9680 9920
rect 9447 9880 9680 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 11882 9908 11888 9920
rect 10459 9880 11888 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12618 9908 12624 9920
rect 12579 9880 12624 9908
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14090 9908 14096 9920
rect 13596 9880 14096 9908
rect 13596 9868 13602 9880
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 15102 9908 15108 9920
rect 15063 9880 15108 9908
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 16776 9908 16804 9948
rect 18049 9945 18061 9979
rect 18095 9976 18107 9979
rect 19150 9976 19156 9988
rect 18095 9948 19156 9976
rect 18095 9945 18107 9948
rect 18049 9939 18107 9945
rect 19150 9936 19156 9948
rect 19208 9936 19214 9988
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 21082 9976 21088 9988
rect 20864 9948 21088 9976
rect 20864 9936 20870 9948
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 16356 9880 16804 9908
rect 16853 9911 16911 9917
rect 16356 9868 16362 9880
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 17034 9908 17040 9920
rect 16899 9880 17040 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18693 9911 18751 9917
rect 18693 9908 18705 9911
rect 17644 9880 18705 9908
rect 17644 9868 17650 9880
rect 18693 9877 18705 9880
rect 18739 9877 18751 9911
rect 18693 9871 18751 9877
rect 19429 9911 19487 9917
rect 19429 9877 19441 9911
rect 19475 9908 19487 9911
rect 19610 9908 19616 9920
rect 19475 9880 19616 9908
rect 19475 9877 19487 9880
rect 19429 9871 19487 9877
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19889 9911 19947 9917
rect 19889 9908 19901 9911
rect 19760 9880 19901 9908
rect 19760 9868 19766 9880
rect 19889 9877 19901 9880
rect 19935 9877 19947 9911
rect 19889 9871 19947 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6052 9676 6745 9704
rect 6052 9664 6058 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 7101 9707 7159 9713
rect 7101 9673 7113 9707
rect 7147 9704 7159 9707
rect 7653 9707 7711 9713
rect 7653 9704 7665 9707
rect 7147 9676 7665 9704
rect 7147 9673 7159 9676
rect 7101 9667 7159 9673
rect 7653 9673 7665 9676
rect 7699 9673 7711 9707
rect 7653 9667 7711 9673
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 9916 9676 10241 9704
rect 9916 9664 9922 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 10229 9667 10287 9673
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10468 9676 10885 9704
rect 10468 9664 10474 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 13906 9704 13912 9716
rect 10873 9667 10931 9673
rect 13464 9676 13912 9704
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 5960 9608 6653 9636
rect 5960 9596 5966 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 8110 9636 8116 9648
rect 6641 9599 6699 9605
rect 7576 9608 8116 9636
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5031 9540 5641 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5629 9537 5641 9540
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5718 9528 5724 9540
rect 5776 9568 5782 9580
rect 5776 9540 7512 9568
rect 5776 9528 5782 9540
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 6270 9500 6276 9512
rect 5583 9472 6276 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 4617 9435 4675 9441
rect 4617 9401 4629 9435
rect 4663 9432 4675 9435
rect 4798 9432 4804 9444
rect 4663 9404 4804 9432
rect 4663 9401 4675 9404
rect 4617 9395 4675 9401
rect 4798 9392 4804 9404
rect 4856 9432 4862 9444
rect 5258 9432 5264 9444
rect 4856 9404 5264 9432
rect 4856 9392 4862 9404
rect 5258 9392 5264 9404
rect 5316 9432 5322 9444
rect 5552 9432 5580 9463
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9500 6607 9503
rect 7282 9500 7288 9512
rect 6595 9472 7288 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 5316 9404 5580 9432
rect 5316 9392 5322 9404
rect 5997 9367 6055 9373
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 7190 9364 7196 9376
rect 6043 9336 7196 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7484 9364 7512 9540
rect 7576 9509 7604 9608
rect 8110 9596 8116 9608
rect 8168 9596 8174 9648
rect 8662 9636 8668 9648
rect 8623 9608 8668 9636
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11609 9639 11667 9645
rect 11609 9636 11621 9639
rect 11296 9608 11621 9636
rect 11296 9596 11302 9608
rect 11609 9605 11621 9608
rect 11655 9636 11667 9639
rect 11698 9636 11704 9648
rect 11655 9608 11704 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 13464 9636 13492 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 14642 9664 14648 9716
rect 14700 9664 14706 9716
rect 14737 9707 14795 9713
rect 14737 9673 14749 9707
rect 14783 9704 14795 9707
rect 15102 9704 15108 9716
rect 14783 9676 15108 9704
rect 14783 9673 14795 9676
rect 14737 9667 14795 9673
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 16666 9704 16672 9716
rect 15620 9676 16672 9704
rect 15620 9664 15626 9676
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 17034 9704 17040 9716
rect 16995 9676 17040 9704
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18417 9707 18475 9713
rect 18417 9704 18429 9707
rect 18012 9676 18429 9704
rect 18012 9664 18018 9676
rect 18417 9673 18429 9676
rect 18463 9673 18475 9707
rect 18690 9704 18696 9716
rect 18651 9676 18696 9704
rect 18417 9667 18475 9673
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 19886 9704 19892 9716
rect 18892 9676 19748 9704
rect 19847 9676 19892 9704
rect 13630 9636 13636 9648
rect 12406 9608 13492 9636
rect 13591 9608 13636 9636
rect 7742 9568 7748 9580
rect 7703 9540 7748 9568
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 8803 9540 9076 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 8352 9472 8493 9500
rect 8352 9460 8358 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 8386 9432 8392 9444
rect 8159 9404 8392 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9048 9364 9076 9540
rect 9214 9528 9220 9580
rect 9272 9568 9278 9580
rect 12406 9568 12434 9608
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 14458 9636 14464 9648
rect 14148 9608 14464 9636
rect 14148 9596 14154 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 14660 9636 14688 9664
rect 18892 9636 18920 9676
rect 14660 9608 14780 9636
rect 9272 9540 12434 9568
rect 12529 9571 12587 9577
rect 9272 9528 9278 9540
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12575 9540 13216 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 10042 9500 10048 9512
rect 10003 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 12894 9500 12900 9512
rect 12851 9472 12900 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 10152 9432 10180 9463
rect 12158 9432 12164 9444
rect 9171 9404 10180 9432
rect 12119 9404 12164 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 7484 9336 9505 9364
rect 9493 9333 9505 9336
rect 9539 9364 9551 9367
rect 9674 9364 9680 9376
rect 9539 9336 9680 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 12636 9364 12664 9463
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13188 9441 13216 9540
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 13320 9540 13553 9568
rect 13320 9528 13326 9540
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 13541 9531 13599 9537
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 14366 9500 14372 9512
rect 13863 9472 14372 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 13173 9435 13231 9441
rect 13173 9401 13185 9435
rect 13219 9401 13231 9435
rect 13173 9395 13231 9401
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14752 9432 14780 9608
rect 17788 9608 18920 9636
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15654 9568 15660 9580
rect 14884 9540 15516 9568
rect 15615 9540 15660 9568
rect 14884 9528 14890 9540
rect 14918 9500 14924 9512
rect 14879 9472 14924 9500
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15160 9472 15393 9500
rect 15160 9460 15166 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15488 9500 15516 9540
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15948 9540 17540 9568
rect 15562 9500 15568 9512
rect 15488 9472 15568 9500
rect 15381 9463 15439 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 14826 9432 14832 9444
rect 14056 9404 14412 9432
rect 14752 9404 14832 9432
rect 14056 9392 14062 9404
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 12636 9336 14289 9364
rect 14277 9333 14289 9336
rect 14323 9333 14335 9367
rect 14384 9364 14412 9404
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 15948 9364 15976 9540
rect 16850 9500 16856 9512
rect 16811 9472 16856 9500
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17000 9472 17045 9500
rect 17000 9460 17006 9472
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 17126 9432 17132 9444
rect 16071 9404 17132 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 14384 9336 15976 9364
rect 14277 9327 14335 9333
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 16666 9364 16672 9376
rect 16172 9336 16672 9364
rect 16172 9324 16178 9336
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17092 9336 17417 9364
rect 17092 9324 17098 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17512 9364 17540 9540
rect 17788 9509 17816 9608
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 19720 9636 19748 9676
rect 19886 9664 19892 9676
rect 19944 9664 19950 9716
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 22094 9704 22100 9716
rect 21140 9676 22100 9704
rect 21140 9664 21146 9676
rect 22094 9664 22100 9676
rect 22152 9704 22158 9716
rect 22278 9704 22284 9716
rect 22152 9676 22284 9704
rect 22152 9664 22158 9676
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 20254 9636 20260 9648
rect 19024 9608 19472 9636
rect 19720 9608 20260 9636
rect 19024 9596 19030 9608
rect 19444 9577 19472 9608
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 20625 9639 20683 9645
rect 20625 9605 20637 9639
rect 20671 9636 20683 9639
rect 22554 9636 22560 9648
rect 20671 9608 22560 9636
rect 20671 9605 20683 9608
rect 20625 9599 20683 9605
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 17957 9572 18015 9577
rect 17880 9571 18015 9572
rect 17880 9544 17969 9571
rect 17773 9503 17831 9509
rect 17773 9469 17785 9503
rect 17819 9469 17831 9503
rect 17773 9463 17831 9469
rect 17880 9432 17908 9544
rect 17957 9537 17969 9544
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18095 9552 18368 9568
rect 18095 9540 18460 9552
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18340 9524 18460 9540
rect 18432 9444 18460 9524
rect 18524 9540 18889 9568
rect 17954 9432 17960 9444
rect 17880 9404 17960 9432
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 18414 9392 18420 9444
rect 18472 9392 18478 9444
rect 18524 9364 18552 9540
rect 18877 9537 18889 9540
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19702 9568 19708 9580
rect 19663 9540 19708 9568
rect 19429 9531 19487 9537
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 19812 9540 20545 9568
rect 19058 9392 19064 9444
rect 19116 9432 19122 9444
rect 19245 9435 19303 9441
rect 19245 9432 19257 9435
rect 19116 9404 19257 9432
rect 19116 9392 19122 9404
rect 19245 9401 19257 9404
rect 19291 9401 19303 9435
rect 19245 9395 19303 9401
rect 19702 9392 19708 9444
rect 19760 9432 19766 9444
rect 19812 9432 19840 9540
rect 20533 9537 20545 9540
rect 20579 9537 20591 9571
rect 21358 9568 21364 9580
rect 21319 9540 21364 9568
rect 20533 9531 20591 9537
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 20254 9460 20260 9512
rect 20312 9500 20318 9512
rect 20717 9503 20775 9509
rect 20717 9500 20729 9503
rect 20312 9472 20729 9500
rect 20312 9460 20318 9472
rect 20717 9469 20729 9472
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 21174 9432 21180 9444
rect 19760 9404 19840 9432
rect 21135 9404 21180 9432
rect 19760 9392 19766 9404
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 17512 9336 18552 9364
rect 17405 9327 17463 9333
rect 19150 9324 19156 9376
rect 19208 9364 19214 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19208 9336 20177 9364
rect 19208 9324 19214 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 5905 9163 5963 9169
rect 5905 9129 5917 9163
rect 5951 9160 5963 9163
rect 6638 9160 6644 9172
rect 5951 9132 6644 9160
rect 5951 9129 5963 9132
rect 5905 9123 5963 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7098 9120 7104 9172
rect 7156 9120 7162 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 9306 9160 9312 9172
rect 7340 9132 9312 9160
rect 7340 9120 7346 9132
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9160 10011 9163
rect 10502 9160 10508 9172
rect 9999 9132 10508 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10735 9132 11069 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 11057 9129 11069 9132
rect 11103 9160 11115 9163
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 11103 9132 11621 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11609 9129 11621 9132
rect 11655 9160 11667 9163
rect 11974 9160 11980 9172
rect 11655 9132 11980 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14366 9160 14372 9172
rect 14231 9132 14372 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14366 9120 14372 9132
rect 14424 9160 14430 9172
rect 14918 9160 14924 9172
rect 14424 9132 14924 9160
rect 14424 9120 14430 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15102 9160 15108 9172
rect 15063 9132 15108 9160
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 18414 9160 18420 9172
rect 15712 9132 18276 9160
rect 18375 9132 18420 9160
rect 15712 9120 15718 9132
rect 7116 9092 7144 9120
rect 6196 9064 7144 9092
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5994 9024 6000 9036
rect 5399 8996 6000 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5994 8984 6000 8996
rect 6052 9024 6058 9036
rect 6196 9024 6224 9064
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7432 9064 10548 9092
rect 7432 9052 7438 9064
rect 10520 9036 10548 9064
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 10652 9064 16896 9092
rect 10652 9052 10658 9064
rect 6052 8996 6224 9024
rect 6917 9027 6975 9033
rect 6052 8984 6058 8996
rect 6917 8993 6929 9027
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 4764 8860 5457 8888
rect 4764 8848 4770 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 6932 8888 6960 8987
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 7064 8996 7113 9024
rect 7064 8984 7070 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7834 9024 7840 9036
rect 7795 8996 7840 9024
rect 7101 8987 7159 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9024 9459 9027
rect 9582 9024 9588 9036
rect 9447 8996 9588 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10134 9024 10140 9036
rect 9916 8996 10140 9024
rect 9916 8984 9922 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 10836 8996 12449 9024
rect 10836 8984 10842 8996
rect 12437 8993 12449 8996
rect 12483 8993 12495 9027
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 12437 8987 12495 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16758 9024 16764 9036
rect 15979 8996 16764 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 7300 8928 9628 8956
rect 7300 8888 7328 8928
rect 9493 8891 9551 8897
rect 9493 8888 9505 8891
rect 6932 8860 7328 8888
rect 7576 8860 9505 8888
rect 5445 8851 5503 8857
rect 6270 8820 6276 8832
rect 6183 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8820 6334 8832
rect 7374 8820 7380 8832
rect 6328 8792 7380 8820
rect 6328 8780 6334 8792
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7576 8829 7604 8860
rect 9493 8857 9505 8860
rect 9539 8857 9551 8891
rect 9600 8888 9628 8928
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 16868 8965 16896 9064
rect 17402 9052 17408 9104
rect 17460 9092 17466 9104
rect 17460 9064 17908 9092
rect 17460 9052 17466 9064
rect 17770 9024 17776 9036
rect 16940 8996 17776 9024
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 9732 8928 12357 8956
rect 9732 8916 9738 8928
rect 12345 8925 12357 8928
rect 12391 8956 12403 8959
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 12391 8928 13645 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 13633 8925 13645 8928
rect 13679 8956 13691 8959
rect 16853 8959 16911 8965
rect 13679 8928 16160 8956
rect 13679 8925 13691 8928
rect 13633 8919 13691 8925
rect 10134 8888 10140 8900
rect 9600 8860 10140 8888
rect 9493 8851 9551 8857
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 11698 8888 11704 8900
rect 10244 8860 11704 8888
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8789 7619 8823
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 7561 8783 7619 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10244 8820 10272 8860
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12768 8860 14780 8888
rect 12768 8848 12774 8860
rect 10100 8792 10272 8820
rect 10321 8823 10379 8829
rect 10100 8780 10106 8792
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 10410 8820 10416 8832
rect 10367 8792 10416 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 11882 8820 11888 8832
rect 11843 8792 11888 8820
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12032 8792 12265 8820
rect 12032 8780 12038 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 12253 8783 12311 8789
rect 14553 8823 14611 8829
rect 14553 8789 14565 8823
rect 14599 8820 14611 8823
rect 14642 8820 14648 8832
rect 14599 8792 14648 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14752 8820 14780 8860
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 16025 8891 16083 8897
rect 16025 8888 16037 8891
rect 14976 8860 16037 8888
rect 14976 8848 14982 8860
rect 16025 8857 16037 8860
rect 16071 8857 16083 8891
rect 16132 8888 16160 8928
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 16940 8888 16968 8996
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 17880 9033 17908 9064
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 18138 9092 18144 9104
rect 18012 9064 18144 9092
rect 18012 9052 18018 9064
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 18248 9092 18276 9132
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 18840 9132 19840 9160
rect 18840 9120 18846 9132
rect 19426 9092 19432 9104
rect 18248 9064 19432 9092
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 9024 17923 9027
rect 18414 9024 18420 9036
rect 17911 8996 18420 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 19702 9024 19708 9036
rect 19663 8996 19708 9024
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 19812 9024 19840 9132
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20404 9132 20453 9160
rect 20404 9120 20410 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 20165 9095 20223 9101
rect 20165 9061 20177 9095
rect 20211 9092 20223 9095
rect 20714 9092 20720 9104
rect 20211 9064 20720 9092
rect 20211 9061 20223 9064
rect 20165 9055 20223 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 20993 9027 21051 9033
rect 20993 9024 21005 9027
rect 19812 8996 21005 9024
rect 20993 8993 21005 8996
rect 21039 8993 21051 9027
rect 20993 8987 21051 8993
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 17460 8928 18705 8956
rect 17460 8916 17466 8928
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 19981 8959 20039 8965
rect 19981 8956 19993 8959
rect 19668 8928 19993 8956
rect 19668 8916 19674 8928
rect 19981 8925 19993 8928
rect 20027 8925 20039 8959
rect 19981 8919 20039 8925
rect 16132 8860 16968 8888
rect 17052 8860 20576 8888
rect 16025 8851 16083 8857
rect 16114 8820 16120 8832
rect 14752 8792 16120 8820
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16942 8820 16948 8832
rect 16531 8792 16948 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17052 8829 17080 8860
rect 17037 8823 17095 8829
rect 17037 8789 17049 8823
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 17494 8820 17500 8832
rect 17451 8792 17500 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18230 8820 18236 8832
rect 18095 8792 18236 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8820 18935 8823
rect 18966 8820 18972 8832
rect 18923 8792 18972 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 20548 8820 20576 8860
rect 20622 8848 20628 8900
rect 20680 8888 20686 8900
rect 20901 8891 20959 8897
rect 20901 8888 20913 8891
rect 20680 8860 20913 8888
rect 20680 8848 20686 8860
rect 20901 8857 20913 8860
rect 20947 8857 20959 8891
rect 20901 8851 20959 8857
rect 20714 8820 20720 8832
rect 20548 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 20809 8823 20867 8829
rect 20809 8789 20821 8823
rect 20855 8820 20867 8823
rect 20990 8820 20996 8832
rect 20855 8792 20996 8820
rect 20855 8789 20867 8792
rect 20809 8783 20867 8789
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 7282 8616 7288 8628
rect 7243 8588 7288 8616
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 9490 8616 9496 8628
rect 7984 8588 9496 8616
rect 7984 8576 7990 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10137 8619 10195 8625
rect 10137 8616 10149 8619
rect 9640 8588 10149 8616
rect 9640 8576 9646 8588
rect 10137 8585 10149 8588
rect 10183 8585 10195 8619
rect 10137 8579 10195 8585
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 11609 8619 11667 8625
rect 10468 8588 11008 8616
rect 10468 8576 10474 8588
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 8352 8520 10517 8548
rect 8352 8508 8358 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 10505 8511 10563 8517
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 9493 8483 9551 8489
rect 8260 8452 9444 8480
rect 8260 8440 8266 8452
rect 5258 8412 5264 8424
rect 5219 8384 5264 8412
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5592 8384 6377 8412
rect 5592 8372 5598 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 6365 8375 6423 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7926 8412 7932 8424
rect 7607 8384 7932 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 9122 8372 9128 8424
rect 9180 8372 9186 8424
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 6696 8316 6929 8344
rect 6696 8304 6702 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 9140 8344 9168 8372
rect 9416 8344 9444 8452
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9539 8452 10088 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9582 8412 9588 8424
rect 9543 8384 9588 8412
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 9732 8384 9777 8412
rect 9732 8372 9738 8384
rect 10060 8356 10088 8452
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10980 8480 11008 8588
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 11698 8616 11704 8628
rect 11655 8588 11704 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12250 8616 12256 8628
rect 12211 8588 12256 8616
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12713 8619 12771 8625
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 13722 8616 13728 8628
rect 12759 8588 13728 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 16298 8616 16304 8628
rect 16259 8588 16304 8616
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17402 8616 17408 8628
rect 17092 8588 17137 8616
rect 17363 8588 17408 8616
rect 17092 8576 17098 8588
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8585 17923 8619
rect 18138 8616 18144 8628
rect 18099 8588 18144 8616
rect 17865 8579 17923 8585
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 17604 8548 17632 8576
rect 14516 8520 17632 8548
rect 17880 8548 17908 8579
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 20622 8616 20628 8628
rect 18432 8588 20392 8616
rect 20583 8588 20628 8616
rect 18432 8548 18460 8588
rect 20254 8548 20260 8560
rect 17880 8520 18460 8548
rect 18524 8520 20260 8548
rect 14516 8508 14522 8520
rect 12986 8480 12992 8492
rect 10284 8452 10732 8480
rect 10980 8452 12992 8480
rect 10284 8440 10290 8452
rect 10594 8412 10600 8424
rect 10555 8384 10600 8412
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10704 8421 10732 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13127 8452 13645 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 11054 8372 11060 8424
rect 11112 8412 11118 8424
rect 13096 8412 13124 8443
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 13780 8452 15025 8480
rect 13780 8440 13786 8452
rect 15013 8449 15025 8452
rect 15059 8480 15071 8483
rect 15102 8480 15108 8492
rect 15059 8452 15108 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 17586 8480 17592 8492
rect 16163 8452 17592 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 11112 8384 13124 8412
rect 13541 8415 13599 8421
rect 11112 8372 11118 8384
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 14274 8412 14280 8424
rect 13587 8384 14280 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 14458 8412 14464 8424
rect 14419 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 14976 8384 15577 8412
rect 14976 8372 14982 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17218 8412 17224 8424
rect 16899 8384 17224 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 17696 8412 17724 8443
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18524 8489 18552 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 20364 8548 20392 8588
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 21082 8548 21088 8560
rect 20364 8520 21088 8548
rect 21082 8508 21088 8520
rect 21140 8508 21146 8560
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18012 8452 18521 8480
rect 18012 8440 18018 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 19058 8480 19064 8492
rect 18647 8452 19064 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8449 19211 8483
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19153 8443 19211 8449
rect 19260 8452 19901 8480
rect 17460 8384 17724 8412
rect 17460 8372 17466 8384
rect 18414 8372 18420 8424
rect 18472 8412 18478 8424
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 18472 8384 18705 8412
rect 18472 8372 18478 8384
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 9140 8316 9352 8344
rect 9416 8316 9996 8344
rect 6917 8307 6975 8313
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 8021 8279 8079 8285
rect 8021 8276 8033 8279
rect 7432 8248 8033 8276
rect 7432 8236 7438 8248
rect 8021 8245 8033 8248
rect 8067 8276 8079 8279
rect 8202 8276 8208 8288
rect 8067 8248 8208 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 9122 8276 9128 8288
rect 9083 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9324 8276 9352 8316
rect 9490 8276 9496 8288
rect 9324 8248 9496 8276
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9968 8276 9996 8316
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 10100 8316 11989 8344
rect 10100 8304 10106 8316
rect 11977 8313 11989 8316
rect 12023 8344 12035 8347
rect 12434 8344 12440 8356
rect 12023 8316 12440 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 19168 8344 19196 8443
rect 15068 8316 19196 8344
rect 15068 8304 15074 8316
rect 11330 8276 11336 8288
rect 9968 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11882 8276 11888 8288
rect 11480 8248 11888 8276
rect 11480 8236 11486 8248
rect 11882 8236 11888 8248
rect 11940 8276 11946 8288
rect 13722 8276 13728 8288
rect 11940 8248 13728 8276
rect 11940 8236 11946 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14366 8276 14372 8288
rect 14139 8248 14372 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 19260 8276 19288 8452
rect 19889 8449 19901 8452
rect 19935 8480 19947 8483
rect 19978 8480 19984 8492
rect 19935 8452 19984 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20346 8480 20352 8492
rect 20307 8452 20352 8480
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21450 8412 21456 8424
rect 21315 8384 21456 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 19337 8347 19395 8353
rect 19337 8313 19349 8347
rect 19383 8344 19395 8347
rect 19794 8344 19800 8356
rect 19383 8316 19800 8344
rect 19383 8313 19395 8316
rect 19337 8307 19395 8313
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 20165 8347 20223 8353
rect 20165 8313 20177 8347
rect 20211 8344 20223 8347
rect 22646 8344 22652 8356
rect 20211 8316 22652 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 22646 8304 22652 8316
rect 22704 8304 22710 8356
rect 16172 8248 19288 8276
rect 16172 8236 16178 8248
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19484 8248 19717 8276
rect 19484 8236 19490 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6788 8044 6837 8072
rect 6788 8032 6794 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 7800 8044 8953 8072
rect 7800 8032 7806 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 10042 8072 10048 8084
rect 8941 8035 8999 8041
rect 9048 8044 9904 8072
rect 10003 8044 10048 8072
rect 4982 7964 4988 8016
rect 5040 8004 5046 8016
rect 7926 8004 7932 8016
rect 5040 7976 7932 8004
rect 5040 7964 5046 7976
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 8202 7964 8208 8016
rect 8260 8004 8266 8016
rect 9048 8004 9076 8044
rect 8260 7976 9076 8004
rect 8260 7964 8266 7976
rect 9306 7964 9312 8016
rect 9364 8004 9370 8016
rect 9876 8004 9904 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10376 8044 10885 8072
rect 10376 8032 10382 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12676 8044 12909 8072
rect 12676 8032 12682 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13044 8044 13277 8072
rect 13044 8032 13050 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 14550 8072 14556 8084
rect 13265 8035 13323 8041
rect 13464 8044 14556 8072
rect 11422 8004 11428 8016
rect 9364 7976 9536 8004
rect 9876 7976 11428 8004
rect 9364 7964 9370 7976
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5350 7936 5356 7948
rect 5307 7908 5356 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6052 7908 6193 7936
rect 6052 7896 6058 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 6638 7936 6644 7948
rect 6411 7908 6644 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9508 7945 9536 7976
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 13464 8004 13492 8044
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 15930 8072 15936 8084
rect 15804 8044 15936 8072
rect 15804 8032 15810 8044
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 17644 8044 18061 8072
rect 17644 8032 17650 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 19886 8072 19892 8084
rect 19847 8044 19892 8072
rect 18049 8035 18107 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20349 8075 20407 8081
rect 20349 8072 20361 8075
rect 20312 8044 20361 8072
rect 20312 8032 20318 8044
rect 20349 8041 20361 8044
rect 20395 8041 20407 8075
rect 21266 8072 21272 8084
rect 21227 8044 21272 8072
rect 20349 8035 20407 8041
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 11532 7976 13492 8004
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9180 7908 9413 7936
rect 9180 7896 9186 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 11330 7936 11336 7948
rect 11291 7908 11336 7936
rect 9493 7899 9551 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11532 7945 11560 7976
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 18414 8004 18420 8016
rect 13780 7976 18420 8004
rect 13780 7964 13786 7976
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 20993 8007 21051 8013
rect 18564 7976 20576 8004
rect 18564 7964 18570 7976
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12618 7936 12624 7948
rect 12391 7908 12624 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 14274 7936 14280 7948
rect 14235 7908 14280 7936
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 16114 7936 16120 7948
rect 14384 7908 16120 7936
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5534 7868 5540 7880
rect 5491 7840 5540 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 11054 7868 11060 7880
rect 8619 7840 11060 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 11348 7868 11376 7896
rect 11974 7868 11980 7880
rect 11348 7840 11980 7868
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12492 7840 12541 7868
rect 12492 7828 12498 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 14384 7868 14412 7908
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 17218 7936 17224 7948
rect 16264 7908 17224 7936
rect 16264 7896 16270 7908
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 18690 7936 18696 7948
rect 18651 7908 18696 7936
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 12529 7831 12587 7837
rect 14200 7840 14412 7868
rect 14476 7840 17049 7868
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 5828 7772 9321 7800
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 4709 7735 4767 7741
rect 4709 7732 4721 7735
rect 4672 7704 4721 7732
rect 4672 7692 4678 7704
rect 4709 7701 4721 7704
rect 4755 7732 4767 7735
rect 5166 7732 5172 7744
rect 4755 7704 5172 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 5166 7692 5172 7704
rect 5224 7732 5230 7744
rect 5828 7741 5856 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 14200 7800 14228 7840
rect 10643 7772 14228 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 14274 7760 14280 7812
rect 14332 7800 14338 7812
rect 14476 7800 14504 7840
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 20070 7868 20076 7880
rect 20031 7840 20076 7868
rect 17037 7831 17095 7837
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20548 7877 20576 7976
rect 20993 7973 21005 8007
rect 21039 8004 21051 8007
rect 21634 8004 21640 8016
rect 21039 7976 21640 8004
rect 21039 7973 21051 7976
rect 20993 7967 21051 7973
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 20772 7840 20821 7868
rect 20772 7828 20778 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 14332 7772 14504 7800
rect 14332 7760 14338 7772
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 14608 7772 14872 7800
rect 14608 7760 14614 7772
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 5224 7704 5365 7732
rect 5224 7692 5230 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5960 7704 6469 7732
rect 5960 7692 5966 7704
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 6457 7695 6515 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 11020 7704 11253 7732
rect 11020 7692 11026 7704
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 11241 7695 11299 7701
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 11756 7704 12449 7732
rect 11756 7692 11762 7704
rect 12437 7701 12449 7704
rect 12483 7732 12495 7735
rect 12710 7732 12716 7744
rect 12483 7704 12716 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7732 13694 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 13688 7704 14381 7732
rect 13688 7692 13694 7704
rect 14369 7701 14381 7704
rect 14415 7701 14427 7735
rect 14369 7695 14427 7701
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 14844 7741 14872 7772
rect 15286 7760 15292 7812
rect 15344 7800 15350 7812
rect 16945 7803 17003 7809
rect 15344 7772 16712 7800
rect 15344 7760 15350 7772
rect 14829 7735 14887 7741
rect 14516 7704 14561 7732
rect 14516 7692 14522 7704
rect 14829 7701 14841 7735
rect 14875 7701 14887 7735
rect 15654 7732 15660 7744
rect 15615 7704 15660 7732
rect 14829 7695 14887 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 16022 7732 16028 7744
rect 15983 7704 16028 7732
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 16172 7704 16589 7732
rect 16172 7692 16178 7704
rect 16577 7701 16589 7704
rect 16623 7701 16635 7735
rect 16684 7732 16712 7772
rect 16945 7769 16957 7803
rect 16991 7800 17003 7803
rect 17126 7800 17132 7812
rect 16991 7772 17132 7800
rect 16991 7769 17003 7772
rect 16945 7763 17003 7769
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 18230 7760 18236 7812
rect 18288 7800 18294 7812
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 18288 7772 19257 7800
rect 18288 7760 18294 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 17402 7732 17408 7744
rect 16684 7704 17408 7732
rect 16577 7695 16635 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17586 7732 17592 7744
rect 17547 7704 17592 7732
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 18564 7704 18609 7732
rect 18564 7692 18570 7704
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 22462 7732 22468 7744
rect 18840 7704 22468 7732
rect 18840 7692 18846 7704
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 5902 7528 5908 7540
rect 5675 7500 5908 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 6733 7531 6791 7537
rect 6733 7497 6745 7531
rect 6779 7528 6791 7531
rect 7098 7528 7104 7540
rect 6779 7500 7104 7528
rect 6779 7497 6791 7500
rect 6733 7491 6791 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 8018 7528 8024 7540
rect 7979 7500 8024 7528
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 9214 7528 9220 7540
rect 8435 7500 9220 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 10594 7528 10600 7540
rect 9815 7500 10600 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 10744 7500 11529 7528
rect 10744 7488 10750 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11940 7500 11989 7528
rect 11940 7488 11946 7500
rect 11977 7497 11989 7500
rect 12023 7528 12035 7531
rect 12342 7528 12348 7540
rect 12023 7500 12348 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 13630 7528 13636 7540
rect 13504 7500 13636 7528
rect 13504 7488 13510 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13872 7500 13921 7528
rect 13872 7488 13878 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 14550 7528 14556 7540
rect 14511 7500 14556 7528
rect 13909 7491 13967 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15010 7528 15016 7540
rect 14967 7500 15016 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 16114 7528 16120 7540
rect 15703 7500 16120 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16942 7528 16948 7540
rect 16347 7500 16948 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17037 7531 17095 7537
rect 17037 7497 17049 7531
rect 17083 7528 17095 7531
rect 17586 7528 17592 7540
rect 17083 7500 17592 7528
rect 17083 7497 17095 7500
rect 17037 7491 17095 7497
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18472 7500 18613 7528
rect 18472 7488 18478 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7497 18935 7531
rect 18877 7491 18935 7497
rect 5997 7463 6055 7469
rect 5997 7429 6009 7463
rect 6043 7460 6055 7463
rect 6086 7460 6092 7472
rect 6043 7432 6092 7460
rect 6043 7429 6055 7432
rect 5997 7423 6055 7429
rect 6086 7420 6092 7432
rect 6144 7460 6150 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6144 7432 6653 7460
rect 6144 7420 6150 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 6822 7460 6828 7472
rect 6687 7432 6828 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7460 9367 7463
rect 9582 7460 9588 7472
rect 9355 7432 9588 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 9582 7420 9588 7432
rect 9640 7460 9646 7472
rect 11698 7460 11704 7472
rect 9640 7432 11704 7460
rect 9640 7420 9646 7432
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 14366 7420 14372 7472
rect 14424 7460 14430 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 14424 7432 14473 7460
rect 14424 7420 14430 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 15160 7432 16160 7460
rect 15160 7420 15166 7432
rect 16132 7404 16160 7432
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18141 7463 18199 7469
rect 18141 7460 18153 7463
rect 18104 7432 18153 7460
rect 18104 7420 18110 7432
rect 18141 7429 18153 7432
rect 18187 7429 18199 7463
rect 18141 7423 18199 7429
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 10042 7392 10048 7404
rect 9447 7364 10048 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10778 7392 10784 7404
rect 10284 7364 10784 7392
rect 10284 7352 10290 7364
rect 10778 7352 10784 7364
rect 10836 7392 10842 7404
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 10836 7364 11069 7392
rect 10836 7352 10842 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11882 7392 11888 7404
rect 11843 7364 11888 7392
rect 11057 7355 11115 7361
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 12768 7364 13553 7392
rect 12768 7352 12774 7364
rect 13541 7361 13553 7364
rect 13587 7361 13599 7395
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 13541 7355 13599 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 17678 7392 17684 7404
rect 16776 7364 17684 7392
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7188 4586 7200
rect 4890 7188 4896 7200
rect 4580 7160 4896 7188
rect 4580 7148 4586 7160
rect 4890 7148 4896 7160
rect 4948 7188 4954 7200
rect 5184 7188 5212 7287
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 5500 7296 6561 7324
rect 5500 7284 5506 7296
rect 6549 7293 6561 7296
rect 6595 7324 6607 7327
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 6595 7296 9137 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 11514 7324 11520 7336
rect 9916 7296 11520 7324
rect 9916 7284 9922 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12124 7296 12169 7324
rect 12268 7296 13216 7324
rect 12124 7284 12130 7296
rect 7101 7259 7159 7265
rect 7101 7225 7113 7259
rect 7147 7256 7159 7259
rect 8294 7256 8300 7268
rect 7147 7228 8300 7256
rect 7147 7225 7159 7228
rect 7101 7219 7159 7225
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7256 8815 7259
rect 12268 7256 12296 7296
rect 8803 7228 12296 7256
rect 8803 7225 8815 7228
rect 8757 7219 8815 7225
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 12400 7228 12541 7256
rect 12400 7216 12406 7228
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 13188 7256 13216 7296
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13446 7324 13452 7336
rect 13320 7296 13365 7324
rect 13407 7296 13452 7324
rect 13320 7284 13326 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 15194 7324 15200 7336
rect 14415 7296 15200 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 15930 7324 15936 7336
rect 15887 7296 15936 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16776 7333 16804 7364
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 18782 7392 18788 7404
rect 18064 7364 18788 7392
rect 18064 7336 18092 7364
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7293 16819 7327
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16761 7287 16819 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 18046 7324 18052 7336
rect 17959 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 18892 7324 18920 7491
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 19576 7500 19809 7528
rect 19576 7488 19582 7500
rect 19797 7497 19809 7500
rect 19843 7497 19855 7531
rect 19797 7491 19855 7497
rect 20257 7531 20315 7537
rect 20257 7497 20269 7531
rect 20303 7528 20315 7531
rect 20438 7528 20444 7540
rect 20303 7500 20444 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20898 7528 20904 7540
rect 20859 7500 20904 7528
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19024 7432 20760 7460
rect 19024 7420 19030 7432
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19334 7392 19340 7404
rect 19295 7364 19340 7392
rect 19061 7355 19119 7361
rect 18656 7296 18920 7324
rect 18656 7284 18662 7296
rect 17405 7259 17463 7265
rect 13188 7228 17356 7256
rect 12529 7219 12587 7225
rect 4948 7160 5212 7188
rect 4948 7148 4954 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10410 7188 10416 7200
rect 9824 7160 10416 7188
rect 9824 7148 9830 7160
rect 10410 7148 10416 7160
rect 10468 7188 10474 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10468 7160 10701 7188
rect 10468 7148 10474 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12250 7188 12256 7200
rect 12032 7160 12256 7188
rect 12032 7148 12038 7160
rect 12250 7148 12256 7160
rect 12308 7188 12314 7200
rect 12986 7188 12992 7200
rect 12308 7160 12992 7188
rect 12308 7148 12314 7160
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 14608 7160 15209 7188
rect 14608 7148 14614 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 17328 7188 17356 7228
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 19076 7256 19104 7355
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 19978 7392 19984 7404
rect 19444 7364 19984 7392
rect 17451 7228 19104 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 19444 7188 19472 7364
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20732 7401 20760 7432
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 22278 7392 22284 7404
rect 21407 7364 22284 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 20456 7324 20484 7355
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 19536 7296 20484 7324
rect 19536 7265 19564 7296
rect 19521 7259 19579 7265
rect 19521 7225 19533 7259
rect 19567 7225 19579 7259
rect 19521 7219 19579 7225
rect 17328 7160 19472 7188
rect 15197 7151 15255 7157
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 21177 7191 21235 7197
rect 21177 7188 21189 7191
rect 20772 7160 21189 7188
rect 20772 7148 20778 7160
rect 21177 7157 21189 7160
rect 21223 7157 21235 7191
rect 21177 7151 21235 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 10778 6984 10784 6996
rect 6880 6956 10784 6984
rect 6880 6944 6886 6956
rect 10778 6944 10784 6956
rect 10836 6984 10842 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 10836 6956 11437 6984
rect 10836 6944 10842 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 11425 6947 11483 6953
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 13446 6984 13452 6996
rect 11572 6956 13452 6984
rect 11572 6944 11578 6956
rect 13446 6944 13452 6956
rect 13504 6984 13510 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13504 6956 13645 6984
rect 13504 6944 13510 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14366 6984 14372 6996
rect 13872 6956 14372 6984
rect 13872 6944 13878 6956
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 15562 6984 15568 6996
rect 15523 6956 15568 6984
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17313 6987 17371 6993
rect 17313 6984 17325 6987
rect 17000 6956 17325 6984
rect 17000 6944 17006 6956
rect 17313 6953 17325 6956
rect 17359 6953 17371 6987
rect 17313 6947 17371 6953
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17460 6956 18000 6984
rect 17460 6944 17466 6956
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6916 10471 6919
rect 10502 6916 10508 6928
rect 10459 6888 10508 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10686 6916 10692 6928
rect 10647 6888 10692 6916
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 12342 6916 12348 6928
rect 11112 6888 12348 6916
rect 11112 6876 11118 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 12894 6916 12900 6928
rect 12584 6888 12900 6916
rect 12584 6876 12590 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 17972 6916 18000 6956
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18564 6956 18613 6984
rect 18564 6944 18570 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18601 6947 18659 6953
rect 20441 6987 20499 6993
rect 20441 6953 20453 6987
rect 20487 6984 20499 6987
rect 20487 6956 20852 6984
rect 20487 6953 20499 6956
rect 20441 6947 20499 6953
rect 19150 6916 19156 6928
rect 13044 6888 17908 6916
rect 17972 6888 19156 6916
rect 13044 6876 13050 6888
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8202 6848 8208 6860
rect 8163 6820 8208 6848
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 10962 6848 10968 6860
rect 8312 6820 10968 6848
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 8312 6780 8340 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 12023 6820 14749 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 14737 6817 14749 6820
rect 14783 6848 14795 6851
rect 14826 6848 14832 6860
rect 14783 6820 14832 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15194 6848 15200 6860
rect 15155 6820 15200 6848
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 15304 6820 16160 6848
rect 9122 6780 9128 6792
rect 6880 6752 8340 6780
rect 9083 6752 9128 6780
rect 6880 6740 6886 6752
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9490 6780 9496 6792
rect 9451 6752 9496 6780
rect 9490 6740 9496 6752
rect 9548 6780 9554 6792
rect 9858 6780 9864 6792
rect 9548 6752 9864 6780
rect 9548 6740 9554 6752
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 13722 6780 13728 6792
rect 10428 6752 13728 6780
rect 8573 6715 8631 6721
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 10428 6712 10456 6752
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 15304 6780 15332 6820
rect 14016 6752 15332 6780
rect 15933 6783 15991 6789
rect 8619 6684 10456 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11057 6715 11115 6721
rect 11057 6712 11069 6715
rect 10928 6684 11069 6712
rect 10928 6672 10934 6684
rect 11057 6681 11069 6684
rect 11103 6712 11115 6715
rect 11974 6712 11980 6724
rect 11103 6684 11980 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11974 6672 11980 6684
rect 12032 6672 12038 6724
rect 12069 6715 12127 6721
rect 12069 6681 12081 6715
rect 12115 6712 12127 6715
rect 12618 6712 12624 6724
rect 12115 6684 12624 6712
rect 12115 6681 12127 6684
rect 12069 6675 12127 6681
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 14016 6712 14044 6752
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16132 6780 16160 6820
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16761 6851 16819 6857
rect 16264 6820 16309 6848
rect 16264 6808 16270 6820
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17310 6848 17316 6860
rect 16807 6820 17316 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16132 6752 16865 6780
rect 16853 6749 16865 6752
rect 16899 6780 16911 6783
rect 17770 6780 17776 6792
rect 16899 6752 17776 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 17880 6780 17908 6888
rect 19150 6876 19156 6888
rect 19208 6876 19214 6928
rect 20717 6919 20775 6925
rect 20717 6885 20729 6919
rect 20763 6885 20775 6919
rect 20717 6879 20775 6885
rect 18046 6848 18052 6860
rect 18007 6820 18052 6848
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 20732 6848 20760 6879
rect 18892 6820 20760 6848
rect 20824 6848 20852 6956
rect 20990 6848 20996 6860
rect 20824 6820 20996 6848
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17880 6752 18245 6780
rect 18233 6749 18245 6752
rect 18279 6780 18291 6783
rect 18782 6780 18788 6792
rect 18279 6752 18788 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 12952 6684 14044 6712
rect 14461 6715 14519 6721
rect 12952 6672 12958 6684
rect 14461 6681 14473 6715
rect 14507 6712 14519 6715
rect 15010 6712 15016 6724
rect 14507 6684 15016 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 15010 6672 15016 6684
rect 15068 6712 15074 6724
rect 18892 6712 18920 6820
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19794 6780 19800 6792
rect 19755 6752 19800 6780
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 20254 6780 20260 6792
rect 20215 6752 20260 6780
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20364 6752 20576 6780
rect 20364 6712 20392 6752
rect 15068 6684 18920 6712
rect 18984 6684 20392 6712
rect 15068 6672 15074 6684
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 10836 6616 12173 6644
rect 10836 6604 10842 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12161 6607 12219 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12986 6644 12992 6656
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13446 6644 13452 6656
rect 13403 6616 13452 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 14826 6644 14832 6656
rect 14599 6616 14832 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 16025 6647 16083 6653
rect 16025 6644 16037 6647
rect 15896 6616 16037 6644
rect 15896 6604 15902 6616
rect 16025 6613 16037 6616
rect 16071 6613 16083 6647
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16025 6607 16083 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18141 6647 18199 6653
rect 18141 6644 18153 6647
rect 18104 6616 18153 6644
rect 18104 6604 18110 6616
rect 18141 6613 18153 6616
rect 18187 6613 18199 6647
rect 18141 6607 18199 6613
rect 18230 6604 18236 6656
rect 18288 6644 18294 6656
rect 18984 6644 19012 6684
rect 18288 6616 19012 6644
rect 18288 6604 18294 6616
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 19337 6647 19395 6653
rect 19337 6644 19349 6647
rect 19116 6616 19349 6644
rect 19116 6604 19122 6616
rect 19337 6613 19349 6616
rect 19383 6613 19395 6647
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19337 6607 19395 6613
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20548 6644 20576 6752
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20864 6752 20913 6780
rect 20864 6740 20870 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 21358 6780 21364 6792
rect 21319 6752 21364 6780
rect 20901 6743 20959 6749
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 20548 6616 21189 6644
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 7984 6412 8401 6440
rect 7984 6400 7990 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 8389 6403 8447 6409
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9539 6412 10057 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12032 6412 12173 6440
rect 12032 6400 12038 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 13538 6400 13544 6452
rect 13596 6440 13602 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13596 6412 14473 6440
rect 13596 6400 13602 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 14599 6412 16681 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17586 6440 17592 6452
rect 17083 6412 17592 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 18012 6412 18061 6440
rect 18012 6400 18018 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 19058 6440 19064 6452
rect 18187 6412 19064 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19889 6443 19947 6449
rect 19889 6409 19901 6443
rect 19935 6440 19947 6443
rect 20346 6440 20352 6452
rect 19935 6412 20352 6440
rect 19935 6409 19947 6412
rect 19889 6403 19947 6409
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21140 6412 21185 6440
rect 21140 6400 21146 6412
rect 9033 6375 9091 6381
rect 9033 6341 9045 6375
rect 9079 6372 9091 6375
rect 10594 6372 10600 6384
rect 9079 6344 10600 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 11072 6344 13400 6372
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6304 1458 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1452 6276 1869 6304
rect 1452 6264 1458 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 9122 6304 9128 6316
rect 9083 6276 9128 6304
rect 1857 6267 1915 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 10134 6304 10140 6316
rect 10095 6276 10140 6304
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 8202 6236 8208 6248
rect 7708 6208 8208 6236
rect 7708 6196 7714 6208
rect 8202 6196 8208 6208
rect 8260 6236 8266 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8260 6208 8861 6236
rect 8260 6196 8266 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 9950 6236 9956 6248
rect 9911 6208 9956 6236
rect 8849 6199 8907 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 1578 6168 1584 6180
rect 1539 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 8113 6171 8171 6177
rect 8113 6137 8125 6171
rect 8159 6168 8171 6171
rect 11072 6168 11100 6344
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 12158 6304 12164 6316
rect 11195 6276 12164 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11992 6245 12020 6276
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13372 6304 13400 6344
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 15102 6372 15108 6384
rect 13504 6344 15108 6372
rect 13504 6332 13510 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 19242 6372 19248 6384
rect 15396 6344 19248 6372
rect 15396 6304 15424 6344
rect 19242 6332 19248 6344
rect 19300 6372 19306 6384
rect 19300 6344 19472 6372
rect 19300 6332 19306 6344
rect 13372 6276 15424 6304
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15930 6304 15936 6316
rect 15519 6276 15936 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16298 6304 16304 6316
rect 16211 6276 16304 6304
rect 16298 6264 16304 6276
rect 16356 6304 16362 6316
rect 18414 6304 18420 6316
rect 16356 6276 18420 6304
rect 16356 6264 16362 6276
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18966 6304 18972 6316
rect 18927 6276 18972 6304
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19444 6313 19472 6344
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19518 6264 19524 6316
rect 19576 6304 19582 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19576 6276 19717 6304
rect 19576 6264 19582 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6304 20407 6307
rect 20438 6304 20444 6316
rect 20395 6276 20444 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 12084 6168 12112 6199
rect 12342 6168 12348 6180
rect 8159 6140 11100 6168
rect 11992 6140 12348 6168
rect 8159 6137 8171 6140
rect 8113 6131 8171 6137
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11992 6100 12020 6140
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12529 6171 12587 6177
rect 12529 6137 12541 6171
rect 12575 6168 12587 6171
rect 12618 6168 12624 6180
rect 12575 6140 12624 6168
rect 12575 6137 12587 6140
rect 12529 6131 12587 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12802 6168 12808 6180
rect 12763 6140 12808 6168
rect 12802 6128 12808 6140
rect 12860 6128 12866 6180
rect 10744 6072 12020 6100
rect 10744 6060 10750 6072
rect 12894 6060 12900 6112
rect 12952 6100 12958 6112
rect 13280 6100 13308 6199
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13412 6208 13457 6236
rect 13412 6196 13418 6208
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 14090 6236 14096 6248
rect 13596 6208 14096 6236
rect 13596 6196 13602 6208
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14642 6236 14648 6248
rect 14603 6208 14648 6236
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 15194 6236 15200 6248
rect 15155 6208 15200 6236
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 16942 6236 16948 6248
rect 15427 6208 16948 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 17402 6236 17408 6248
rect 17359 6208 17408 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 14826 6128 14832 6180
rect 14884 6168 14890 6180
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 14884 6140 16129 6168
rect 14884 6128 14890 6140
rect 16117 6137 16129 6140
rect 16163 6137 16175 6171
rect 17144 6168 17172 6199
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18230 6236 18236 6248
rect 18191 6208 18236 6236
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18340 6208 19334 6236
rect 16117 6131 16175 6137
rect 16408 6140 17172 6168
rect 12952 6072 13308 6100
rect 12952 6060 12958 6072
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 13872 6072 14105 6100
rect 13872 6060 13878 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 14093 6063 14151 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 16408 6100 16436 6140
rect 17218 6128 17224 6180
rect 17276 6168 17282 6180
rect 18340 6168 18368 6208
rect 17276 6140 18368 6168
rect 19306 6168 19334 6208
rect 21082 6196 21088 6248
rect 21140 6236 21146 6248
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 21140 6208 21189 6236
rect 21140 6196 21146 6208
rect 21177 6205 21189 6208
rect 21223 6236 21235 6239
rect 22738 6236 22744 6248
rect 21223 6208 22744 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 22738 6196 22744 6208
rect 22796 6196 22802 6248
rect 20165 6171 20223 6177
rect 20165 6168 20177 6171
rect 19306 6140 20177 6168
rect 17276 6128 17282 6140
rect 20165 6137 20177 6140
rect 20211 6137 20223 6171
rect 20165 6131 20223 6137
rect 16080 6072 16436 6100
rect 16080 6060 16086 6072
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 16540 6072 17693 6100
rect 16540 6060 16546 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 18785 6103 18843 6109
rect 18785 6100 18797 6103
rect 18656 6072 18797 6100
rect 18656 6060 18662 6072
rect 18785 6069 18797 6072
rect 18831 6069 18843 6103
rect 18785 6063 18843 6069
rect 18966 6060 18972 6112
rect 19024 6100 19030 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 19024 6072 19257 6100
rect 19024 6060 19030 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 20622 6100 20628 6112
rect 20583 6072 20628 6100
rect 19245 6063 19303 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8720 5868 8953 5896
rect 8720 5856 8726 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 10045 5899 10103 5905
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 10134 5896 10140 5908
rect 10091 5868 10140 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 10686 5896 10692 5908
rect 10459 5868 10692 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 10686 5856 10692 5868
rect 10744 5896 10750 5908
rect 11238 5896 11244 5908
rect 10744 5868 11244 5896
rect 10744 5856 10750 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11756 5868 11897 5896
rect 11756 5856 11762 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 15930 5896 15936 5908
rect 12032 5868 13400 5896
rect 15891 5868 15936 5896
rect 12032 5856 12038 5868
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 12802 5828 12808 5840
rect 4120 5800 10824 5828
rect 4120 5788 4126 5800
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 10796 5769 10824 5800
rect 11072 5800 12808 5828
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 8260 5732 9413 5760
rect 8260 5720 8266 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 9490 5692 9496 5704
rect 5132 5664 9496 5692
rect 5132 5652 5138 5664
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5692 9643 5695
rect 9674 5692 9680 5704
rect 9631 5664 9680 5692
rect 9631 5661 9643 5664
rect 9585 5655 9643 5661
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 11072 5701 11100 5800
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 12952 5800 12997 5828
rect 12952 5788 12958 5800
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 11204 5732 12449 5760
rect 11204 5720 11210 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 13372 5760 13400 5868
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 16942 5896 16948 5908
rect 16903 5868 16948 5896
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 13722 5788 13728 5840
rect 13780 5788 13786 5840
rect 14185 5831 14243 5837
rect 14185 5797 14197 5831
rect 14231 5828 14243 5831
rect 16298 5828 16304 5840
rect 14231 5800 16304 5828
rect 14231 5797 14243 5800
rect 14185 5791 14243 5797
rect 16298 5788 16304 5800
rect 16356 5788 16362 5840
rect 18874 5828 18880 5840
rect 16408 5800 18276 5828
rect 13449 5763 13507 5769
rect 13449 5760 13461 5763
rect 13372 5732 13461 5760
rect 12437 5723 12495 5729
rect 13449 5729 13461 5732
rect 13495 5760 13507 5763
rect 13538 5760 13544 5772
rect 13495 5732 13544 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13740 5760 13768 5788
rect 16408 5772 16436 5800
rect 15565 5763 15623 5769
rect 13740 5732 13860 5760
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12526 5692 12532 5704
rect 12299 5664 12532 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13722 5692 13728 5704
rect 13311 5664 13728 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 10870 5624 10876 5636
rect 8628 5596 10876 5624
rect 8628 5584 8634 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 10965 5627 11023 5633
rect 10965 5593 10977 5627
rect 11011 5624 11023 5627
rect 11698 5624 11704 5636
rect 11011 5596 11704 5624
rect 11011 5593 11023 5596
rect 10965 5587 11023 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12345 5627 12403 5633
rect 12345 5593 12357 5627
rect 12391 5624 12403 5627
rect 13446 5624 13452 5636
rect 12391 5596 13452 5624
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 13446 5584 13452 5596
rect 13504 5584 13510 5636
rect 13832 5624 13860 5732
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 15746 5760 15752 5772
rect 15611 5732 15752 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 16390 5760 16396 5772
rect 16351 5732 16396 5760
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 16623 5732 17601 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 17589 5729 17601 5732
rect 17635 5760 17647 5763
rect 17678 5760 17684 5772
rect 17635 5732 17684 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 15160 5664 15301 5692
rect 15160 5652 15166 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 13740 5596 13860 5624
rect 14645 5627 14703 5633
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 8386 5556 8392 5568
rect 4304 5528 8392 5556
rect 4304 5516 4310 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 9766 5556 9772 5568
rect 9723 5528 9772 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 11296 5528 11437 5556
rect 11296 5516 11302 5528
rect 11425 5525 11437 5528
rect 11471 5525 11483 5559
rect 11425 5519 11483 5525
rect 13357 5559 13415 5565
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13740 5556 13768 5596
rect 14645 5593 14657 5627
rect 14691 5624 14703 5627
rect 16316 5624 16344 5655
rect 17218 5652 17224 5704
rect 17276 5692 17282 5704
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17276 5664 17325 5692
rect 17276 5652 17282 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 18248 5692 18276 5800
rect 18340 5800 18880 5828
rect 18340 5769 18368 5800
rect 18874 5788 18880 5800
rect 18932 5828 18938 5840
rect 19886 5828 19892 5840
rect 18932 5800 19892 5828
rect 18932 5788 18938 5800
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 20162 5760 20168 5772
rect 19751 5732 20168 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 20162 5720 20168 5732
rect 20220 5760 20226 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20220 5732 21097 5760
rect 20220 5720 20226 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 19889 5695 19947 5701
rect 18248 5664 19840 5692
rect 17313 5655 17371 5661
rect 14691 5596 16344 5624
rect 14691 5593 14703 5596
rect 14645 5587 14703 5593
rect 18138 5584 18144 5636
rect 18196 5624 18202 5636
rect 18414 5624 18420 5636
rect 18196 5596 18420 5624
rect 18196 5584 18202 5596
rect 18414 5584 18420 5596
rect 18472 5584 18478 5636
rect 18509 5627 18567 5633
rect 18509 5593 18521 5627
rect 18555 5624 18567 5627
rect 19610 5624 19616 5636
rect 18555 5596 19616 5624
rect 18555 5593 18567 5596
rect 18509 5587 18567 5593
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 19812 5624 19840 5664
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 20622 5692 20628 5704
rect 19935 5664 20628 5692
rect 19935 5661 19947 5664
rect 19889 5655 19947 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5692 21051 5695
rect 21174 5692 21180 5704
rect 21039 5664 21180 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 20714 5624 20720 5636
rect 19812 5596 20720 5624
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 14918 5556 14924 5568
rect 13403 5528 13768 5556
rect 14879 5528 14924 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15381 5559 15439 5565
rect 15381 5525 15393 5559
rect 15427 5556 15439 5559
rect 15562 5556 15568 5568
rect 15427 5528 15568 5556
rect 15427 5525 15439 5528
rect 15381 5519 15439 5525
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 16114 5516 16120 5568
rect 16172 5556 16178 5568
rect 17405 5559 17463 5565
rect 17405 5556 17417 5559
rect 16172 5528 17417 5556
rect 16172 5516 16178 5528
rect 17405 5525 17417 5528
rect 17451 5525 17463 5559
rect 18874 5556 18880 5568
rect 18835 5528 18880 5556
rect 17405 5519 17463 5525
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20530 5556 20536 5568
rect 20491 5528 20536 5556
rect 20530 5516 20536 5528
rect 20588 5516 20594 5568
rect 20622 5516 20628 5568
rect 20680 5556 20686 5568
rect 20901 5559 20959 5565
rect 20901 5556 20913 5559
rect 20680 5528 20913 5556
rect 20680 5516 20686 5528
rect 20901 5525 20913 5528
rect 20947 5525 20959 5559
rect 20901 5519 20959 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8720 5324 8769 5352
rect 8720 5312 8726 5324
rect 8757 5321 8769 5324
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9674 5352 9680 5364
rect 9539 5324 9680 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 10686 5352 10692 5364
rect 10643 5324 10692 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 10042 5284 10048 5296
rect 8159 5256 10048 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 9125 5083 9183 5089
rect 9125 5080 9137 5083
rect 6788 5052 9137 5080
rect 6788 5040 6794 5052
rect 9125 5049 9137 5052
rect 9171 5080 9183 5083
rect 9876 5080 9904 5179
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 9171 5052 9904 5080
rect 9968 5080 9996 5111
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10612 5148 10640 5315
rect 10686 5312 10692 5324
rect 10744 5352 10750 5364
rect 11057 5355 11115 5361
rect 11057 5352 11069 5355
rect 10744 5324 11069 5352
rect 10744 5312 10750 5324
rect 11057 5321 11069 5324
rect 11103 5321 11115 5355
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11057 5315 11115 5321
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 13449 5355 13507 5361
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 13814 5352 13820 5364
rect 13495 5324 13820 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14826 5352 14832 5364
rect 14787 5324 14832 5352
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15010 5352 15016 5364
rect 14967 5324 15016 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15120 5324 16068 5352
rect 12069 5287 12127 5293
rect 12069 5253 12081 5287
rect 12115 5284 12127 5287
rect 15120 5284 15148 5324
rect 12115 5256 15148 5284
rect 16040 5284 16068 5324
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16666 5352 16672 5364
rect 16172 5324 16672 5352
rect 16172 5312 16178 5324
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 17773 5355 17831 5361
rect 17773 5321 17785 5355
rect 17819 5352 17831 5355
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17819 5324 18337 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 18693 5355 18751 5361
rect 18693 5321 18705 5355
rect 18739 5352 18751 5355
rect 18874 5352 18880 5364
rect 18739 5324 18880 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 19978 5352 19984 5364
rect 19751 5324 19984 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20588 5324 20729 5352
rect 20588 5312 20594 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 16390 5284 16396 5296
rect 16040 5256 16396 5284
rect 12115 5253 12127 5256
rect 12069 5247 12127 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 19794 5284 19800 5296
rect 16500 5256 19800 5284
rect 13354 5216 13360 5228
rect 12360 5188 13360 5216
rect 12158 5148 12164 5160
rect 10192 5120 10640 5148
rect 12119 5120 12164 5148
rect 10192 5108 10198 5120
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12360 5157 12388 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 15841 5220 15899 5225
rect 15764 5219 15899 5220
rect 15764 5216 15853 5219
rect 14200 5192 15853 5216
rect 14200 5188 15792 5192
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 12986 5148 12992 5160
rect 12943 5120 12992 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13262 5148 13268 5160
rect 13223 5120 13268 5148
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 12250 5080 12256 5092
rect 9968 5052 12256 5080
rect 9171 5049 9183 5052
rect 9125 5043 9183 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14200 5089 14228 5188
rect 15841 5185 15853 5192
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5148 14795 5151
rect 15194 5148 15200 5160
rect 14783 5120 15200 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15194 5108 15200 5120
rect 15252 5148 15258 5160
rect 15378 5148 15384 5160
rect 15252 5120 15384 5148
rect 15252 5108 15258 5120
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 14185 5083 14243 5089
rect 14185 5080 14197 5083
rect 13872 5052 14197 5080
rect 13872 5040 13878 5052
rect 14185 5049 14197 5052
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14274 5012 14280 5024
rect 13955 4984 14280 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 15252 4984 15301 5012
rect 15252 4972 15258 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15764 5012 15792 5111
rect 15856 5080 15884 5179
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 16298 5216 16304 5228
rect 15988 5188 16304 5216
rect 15988 5176 15994 5188
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16390 5080 16396 5092
rect 15856 5052 16396 5080
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 16022 5012 16028 5024
rect 15764 4984 16028 5012
rect 15289 4975 15347 4981
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16500 5012 16528 5256
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20809 5287 20867 5293
rect 20809 5284 20821 5287
rect 20312 5256 20821 5284
rect 20312 5244 20318 5256
rect 20809 5253 20821 5256
rect 20855 5253 20867 5287
rect 20809 5247 20867 5253
rect 16666 5216 16672 5228
rect 16627 5188 16672 5216
rect 16666 5176 16672 5188
rect 16724 5176 16730 5228
rect 17678 5216 17684 5228
rect 17639 5188 17684 5216
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 17862 5148 17868 5160
rect 17823 5120 17868 5148
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 16853 5083 16911 5089
rect 16853 5049 16865 5083
rect 16899 5080 16911 5083
rect 18138 5080 18144 5092
rect 16899 5052 18144 5080
rect 16899 5049 16911 5052
rect 16853 5043 16911 5049
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 18800 5080 18828 5111
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19794 5148 19800 5160
rect 19024 5120 19656 5148
rect 19755 5120 19800 5148
rect 19024 5108 19030 5120
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 18800 5052 19349 5080
rect 19337 5049 19349 5052
rect 19383 5049 19395 5083
rect 19628 5080 19656 5120
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 19886 5108 19892 5160
rect 19944 5148 19950 5160
rect 20993 5151 21051 5157
rect 19944 5120 19989 5148
rect 19944 5108 19950 5120
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 21542 5148 21548 5160
rect 21039 5120 21548 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 21542 5108 21548 5120
rect 21600 5108 21606 5160
rect 22922 5080 22928 5092
rect 19628 5052 22928 5080
rect 19337 5043 19395 5049
rect 22922 5040 22928 5052
rect 22980 5040 22986 5092
rect 16347 4984 16528 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17000 4984 17325 5012
rect 17000 4972 17006 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 17313 4975 17371 4981
rect 17586 4972 17592 5024
rect 17644 5012 17650 5024
rect 18874 5012 18880 5024
rect 17644 4984 18880 5012
rect 17644 4972 17650 4984
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9180 4780 9505 4808
rect 9180 4768 9186 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 9493 4771 9551 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 13446 4808 13452 4820
rect 10836 4780 13452 4808
rect 10836 4768 10842 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13596 4780 14105 4808
rect 13596 4768 13602 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 14274 4768 14280 4820
rect 14332 4808 14338 4820
rect 14332 4780 15240 4808
rect 14332 4768 14338 4780
rect 7837 4743 7895 4749
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 15102 4740 15108 4752
rect 7883 4712 15108 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 15212 4740 15240 4780
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 17586 4808 17592 4820
rect 15988 4780 17592 4808
rect 15988 4768 15994 4780
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 17678 4768 17684 4820
rect 17736 4808 17742 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 17736 4780 17877 4808
rect 17736 4768 17742 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 18840 4780 20116 4808
rect 18840 4768 18846 4780
rect 19518 4740 19524 4752
rect 15212 4712 19524 4740
rect 19518 4700 19524 4712
rect 19576 4700 19582 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19852 4712 19993 4740
rect 19852 4700 19858 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 20088 4740 20116 4780
rect 20088 4712 20852 4740
rect 19981 4703 20039 4709
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 7984 4644 9536 4672
rect 7984 4632 7990 4644
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8619 4576 9045 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9033 4573 9045 4576
rect 9079 4604 9091 4607
rect 9398 4604 9404 4616
rect 9079 4576 9404 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9508 4604 9536 4644
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 9950 4672 9956 4684
rect 9732 4644 9956 4672
rect 9732 4632 9738 4644
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4672 10198 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 10192 4644 11161 4672
rect 10192 4632 10198 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11149 4635 11207 4641
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11848 4644 12173 4672
rect 11848 4632 11854 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13173 4675 13231 4681
rect 13173 4672 13185 4675
rect 12952 4644 13185 4672
rect 12952 4632 12958 4644
rect 13173 4641 13185 4644
rect 13219 4672 13231 4675
rect 13538 4672 13544 4684
rect 13219 4644 13544 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 14642 4672 14648 4684
rect 14603 4644 14648 4672
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 15344 4644 15577 4672
rect 15344 4632 15350 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15565 4635 15623 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 18322 4672 18328 4684
rect 15896 4644 17356 4672
rect 18283 4644 18328 4672
rect 15896 4632 15902 4644
rect 9861 4607 9919 4613
rect 9508 4576 9674 4604
rect 8205 4539 8263 4545
rect 8205 4505 8217 4539
rect 8251 4536 8263 4539
rect 9306 4536 9312 4548
rect 8251 4508 9312 4536
rect 8251 4505 8263 4508
rect 8205 4499 8263 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 9490 4468 9496 4480
rect 9263 4440 9496 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9646 4468 9674 4576
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 10962 4604 10968 4616
rect 9907 4576 10968 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12710 4604 12716 4616
rect 12115 4576 12716 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12986 4604 12992 4616
rect 12947 4576 12992 4604
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13446 4564 13452 4616
rect 13504 4604 13510 4616
rect 15470 4604 15476 4616
rect 13504 4576 15332 4604
rect 15431 4576 15476 4604
rect 13504 4564 13510 4576
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 11057 4539 11115 4545
rect 11057 4536 11069 4539
rect 10928 4508 11069 4536
rect 10928 4496 10934 4508
rect 11057 4505 11069 4508
rect 11103 4505 11115 4539
rect 11057 4499 11115 4505
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 13081 4539 13139 4545
rect 12023 4508 12434 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 10965 4471 11023 4477
rect 10965 4468 10977 4471
rect 9646 4440 10977 4468
rect 10965 4437 10977 4440
rect 11011 4468 11023 4471
rect 11146 4468 11152 4480
rect 11011 4440 11152 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 11698 4468 11704 4480
rect 11655 4440 11704 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 12406 4468 12434 4508
rect 13081 4505 13093 4539
rect 13127 4536 13139 4539
rect 15304 4536 15332 4576
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 16942 4604 16948 4616
rect 16899 4576 16948 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 16408 4536 16436 4567
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17328 4613 17356 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4672 18567 4675
rect 18966 4672 18972 4684
rect 18555 4644 18972 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 20622 4672 20628 4684
rect 19751 4644 20628 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 20824 4681 20852 4712
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4641 20867 4675
rect 20809 4635 20867 4641
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 20533 4607 20591 4613
rect 20533 4604 20545 4607
rect 19208 4576 20545 4604
rect 19208 4564 19214 4576
rect 20533 4573 20545 4576
rect 20579 4604 20591 4607
rect 20714 4604 20720 4616
rect 20579 4576 20720 4604
rect 20579 4573 20591 4576
rect 20533 4567 20591 4573
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 17954 4536 17960 4548
rect 13127 4508 15148 4536
rect 15304 4508 17960 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 12406 4440 12633 4468
rect 12621 4437 12633 4440
rect 12667 4437 12679 4471
rect 12621 4431 12679 4437
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 13814 4468 13820 4480
rect 13771 4440 13820 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14240 4440 14473 4468
rect 14240 4428 14246 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14461 4431 14519 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15120 4477 15148 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 19242 4496 19248 4548
rect 19300 4536 19306 4548
rect 20165 4539 20223 4545
rect 20165 4536 20177 4539
rect 19300 4508 20177 4536
rect 19300 4496 19306 4508
rect 20165 4505 20177 4508
rect 20211 4505 20223 4539
rect 20165 4499 20223 4505
rect 15105 4471 15163 4477
rect 14608 4440 14653 4468
rect 14608 4428 14614 4440
rect 15105 4437 15117 4471
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 15286 4428 15292 4480
rect 15344 4468 15350 4480
rect 15746 4468 15752 4480
rect 15344 4440 15752 4468
rect 15344 4428 15350 4440
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16577 4471 16635 4477
rect 16577 4437 16589 4471
rect 16623 4468 16635 4471
rect 16942 4468 16948 4480
rect 16623 4440 16948 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17037 4471 17095 4477
rect 17037 4437 17049 4471
rect 17083 4468 17095 4471
rect 17126 4468 17132 4480
rect 17083 4440 17132 4468
rect 17083 4437 17095 4440
rect 17037 4431 17095 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17497 4471 17555 4477
rect 17497 4437 17509 4471
rect 17543 4468 17555 4471
rect 17586 4468 17592 4480
rect 17543 4440 17592 4468
rect 17543 4437 17555 4440
rect 17497 4431 17555 4437
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 10413 4267 10471 4273
rect 10413 4233 10425 4267
rect 10459 4264 10471 4267
rect 11054 4264 11060 4276
rect 10459 4236 11060 4264
rect 10459 4233 10471 4236
rect 10413 4227 10471 4233
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11204 4236 12112 4264
rect 11204 4224 11210 4236
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 9677 4199 9735 4205
rect 9456 4168 9628 4196
rect 9456 4156 9462 4168
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9600 4128 9628 4168
rect 9677 4165 9689 4199
rect 9723 4196 9735 4199
rect 10778 4196 10784 4208
rect 9723 4168 10784 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11440 4168 11897 4196
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 9600 4100 10701 4128
rect 10689 4097 10701 4100
rect 10735 4128 10747 4131
rect 11440 4128 11468 4168
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 12084 4196 12112 4236
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 12253 4267 12311 4273
rect 12253 4264 12265 4267
rect 12216 4236 12265 4264
rect 12216 4224 12222 4236
rect 12253 4233 12265 4236
rect 12299 4233 12311 4267
rect 12253 4227 12311 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 12989 4267 13047 4273
rect 12989 4264 13001 4267
rect 12768 4236 13001 4264
rect 12768 4224 12774 4236
rect 12989 4233 13001 4236
rect 13035 4233 13047 4267
rect 14182 4264 14188 4276
rect 14143 4236 14188 4264
rect 12989 4227 13047 4233
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 15286 4264 15292 4276
rect 14424 4236 15292 4264
rect 14424 4224 14430 4236
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15749 4267 15807 4273
rect 15749 4264 15761 4267
rect 15528 4236 15761 4264
rect 15528 4224 15534 4236
rect 15749 4233 15761 4236
rect 15795 4233 15807 4267
rect 15749 4227 15807 4233
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 18230 4264 18236 4276
rect 17000 4236 18000 4264
rect 18191 4236 18236 4264
rect 17000 4224 17006 4236
rect 13357 4199 13415 4205
rect 12084 4168 13308 4196
rect 11885 4159 11943 4165
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 10735 4100 11468 4128
rect 11624 4100 11805 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 8846 4060 8852 4072
rect 8807 4032 8852 4060
rect 8846 4020 8852 4032
rect 8904 4060 8910 4072
rect 9766 4060 9772 4072
rect 8904 4032 9772 4060
rect 8904 4020 8910 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10962 4060 10968 4072
rect 10091 4032 10968 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 10962 4020 10968 4032
rect 11020 4060 11026 4072
rect 11624 4060 11652 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 12618 4128 12624 4140
rect 11793 4091 11851 4097
rect 12360 4100 12624 4128
rect 11020 4032 11652 4060
rect 11701 4063 11759 4069
rect 11020 4020 11026 4032
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 11974 4060 11980 4072
rect 11747 4032 11980 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 7469 3995 7527 4001
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 12360 3992 12388 4100
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 13078 4128 13084 4140
rect 12759 4100 13084 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13280 4128 13308 4168
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 14918 4196 14924 4208
rect 13403 4168 14924 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 15105 4199 15163 4205
rect 15105 4165 15117 4199
rect 15151 4196 15163 4199
rect 16574 4196 16580 4208
rect 15151 4168 16580 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 16574 4156 16580 4168
rect 16632 4156 16638 4208
rect 17972 4196 18000 4236
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 18693 4267 18751 4273
rect 18693 4233 18705 4267
rect 18739 4233 18751 4267
rect 18693 4227 18751 4233
rect 18414 4196 18420 4208
rect 17972 4168 18420 4196
rect 18414 4156 18420 4168
rect 18472 4156 18478 4208
rect 13280 4100 13768 4128
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 13740 4060 13768 4100
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 13872 4100 14473 4128
rect 13872 4088 13878 4100
rect 14461 4097 14473 4100
rect 14507 4128 14519 4131
rect 14642 4128 14648 4140
rect 14507 4100 14648 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15930 4128 15936 4140
rect 14752 4100 15936 4128
rect 14752 4060 14780 4100
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16448 4100 16681 4128
rect 16448 4088 16454 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 13596 4032 13641 4060
rect 13740 4032 14780 4060
rect 13596 4020 13602 4032
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15436 4032 15485 4060
rect 15436 4020 15442 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15654 4060 15660 4072
rect 15615 4032 15660 4060
rect 15473 4023 15531 4029
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 17328 4060 17356 4091
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17736 4100 17785 4128
rect 17736 4088 17742 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 18708 4060 18736 4227
rect 20165 4199 20223 4205
rect 20165 4165 20177 4199
rect 20211 4196 20223 4199
rect 20438 4196 20444 4208
rect 20211 4168 20444 4196
rect 20211 4165 20223 4168
rect 20165 4159 20223 4165
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 17328 4032 18736 4060
rect 18892 4060 18920 4091
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19024 4100 19441 4128
rect 19024 4088 19030 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 19429 4091 19487 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20680 4100 20821 4128
rect 20680 4088 20686 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 20346 4060 20352 4072
rect 18892 4032 20352 4060
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 7515 3964 12388 3992
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 14826 3992 14832 4004
rect 12676 3964 14832 3992
rect 12676 3952 12682 3964
rect 14826 3952 14832 3964
rect 14884 3952 14890 4004
rect 16853 3995 16911 4001
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 17218 3992 17224 4004
rect 16899 3964 17224 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 17218 3952 17224 3964
rect 17276 3952 17282 4004
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 19613 3995 19671 4001
rect 17828 3964 19334 3992
rect 17828 3952 17834 3964
rect 1394 3924 1400 3936
rect 1355 3896 1400 3924
rect 1394 3884 1400 3896
rect 1452 3884 1458 3936
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 8076 3896 8125 3924
rect 8076 3884 8082 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 8113 3887 8171 3893
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 9214 3924 9220 3936
rect 8628 3896 9220 3924
rect 8628 3884 8634 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 14645 3927 14703 3933
rect 12584 3896 12629 3924
rect 12584 3884 12590 3896
rect 14645 3893 14657 3927
rect 14691 3924 14703 3927
rect 15930 3924 15936 3936
rect 14691 3896 15936 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16666 3924 16672 3936
rect 16163 3896 16672 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17497 3927 17555 3933
rect 17497 3893 17509 3927
rect 17543 3924 17555 3927
rect 17678 3924 17684 3936
rect 17543 3896 17684 3924
rect 17543 3893 17555 3896
rect 17497 3887 17555 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17957 3927 18015 3933
rect 17957 3893 17969 3927
rect 18003 3924 18015 3927
rect 19058 3924 19064 3936
rect 18003 3896 19064 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19306 3924 19334 3964
rect 19613 3961 19625 3995
rect 19659 3992 19671 3995
rect 22462 3992 22468 4004
rect 19659 3964 22468 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 22462 3952 22468 3964
rect 22520 3952 22526 4004
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 19306 3896 20085 3924
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 6822 3720 6828 3732
rect 1627 3692 6828 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 18233 3723 18291 3729
rect 7147 3692 18184 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7837 3655 7895 3661
rect 7837 3621 7849 3655
rect 7883 3652 7895 3655
rect 8202 3652 8208 3664
rect 7883 3624 8208 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9858 3652 9864 3664
rect 9819 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10502 3652 10508 3664
rect 10008 3624 10508 3652
rect 10008 3612 10014 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 10962 3652 10968 3664
rect 10923 3624 10968 3652
rect 10962 3612 10968 3624
rect 11020 3652 11026 3664
rect 12986 3652 12992 3664
rect 11020 3624 12992 3652
rect 11020 3612 11026 3624
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 18156 3652 18184 3692
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 18966 3720 18972 3732
rect 18279 3692 18972 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 18598 3652 18604 3664
rect 15620 3624 16804 3652
rect 18156 3624 18604 3652
rect 15620 3612 15626 3624
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3584 7527 3587
rect 14829 3587 14887 3593
rect 7515 3556 14780 3584
rect 7515 3553 7527 3556
rect 7469 3547 7527 3553
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3516 1455 3519
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1443 3488 1869 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 1857 3485 1869 3488
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 5776 3488 8493 3516
rect 5776 3476 5782 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 10962 3516 10968 3528
rect 9539 3488 10968 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 2225 3451 2283 3457
rect 2225 3448 2237 3451
rect 1544 3420 2237 3448
rect 1544 3408 1550 3420
rect 2225 3417 2237 3420
rect 2271 3417 2283 3451
rect 2225 3411 2283 3417
rect 6733 3451 6791 3457
rect 6733 3417 6745 3451
rect 6779 3448 6791 3451
rect 8294 3448 8300 3460
rect 6779 3420 8300 3448
rect 6779 3417 6791 3420
rect 6733 3411 6791 3417
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4890 3380 4896 3392
rect 4847 3352 4896 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5902 3340 5908 3392
rect 5960 3380 5966 3392
rect 6089 3383 6147 3389
rect 6089 3380 6101 3383
rect 5960 3352 6101 3380
rect 5960 3340 5966 3352
rect 6089 3349 6101 3352
rect 6135 3349 6147 3383
rect 6089 3343 6147 3349
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8386 3380 8392 3392
rect 8251 3352 8392 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8496 3380 8524 3479
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 11296 3488 11345 3516
rect 11296 3476 11302 3488
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 11333 3479 11391 3485
rect 11532 3488 11805 3516
rect 9125 3451 9183 3457
rect 9125 3417 9137 3451
rect 9171 3448 9183 3451
rect 9950 3448 9956 3460
rect 9171 3420 9956 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 8496 3352 10149 3380
rect 10137 3349 10149 3352
rect 10183 3380 10195 3383
rect 11238 3380 11244 3392
rect 10183 3352 11244 3380
rect 10183 3349 10195 3352
rect 10137 3343 10195 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11532 3389 11560 3488
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12526 3516 12532 3528
rect 12299 3488 12532 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 14752 3516 14780 3556
rect 14829 3553 14841 3587
rect 14875 3584 14887 3587
rect 14918 3584 14924 3596
rect 14875 3556 14924 3584
rect 14875 3553 14887 3556
rect 14829 3547 14887 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 15436 3556 15761 3584
rect 15436 3544 15442 3556
rect 15749 3553 15761 3556
rect 15795 3553 15807 3587
rect 16666 3584 16672 3596
rect 16627 3556 16672 3584
rect 15749 3547 15807 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 16776 3593 16804 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 19150 3652 19156 3664
rect 18748 3624 19156 3652
rect 18748 3612 18754 3624
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 19613 3655 19671 3661
rect 19613 3621 19625 3655
rect 19659 3652 19671 3655
rect 21542 3652 21548 3664
rect 19659 3624 21548 3652
rect 19659 3621 19671 3624
rect 19613 3615 19671 3621
rect 21542 3612 21548 3624
rect 21600 3612 21606 3664
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3553 16819 3587
rect 16761 3547 16819 3553
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 17368 3556 17724 3584
rect 17368 3544 17374 3556
rect 16574 3516 16580 3528
rect 13219 3488 14228 3516
rect 14752 3488 16436 3516
rect 16535 3488 16580 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 12728 3448 12756 3479
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 12400 3420 13645 3448
rect 12400 3408 12406 3420
rect 13633 3417 13645 3420
rect 13679 3417 13691 3451
rect 13633 3411 13691 3417
rect 11517 3383 11575 3389
rect 11517 3349 11529 3383
rect 11563 3349 11575 3383
rect 11517 3343 11575 3349
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3380 12035 3383
rect 12066 3380 12072 3392
rect 12023 3352 12072 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12618 3380 12624 3392
rect 12483 3352 12624 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12894 3380 12900 3392
rect 12855 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13354 3380 13360 3392
rect 13315 3352 13360 3380
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14200 3389 14228 3488
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 16408 3448 16436 3488
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17460 3488 17601 3516
rect 17460 3476 17466 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17696 3516 17724 3556
rect 17954 3544 17960 3596
rect 18012 3584 18018 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 18012 3556 19993 3584
rect 18012 3544 18018 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17696 3488 18061 3516
rect 17589 3479 17647 3485
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 18049 3479 18107 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20530 3516 20536 3528
rect 19536 3488 20536 3516
rect 14599 3420 16252 3448
rect 16408 3420 17908 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14185 3383 14243 3389
rect 14185 3349 14197 3383
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 14826 3380 14832 3392
rect 14691 3352 14832 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 15286 3380 15292 3392
rect 15243 3352 15292 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 15565 3383 15623 3389
rect 15565 3380 15577 3383
rect 15528 3352 15577 3380
rect 15528 3340 15534 3352
rect 15565 3349 15577 3352
rect 15611 3349 15623 3383
rect 15565 3343 15623 3349
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 16224 3389 16252 3420
rect 16209 3383 16267 3389
rect 15712 3352 15757 3380
rect 15712 3340 15718 3352
rect 16209 3349 16221 3383
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 16356 3352 17233 3380
rect 16356 3340 16362 3352
rect 17221 3349 17233 3352
rect 17267 3380 17279 3383
rect 17310 3380 17316 3392
rect 17267 3352 17316 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17770 3380 17776 3392
rect 17731 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 17880 3380 17908 3420
rect 18598 3408 18604 3460
rect 18656 3448 18662 3460
rect 19536 3448 19564 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 20162 3448 20168 3460
rect 18656 3420 19564 3448
rect 20123 3420 20168 3448
rect 18656 3408 18662 3420
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 18506 3380 18512 3392
rect 17880 3352 18512 3380
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 18690 3380 18696 3392
rect 18651 3352 18696 3380
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 20824 3380 20852 3479
rect 18840 3352 20852 3380
rect 18840 3340 18846 3352
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3145 1823 3179
rect 7282 3176 7288 3188
rect 1765 3139 1823 3145
rect 2746 3148 7288 3176
rect 1780 3108 1808 3139
rect 2746 3108 2774 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 9493 3179 9551 3185
rect 9493 3145 9505 3179
rect 9539 3176 9551 3179
rect 11146 3176 11152 3188
rect 9539 3148 11152 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 11839 3148 12434 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 1780 3080 2774 3108
rect 5350 3068 5356 3120
rect 5408 3108 5414 3120
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 5408 3080 5549 3108
rect 5408 3068 5414 3080
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 5718 3108 5724 3120
rect 5679 3080 5724 3108
rect 5537 3071 5595 3077
rect 5718 3068 5724 3080
rect 5776 3108 5782 3120
rect 8478 3108 8484 3120
rect 5776 3080 8484 3108
rect 5776 3068 5782 3080
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 9033 3111 9091 3117
rect 9033 3077 9045 3111
rect 9079 3108 9091 3111
rect 9079 3080 10088 3108
rect 9079 3077 9091 3080
rect 9033 3071 9091 3077
rect 10060 3052 10088 3080
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1544 3012 1593 3040
rect 1544 3000 1550 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4522 3040 4528 3052
rect 4111 3012 4528 3040
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4890 3040 4896 3052
rect 4851 3012 4896 3040
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8110 3040 8116 3052
rect 7607 3012 8116 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 9214 3040 9220 3052
rect 8343 3012 9220 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 9214 3000 9220 3012
rect 9272 3040 9278 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 9272 3012 9321 3040
rect 9272 3000 9278 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9824 3012 9873 3040
rect 9824 3000 9830 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10100 3012 10977 3040
rect 10100 3000 10106 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11609 3043 11667 3049
rect 11609 3009 11621 3043
rect 11655 3040 11667 3043
rect 11698 3040 11704 3052
rect 11655 3012 11704 3040
rect 11655 3009 11667 3012
rect 11609 3003 11667 3009
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12406 3040 12434 3148
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13504 3148 13829 3176
rect 13504 3136 13510 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 13817 3139 13875 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14826 3176 14832 3188
rect 14787 3148 14832 3176
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15286 3176 15292 3188
rect 15247 3148 15292 3176
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 18969 3179 19027 3185
rect 18969 3176 18981 3179
rect 18932 3148 18981 3176
rect 18932 3136 18938 3148
rect 18969 3145 18981 3148
rect 19015 3145 19027 3179
rect 18969 3139 19027 3145
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 19208 3148 20852 3176
rect 19208 3136 19214 3148
rect 13354 3068 13360 3120
rect 13412 3108 13418 3120
rect 15194 3108 15200 3120
rect 13412 3080 14780 3108
rect 15155 3080 15200 3108
rect 13412 3068 13418 3080
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12406 3012 12541 3040
rect 12069 3003 12127 3009
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12529 3003 12587 3009
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3476 2944 3525 2972
rect 3476 2932 3482 2944
rect 3513 2941 3525 2944
rect 3559 2972 3571 2975
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3559 2944 3801 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 9732 2944 10241 2972
rect 9732 2932 9738 2944
rect 10229 2941 10241 2944
rect 10275 2972 10287 2975
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10275 2944 10609 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 10597 2941 10609 2944
rect 10643 2972 10655 2975
rect 12084 2972 12112 3003
rect 12986 3000 12992 3012
rect 13044 3040 13050 3052
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13044 3012 13461 3040
rect 13044 3000 13050 3012
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 14752 3040 14780 3080
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 15988 3080 19472 3108
rect 15988 3068 15994 3080
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 14752 3012 16037 3040
rect 13449 3003 13507 3009
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 16853 3003 16911 3009
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 10643 2944 14289 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 15473 2975 15531 2981
rect 14424 2944 14469 2972
rect 14424 2932 14430 2944
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 15562 2972 15568 2984
rect 15519 2944 15568 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 16868 2972 16896 3003
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 17862 3040 17868 3052
rect 17696 3012 17868 3040
rect 15672 2944 16896 2972
rect 15672 2916 15700 2944
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 17696 2972 17724 3012
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18874 3040 18880 3052
rect 18564 3012 18880 3040
rect 18564 3000 18570 3012
rect 18874 3000 18880 3012
rect 18932 3040 18938 3052
rect 19444 3049 19472 3080
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18932 3012 19073 3040
rect 18932 3000 18938 3012
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 20530 3040 20536 3052
rect 20491 3012 20536 3040
rect 19981 3003 20039 3009
rect 19996 2972 20024 3003
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 20824 3049 20852 3148
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 17276 2944 17724 2972
rect 17788 2944 20024 2972
rect 17276 2932 17282 2944
rect 5074 2904 5080 2916
rect 5035 2876 5080 2904
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 7558 2904 7564 2916
rect 7239 2876 7564 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8665 2907 8723 2913
rect 8665 2873 8677 2907
rect 8711 2904 8723 2907
rect 10502 2904 10508 2916
rect 8711 2876 10508 2904
rect 8711 2873 8723 2876
rect 8665 2867 8723 2873
rect 10502 2864 10508 2876
rect 10560 2864 10566 2916
rect 11146 2904 11152 2916
rect 11107 2876 11152 2904
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 11238 2864 11244 2916
rect 11296 2904 11302 2916
rect 15654 2904 15660 2916
rect 11296 2876 15660 2904
rect 11296 2864 11302 2876
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 17788 2913 17816 2944
rect 17773 2907 17831 2913
rect 16264 2876 17448 2904
rect 16264 2864 16270 2876
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 2096 2808 2329 2836
rect 2096 2796 2102 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2317 2799 2375 2805
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3142 2836 3148 2848
rect 2832 2808 2877 2836
rect 3103 2808 3148 2836
rect 2832 2796 2838 2808
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 6546 2836 6552 2848
rect 6503 2808 6552 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 6825 2839 6883 2845
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 7006 2836 7012 2848
rect 6871 2808 7012 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8478 2836 8484 2848
rect 7975 2808 8484 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12342 2836 12348 2848
rect 12299 2808 12348 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 12710 2836 12716 2848
rect 12671 2808 12716 2836
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 13173 2839 13231 2845
rect 13173 2805 13185 2839
rect 13219 2836 13231 2839
rect 13354 2836 13360 2848
rect 13219 2808 13360 2836
rect 13219 2805 13231 2808
rect 13173 2799 13231 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15841 2839 15899 2845
rect 15841 2836 15853 2839
rect 15252 2808 15853 2836
rect 15252 2796 15258 2808
rect 15841 2805 15853 2808
rect 15887 2805 15899 2839
rect 16666 2836 16672 2848
rect 16627 2808 16672 2836
rect 15841 2799 15899 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 17276 2808 17325 2836
rect 17276 2796 17282 2808
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 17420 2836 17448 2876
rect 17773 2873 17785 2907
rect 17819 2873 17831 2907
rect 18782 2904 18788 2916
rect 17773 2867 17831 2873
rect 17880 2876 18788 2904
rect 17880 2836 17908 2876
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 19613 2907 19671 2913
rect 19613 2873 19625 2907
rect 19659 2904 19671 2907
rect 21358 2904 21364 2916
rect 19659 2876 21364 2904
rect 19659 2873 19671 2876
rect 19613 2867 19671 2873
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 17420 2808 17908 2836
rect 17313 2799 17371 2805
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18325 2839 18383 2845
rect 18325 2836 18337 2839
rect 18104 2808 18337 2836
rect 18104 2796 18110 2808
rect 18325 2805 18337 2808
rect 18371 2805 18383 2839
rect 18325 2799 18383 2805
rect 20165 2839 20223 2845
rect 20165 2805 20177 2839
rect 20211 2836 20223 2839
rect 20806 2836 20812 2848
rect 20211 2808 20812 2836
rect 20211 2805 20223 2808
rect 20165 2799 20223 2805
rect 20806 2796 20812 2808
rect 20864 2796 20870 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 5776 2604 6745 2632
rect 5776 2592 5782 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7708 2604 7849 2632
rect 7708 2592 7714 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 7984 2604 8401 2632
rect 7984 2592 7990 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 8389 2595 8447 2601
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10284 2604 10609 2632
rect 10284 2592 10290 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 14550 2632 14556 2644
rect 11195 2604 14556 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 14700 2604 16896 2632
rect 14700 2592 14706 2604
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 10137 2567 10195 2573
rect 3283 2536 9444 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4614 2496 4620 2508
rect 4111 2468 4476 2496
rect 4575 2468 4620 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 382 2388 388 2440
rect 440 2428 446 2440
rect 1394 2428 1400 2440
rect 440 2400 1400 2428
rect 440 2388 446 2400
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2832 2400 3065 2428
rect 2832 2388 2838 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4304 2400 4353 2428
rect 4304 2388 4310 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4448 2428 4476 2468
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5684 2468 5733 2496
rect 5684 2456 5690 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9306 2496 9312 2508
rect 9263 2468 9312 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 5994 2428 6000 2440
rect 4448 2400 6000 2428
rect 4341 2391 4399 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 7064 2400 7113 2428
rect 7064 2388 7070 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8662 2428 8668 2440
rect 8536 2400 8668 2428
rect 8536 2388 8542 2400
rect 8662 2388 8668 2400
rect 8720 2428 8726 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8720 2400 9045 2428
rect 8720 2388 8726 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 2038 2320 2044 2372
rect 2096 2360 2102 2372
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 2096 2332 2605 2360
rect 2096 2320 2102 2332
rect 2593 2329 2605 2332
rect 2639 2329 2651 2363
rect 2593 2323 2651 2329
rect 3142 2320 3148 2372
rect 3200 2360 3206 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3200 2332 3893 2360
rect 3200 2320 3206 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 5902 2360 5908 2372
rect 5863 2332 5908 2360
rect 3881 2323 3939 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 6604 2332 6653 2360
rect 6604 2320 6610 2332
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 6641 2323 6699 2329
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 7745 2363 7803 2369
rect 7745 2360 7757 2363
rect 7616 2332 7757 2360
rect 7616 2320 7622 2332
rect 7745 2329 7757 2332
rect 7791 2329 7803 2363
rect 8294 2360 8300 2372
rect 8255 2332 8300 2360
rect 7745 2323 7803 2329
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 9416 2360 9444 2536
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 10410 2564 10416 2576
rect 10183 2536 10416 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 11793 2567 11851 2573
rect 11793 2533 11805 2567
rect 11839 2564 11851 2567
rect 13630 2564 13636 2576
rect 11839 2536 13636 2564
rect 11839 2533 11851 2536
rect 11793 2527 11851 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 14182 2524 14188 2576
rect 14240 2564 14246 2576
rect 14737 2567 14795 2573
rect 14737 2564 14749 2567
rect 14240 2536 14749 2564
rect 14240 2524 14246 2536
rect 14737 2533 14749 2536
rect 14783 2533 14795 2567
rect 14737 2527 14795 2533
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15344 2536 15945 2564
rect 15344 2524 15350 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 16080 2536 16804 2564
rect 16080 2524 16086 2536
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 10870 2496 10876 2508
rect 9631 2468 10876 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 10870 2456 10876 2468
rect 10928 2496 10934 2508
rect 12802 2496 12808 2508
rect 10928 2468 11652 2496
rect 10928 2456 10934 2468
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11624 2437 11652 2468
rect 11716 2468 12808 2496
rect 11609 2431 11667 2437
rect 11609 2397 11621 2431
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 11514 2360 11520 2372
rect 9416 2332 11520 2360
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 2685 2295 2743 2301
rect 2685 2261 2697 2295
rect 2731 2292 2743 2295
rect 6730 2292 6736 2304
rect 2731 2264 6736 2292
rect 2731 2261 2743 2264
rect 2685 2255 2743 2261
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2292 7343 2295
rect 11716 2292 11744 2468
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 12894 2456 12900 2508
rect 12952 2496 12958 2508
rect 12952 2468 15240 2496
rect 12952 2456 12958 2468
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12768 2400 13185 2428
rect 12768 2388 12774 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13354 2388 13360 2440
rect 13412 2428 13418 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13412 2400 14105 2428
rect 13412 2388 13418 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2424 14979 2431
rect 15102 2428 15108 2440
rect 15028 2424 15108 2428
rect 14967 2400 15108 2424
rect 14967 2397 15056 2400
rect 14921 2396 15056 2397
rect 14921 2391 14979 2396
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15212 2437 15240 2468
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 15749 2391 15807 2397
rect 12342 2320 12348 2372
rect 12400 2360 12406 2372
rect 15764 2360 15792 2391
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 16776 2428 16804 2536
rect 16868 2496 16896 2604
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17957 2635 18015 2641
rect 17957 2632 17969 2635
rect 17000 2604 17969 2632
rect 17000 2592 17006 2604
rect 17957 2601 17969 2604
rect 18003 2601 18015 2635
rect 17957 2595 18015 2601
rect 17494 2524 17500 2576
rect 17552 2564 17558 2576
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 17552 2536 18521 2564
rect 17552 2524 17558 2536
rect 18509 2533 18521 2536
rect 18555 2533 18567 2567
rect 18509 2527 18567 2533
rect 19150 2524 19156 2576
rect 19208 2564 19214 2576
rect 19981 2567 20039 2573
rect 19981 2564 19993 2567
rect 19208 2536 19993 2564
rect 19208 2524 19214 2536
rect 19981 2533 19993 2536
rect 20027 2533 20039 2567
rect 19981 2527 20039 2533
rect 20254 2524 20260 2576
rect 20312 2564 20318 2576
rect 21085 2567 21143 2573
rect 21085 2564 21097 2567
rect 20312 2536 21097 2564
rect 20312 2524 20318 2536
rect 21085 2533 21097 2536
rect 21131 2533 21143 2567
rect 21085 2527 21143 2533
rect 16868 2468 17540 2496
rect 17034 2428 17040 2440
rect 16776 2400 17040 2428
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 17218 2428 17224 2440
rect 17179 2400 17224 2428
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 12400 2332 15792 2360
rect 12400 2320 12406 2332
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 17512 2360 17540 2468
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17736 2468 18460 2496
rect 17736 2456 17742 2468
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17920 2400 18337 2428
rect 17920 2388 17926 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18432 2428 18460 2468
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 18748 2468 20392 2496
rect 18748 2456 18754 2468
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18432 2400 19257 2428
rect 18325 2391 18383 2397
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19794 2428 19800 2440
rect 19755 2400 19800 2428
rect 19245 2391 19303 2397
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 20364 2437 20392 2468
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 18966 2360 18972 2372
rect 16448 2332 17448 2360
rect 17512 2332 18972 2360
rect 16448 2320 16454 2332
rect 7331 2264 11744 2292
rect 7331 2261 7343 2264
rect 7285 2255 7343 2261
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12032 2264 12265 2292
rect 12032 2252 12038 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12253 2255 12311 2261
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12584 2264 12817 2292
rect 12584 2252 12590 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13136 2264 13369 2292
rect 13136 2252 13142 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13688 2264 14289 2292
rect 13688 2252 13694 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 14792 2264 15393 2292
rect 14792 2252 14798 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 17420 2301 17448 2332
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 19058 2320 19064 2372
rect 19116 2360 19122 2372
rect 20916 2360 20944 2391
rect 19116 2332 20944 2360
rect 19116 2320 19122 2332
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 15896 2264 16865 2292
rect 15896 2252 15902 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18656 2264 19441 2292
rect 18656 2252 18662 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 20533 2295 20591 2301
rect 20533 2292 20545 2295
rect 19760 2264 20545 2292
rect 19760 2252 19766 2264
rect 20533 2261 20545 2264
rect 20579 2261 20591 2295
rect 20533 2255 20591 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 8018 2048 8024 2100
rect 8076 2088 8082 2100
rect 16022 2088 16028 2100
rect 8076 2060 16028 2088
rect 8076 2048 8082 2060
rect 16022 2048 16028 2060
rect 16080 2048 16086 2100
rect 19794 2088 19800 2100
rect 16546 2060 19800 2088
rect 7834 1980 7840 2032
rect 7892 2020 7898 2032
rect 14642 2020 14648 2032
rect 7892 1992 14648 2020
rect 7892 1980 7898 1992
rect 14642 1980 14648 1992
rect 14700 1980 14706 2032
rect 16546 2020 16574 2060
rect 19794 2048 19800 2060
rect 19852 2048 19858 2100
rect 14844 1992 16574 2020
rect 9490 1912 9496 1964
rect 9548 1952 9554 1964
rect 14844 1952 14872 1992
rect 17034 1980 17040 2032
rect 17092 2020 17098 2032
rect 20438 2020 20444 2032
rect 17092 1992 20444 2020
rect 17092 1980 17098 1992
rect 20438 1980 20444 1992
rect 20496 1980 20502 2032
rect 9548 1924 14872 1952
rect 9548 1912 9554 1924
rect 14918 1912 14924 1964
rect 14976 1952 14982 1964
rect 22646 1952 22652 1964
rect 14976 1924 22652 1952
rect 14976 1912 14982 1924
rect 22646 1912 22652 1924
rect 22704 1912 22710 1964
rect 1670 1708 1676 1760
rect 1728 1748 1734 1760
rect 13722 1748 13728 1760
rect 1728 1720 13728 1748
rect 1728 1708 1734 1720
rect 13722 1708 13728 1720
rect 13780 1708 13786 1760
<< via1 >>
rect 14556 20816 14608 20868
rect 17960 20816 18012 20868
rect 2320 20748 2372 20800
rect 20352 20748 20404 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 12532 20544 12584 20596
rect 13084 20544 13136 20596
rect 13820 20544 13872 20596
rect 14740 20544 14792 20596
rect 15844 20544 15896 20596
rect 17500 20544 17552 20596
rect 18604 20544 18656 20596
rect 3884 20476 3936 20528
rect 10324 20476 10376 20528
rect 11704 20476 11756 20528
rect 388 20408 440 20460
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 3056 20408 3108 20460
rect 3700 20408 3752 20460
rect 4252 20408 4304 20460
rect 4988 20451 5040 20460
rect 4988 20417 4997 20451
rect 4997 20417 5031 20451
rect 5031 20417 5040 20451
rect 4988 20408 5040 20417
rect 5080 20408 5132 20460
rect 5356 20408 5408 20460
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 2136 20340 2188 20392
rect 3240 20340 3292 20392
rect 4436 20340 4488 20392
rect 6000 20340 6052 20392
rect 6552 20383 6604 20392
rect 6552 20349 6561 20383
rect 6561 20349 6595 20383
rect 6595 20349 6604 20383
rect 6552 20340 6604 20349
rect 6920 20340 6972 20392
rect 7656 20383 7708 20392
rect 7656 20349 7665 20383
rect 7665 20349 7699 20383
rect 7699 20349 7708 20383
rect 7656 20340 7708 20349
rect 4712 20272 4764 20324
rect 9312 20340 9364 20392
rect 10324 20340 10376 20392
rect 11060 20340 11112 20392
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 11612 20340 11664 20392
rect 12072 20340 12124 20392
rect 13268 20408 13320 20460
rect 15200 20451 15252 20460
rect 13544 20340 13596 20392
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15384 20408 15436 20460
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18512 20408 18564 20460
rect 20076 20408 20128 20460
rect 16764 20340 16816 20392
rect 20260 20340 20312 20392
rect 3424 20204 3476 20256
rect 11888 20272 11940 20324
rect 4896 20204 4948 20256
rect 5540 20204 5592 20256
rect 8668 20204 8720 20256
rect 10692 20204 10744 20256
rect 12532 20272 12584 20324
rect 14188 20272 14240 20324
rect 15292 20272 15344 20324
rect 16396 20272 16448 20324
rect 18144 20272 18196 20324
rect 19156 20272 19208 20324
rect 16948 20204 17000 20256
rect 18696 20204 18748 20256
rect 20720 20204 20772 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 3424 20043 3476 20052
rect 3424 20009 3433 20043
rect 3433 20009 3467 20043
rect 3467 20009 3476 20043
rect 3424 20000 3476 20009
rect 3884 20043 3936 20052
rect 3884 20009 3893 20043
rect 3893 20009 3927 20043
rect 3927 20009 3936 20043
rect 3884 20000 3936 20009
rect 10692 20000 10744 20052
rect 3976 19932 4028 19984
rect 5724 19975 5776 19984
rect 5724 19941 5733 19975
rect 5733 19941 5767 19975
rect 5767 19941 5776 19975
rect 5724 19932 5776 19941
rect 1492 19796 1544 19848
rect 2044 19796 2096 19848
rect 2596 19796 2648 19848
rect 4528 19796 4580 19848
rect 6552 19864 6604 19916
rect 7288 19864 7340 19916
rect 7564 19864 7616 19916
rect 8116 19864 8168 19916
rect 8392 19864 8444 19916
rect 9588 19864 9640 19916
rect 11612 20000 11664 20052
rect 11980 20000 12032 20052
rect 17960 20000 18012 20052
rect 18052 20000 18104 20052
rect 12164 19932 12216 19984
rect 14464 19932 14516 19984
rect 2780 19728 2832 19780
rect 4252 19728 4304 19780
rect 5632 19796 5684 19848
rect 5908 19796 5960 19848
rect 6644 19796 6696 19848
rect 11888 19864 11940 19916
rect 14372 19864 14424 19916
rect 18144 19932 18196 19984
rect 6736 19728 6788 19780
rect 4344 19703 4396 19712
rect 4344 19669 4353 19703
rect 4353 19669 4387 19703
rect 4387 19669 4396 19703
rect 4344 19660 4396 19669
rect 7288 19771 7340 19780
rect 7288 19737 7297 19771
rect 7297 19737 7331 19771
rect 7331 19737 7340 19771
rect 7288 19728 7340 19737
rect 7472 19728 7524 19780
rect 8208 19728 8260 19780
rect 8392 19771 8444 19780
rect 8392 19737 8401 19771
rect 8401 19737 8435 19771
rect 8435 19737 8444 19771
rect 8392 19728 8444 19737
rect 9404 19728 9456 19780
rect 10324 19771 10376 19780
rect 10324 19737 10342 19771
rect 10342 19737 10376 19771
rect 10324 19728 10376 19737
rect 11152 19771 11204 19780
rect 11152 19737 11186 19771
rect 11186 19737 11204 19771
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 13452 19839 13504 19848
rect 12532 19796 12584 19805
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 11152 19728 11204 19737
rect 16028 19796 16080 19848
rect 15108 19728 15160 19780
rect 16304 19796 16356 19848
rect 18052 19864 18104 19916
rect 18144 19839 18196 19848
rect 7380 19703 7432 19712
rect 7380 19669 7389 19703
rect 7389 19669 7423 19703
rect 7423 19669 7432 19703
rect 7380 19660 7432 19669
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 8484 19660 8536 19712
rect 9496 19660 9548 19712
rect 9864 19660 9916 19712
rect 10876 19660 10928 19712
rect 11520 19660 11572 19712
rect 12624 19660 12676 19712
rect 14280 19660 14332 19712
rect 14464 19660 14516 19712
rect 17040 19728 17092 19780
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 20720 19796 20772 19848
rect 20904 19796 20956 19848
rect 19800 19771 19852 19780
rect 16764 19660 16816 19712
rect 19800 19737 19834 19771
rect 19834 19737 19852 19771
rect 19800 19728 19852 19737
rect 19984 19728 20036 19780
rect 19708 19660 19760 19712
rect 20996 19660 21048 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 4068 19456 4120 19508
rect 5816 19456 5868 19508
rect 6644 19456 6696 19508
rect 4160 19431 4212 19440
rect 4160 19397 4169 19431
rect 4169 19397 4203 19431
rect 4203 19397 4212 19431
rect 4160 19388 4212 19397
rect 7012 19456 7064 19508
rect 7196 19456 7248 19508
rect 8116 19499 8168 19508
rect 8116 19465 8125 19499
rect 8125 19465 8159 19499
rect 8159 19465 8168 19499
rect 8116 19456 8168 19465
rect 9312 19456 9364 19508
rect 9496 19456 9548 19508
rect 11336 19456 11388 19508
rect 11888 19456 11940 19508
rect 12164 19499 12216 19508
rect 12164 19465 12173 19499
rect 12173 19465 12207 19499
rect 12207 19465 12216 19499
rect 12164 19456 12216 19465
rect 14556 19456 14608 19508
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 14832 19456 14884 19508
rect 16304 19456 16356 19508
rect 940 19252 992 19304
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 5540 19320 5592 19372
rect 5724 19320 5776 19372
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 7104 19388 7156 19440
rect 3148 19184 3200 19236
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 4344 19184 4396 19236
rect 3884 19116 3936 19168
rect 4160 19116 4212 19168
rect 5172 19116 5224 19168
rect 10324 19388 10376 19440
rect 12992 19388 13044 19440
rect 13728 19388 13780 19440
rect 18788 19456 18840 19508
rect 20444 19456 20496 19508
rect 19708 19388 19760 19440
rect 7748 19320 7800 19372
rect 9588 19320 9640 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 8392 19252 8444 19304
rect 7472 19116 7524 19168
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 8576 19116 8628 19168
rect 10968 19252 11020 19304
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 13820 19320 13872 19372
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 16856 19320 16908 19372
rect 20168 19320 20220 19372
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 10784 19184 10836 19236
rect 13268 19184 13320 19236
rect 12992 19159 13044 19168
rect 12992 19125 13001 19159
rect 13001 19125 13035 19159
rect 13035 19125 13044 19159
rect 12992 19116 13044 19125
rect 13728 19116 13780 19168
rect 16580 19116 16632 19168
rect 18236 19116 18288 19168
rect 18604 19116 18656 19168
rect 21548 19116 21600 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 2044 18912 2096 18964
rect 4804 18912 4856 18964
rect 8208 18912 8260 18964
rect 9220 18912 9272 18964
rect 9588 18912 9640 18964
rect 13452 18912 13504 18964
rect 2596 18844 2648 18896
rect 5080 18844 5132 18896
rect 6736 18887 6788 18896
rect 6736 18853 6745 18887
rect 6745 18853 6779 18887
rect 6779 18853 6788 18887
rect 6736 18844 6788 18853
rect 6920 18844 6972 18896
rect 7380 18844 7432 18896
rect 8944 18887 8996 18896
rect 8944 18853 8953 18887
rect 8953 18853 8987 18887
rect 8987 18853 8996 18887
rect 8944 18844 8996 18853
rect 12808 18844 12860 18896
rect 15200 18912 15252 18964
rect 17960 18912 18012 18964
rect 21364 18912 21416 18964
rect 4528 18776 4580 18828
rect 7288 18776 7340 18828
rect 4436 18751 4488 18760
rect 4436 18717 4445 18751
rect 4445 18717 4479 18751
rect 4479 18717 4488 18751
rect 4436 18708 4488 18717
rect 4160 18640 4212 18692
rect 5264 18640 5316 18692
rect 6644 18708 6696 18760
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 10692 18708 10744 18760
rect 12532 18751 12584 18760
rect 7104 18640 7156 18692
rect 8944 18640 8996 18692
rect 3884 18572 3936 18624
rect 5632 18572 5684 18624
rect 6828 18572 6880 18624
rect 7288 18572 7340 18624
rect 7656 18572 7708 18624
rect 12532 18717 12550 18751
rect 12550 18717 12584 18751
rect 12532 18708 12584 18717
rect 13084 18776 13136 18828
rect 16856 18819 16908 18828
rect 13544 18708 13596 18760
rect 13636 18708 13688 18760
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 14372 18708 14424 18760
rect 12992 18640 13044 18692
rect 15108 18708 15160 18760
rect 15752 18640 15804 18692
rect 16856 18785 16865 18819
rect 16865 18785 16899 18819
rect 16899 18785 16908 18819
rect 16856 18776 16908 18785
rect 20720 18776 20772 18828
rect 21272 18776 21324 18828
rect 18236 18708 18288 18760
rect 18696 18708 18748 18760
rect 19800 18640 19852 18692
rect 20444 18640 20496 18692
rect 20904 18708 20956 18760
rect 22560 18640 22612 18692
rect 12256 18572 12308 18624
rect 13728 18572 13780 18624
rect 15844 18615 15896 18624
rect 15844 18581 15853 18615
rect 15853 18581 15887 18615
rect 15887 18581 15896 18615
rect 15844 18572 15896 18581
rect 17960 18572 18012 18624
rect 18420 18572 18472 18624
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 19708 18572 19760 18624
rect 21456 18572 21508 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 940 18368 992 18420
rect 1492 18368 1544 18420
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 4160 18368 4212 18420
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 7012 18411 7064 18420
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 10784 18368 10836 18420
rect 12440 18368 12492 18420
rect 12624 18368 12676 18420
rect 13360 18368 13412 18420
rect 13544 18368 13596 18420
rect 15568 18368 15620 18420
rect 16856 18368 16908 18420
rect 16948 18368 17000 18420
rect 17132 18368 17184 18420
rect 22192 18368 22244 18420
rect 3240 18300 3292 18352
rect 4988 18300 5040 18352
rect 9220 18300 9272 18352
rect 5908 18232 5960 18284
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 7380 18232 7432 18284
rect 8024 18232 8076 18284
rect 9772 18232 9824 18284
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 7564 18164 7616 18216
rect 8944 18164 8996 18216
rect 5540 18096 5592 18148
rect 5724 18096 5776 18148
rect 7012 18028 7064 18080
rect 11152 18096 11204 18148
rect 10600 18028 10652 18080
rect 10968 18028 11020 18080
rect 12716 18300 12768 18352
rect 12256 18232 12308 18284
rect 13360 18232 13412 18284
rect 14188 18232 14240 18284
rect 14372 18232 14424 18284
rect 17868 18300 17920 18352
rect 20996 18300 21048 18352
rect 21548 18300 21600 18352
rect 15844 18164 15896 18216
rect 18972 18232 19024 18284
rect 21272 18232 21324 18284
rect 15568 18096 15620 18148
rect 16304 18096 16356 18148
rect 18328 18096 18380 18148
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 18696 18028 18748 18080
rect 18972 18028 19024 18080
rect 21088 18028 21140 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 4160 17867 4212 17876
rect 4160 17833 4169 17867
rect 4169 17833 4203 17867
rect 4203 17833 4212 17867
rect 4160 17824 4212 17833
rect 5356 17824 5408 17876
rect 7104 17824 7156 17876
rect 12164 17824 12216 17876
rect 12440 17824 12492 17876
rect 13820 17824 13872 17876
rect 14832 17867 14884 17876
rect 6000 17756 6052 17808
rect 7840 17756 7892 17808
rect 8024 17756 8076 17808
rect 9496 17756 9548 17808
rect 10876 17756 10928 17808
rect 11796 17756 11848 17808
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 17224 17824 17276 17876
rect 17408 17824 17460 17876
rect 22468 17824 22520 17876
rect 2044 17731 2096 17740
rect 2044 17697 2053 17731
rect 2053 17697 2087 17731
rect 2087 17697 2096 17731
rect 2044 17688 2096 17697
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 4160 17484 4212 17536
rect 5448 17484 5500 17536
rect 5908 17484 5960 17536
rect 7380 17688 7432 17740
rect 15016 17688 15068 17740
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 9312 17620 9364 17672
rect 11888 17620 11940 17672
rect 14464 17620 14516 17672
rect 14740 17620 14792 17672
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 17868 17620 17920 17672
rect 18880 17620 18932 17672
rect 21272 17620 21324 17672
rect 7288 17552 7340 17604
rect 10784 17552 10836 17604
rect 12164 17552 12216 17604
rect 15200 17552 15252 17604
rect 8576 17484 8628 17536
rect 9312 17484 9364 17536
rect 9496 17484 9548 17536
rect 10876 17484 10928 17536
rect 10968 17484 11020 17536
rect 12440 17484 12492 17536
rect 12532 17484 12584 17536
rect 15568 17552 15620 17604
rect 16396 17552 16448 17604
rect 17132 17552 17184 17604
rect 18052 17552 18104 17604
rect 20996 17552 21048 17604
rect 21088 17595 21140 17604
rect 21088 17561 21128 17595
rect 21128 17561 21140 17595
rect 21088 17552 21140 17561
rect 22100 17552 22152 17604
rect 15476 17484 15528 17536
rect 17224 17484 17276 17536
rect 17316 17484 17368 17536
rect 18604 17484 18656 17536
rect 19248 17484 19300 17536
rect 19524 17484 19576 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 4252 17280 4304 17332
rect 7748 17280 7800 17332
rect 8208 17280 8260 17332
rect 12164 17280 12216 17332
rect 8576 17212 8628 17264
rect 4896 17144 4948 17196
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 9864 17144 9916 17196
rect 10140 17187 10192 17196
rect 14740 17212 14792 17264
rect 15752 17212 15804 17264
rect 10140 17153 10158 17187
rect 10158 17153 10192 17187
rect 10140 17144 10192 17153
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 5540 17076 5592 17128
rect 9312 17076 9364 17128
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15568 17187 15620 17196
rect 15108 17144 15160 17153
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 17316 17280 17368 17332
rect 18420 17323 18472 17332
rect 17408 17212 17460 17264
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 20812 17212 20864 17264
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 17316 17144 17368 17196
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 20352 17144 20404 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 21640 17144 21692 17196
rect 15292 17076 15344 17128
rect 5356 17008 5408 17060
rect 8576 17008 8628 17060
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 10232 16940 10284 16992
rect 12440 16940 12492 16992
rect 18512 17076 18564 17128
rect 21272 17076 21324 17128
rect 19064 17008 19116 17060
rect 17960 16940 18012 16992
rect 18512 16940 18564 16992
rect 20628 16940 20680 16992
rect 21364 16940 21416 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 7196 16736 7248 16788
rect 4896 16600 4948 16652
rect 6828 16600 6880 16652
rect 13544 16736 13596 16788
rect 16672 16736 16724 16788
rect 15292 16668 15344 16720
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 8576 16600 8628 16652
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 12348 16600 12400 16652
rect 13452 16600 13504 16652
rect 15752 16643 15804 16652
rect 5540 16464 5592 16516
rect 8944 16464 8996 16516
rect 13084 16532 13136 16584
rect 4160 16396 4212 16448
rect 5724 16396 5776 16448
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 8116 16396 8168 16448
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 15200 16532 15252 16584
rect 13360 16464 13412 16516
rect 16212 16464 16264 16516
rect 19524 16736 19576 16788
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 17592 16532 17644 16584
rect 20812 16532 20864 16584
rect 18512 16464 18564 16516
rect 12808 16396 12860 16405
rect 15936 16396 15988 16448
rect 17684 16396 17736 16448
rect 20352 16396 20404 16448
rect 21456 16396 21508 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 5816 16192 5868 16244
rect 7012 16192 7064 16244
rect 9128 16192 9180 16244
rect 15660 16192 15712 16244
rect 4896 16056 4948 16108
rect 4620 15988 4672 16040
rect 5816 16056 5868 16108
rect 6828 16056 6880 16108
rect 8576 16124 8628 16176
rect 10232 16124 10284 16176
rect 13636 16124 13688 16176
rect 16856 16192 16908 16244
rect 7012 15988 7064 16040
rect 7288 15988 7340 16040
rect 10692 16056 10744 16108
rect 12716 16056 12768 16108
rect 13452 16056 13504 16108
rect 13820 16099 13872 16108
rect 13820 16065 13854 16099
rect 13854 16065 13872 16099
rect 13820 16056 13872 16065
rect 7196 15920 7248 15972
rect 16488 16056 16540 16108
rect 17868 16124 17920 16176
rect 16948 16099 17000 16108
rect 16948 16065 16982 16099
rect 16982 16065 17000 16099
rect 16580 15988 16632 16040
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 6368 15852 6420 15904
rect 7932 15852 7984 15904
rect 8300 15852 8352 15904
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 9956 15852 10008 15904
rect 10692 15852 10744 15904
rect 11704 15852 11756 15904
rect 11980 15852 12032 15904
rect 12624 15852 12676 15904
rect 15752 15920 15804 15972
rect 16948 16056 17000 16065
rect 20076 16124 20128 16176
rect 17684 15988 17736 16040
rect 19892 16056 19944 16108
rect 21180 16056 21232 16108
rect 19524 15920 19576 15972
rect 17316 15852 17368 15904
rect 19800 15852 19852 15904
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21364 15852 21416 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 7012 15648 7064 15700
rect 7104 15580 7156 15632
rect 8576 15648 8628 15700
rect 9036 15648 9088 15700
rect 10048 15648 10100 15700
rect 8208 15580 8260 15632
rect 9772 15623 9824 15632
rect 9772 15589 9781 15623
rect 9781 15589 9815 15623
rect 9815 15589 9824 15623
rect 9772 15580 9824 15589
rect 13544 15648 13596 15700
rect 14372 15648 14424 15700
rect 16488 15648 16540 15700
rect 17776 15648 17828 15700
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 18604 15648 18656 15700
rect 19616 15691 19668 15700
rect 19616 15657 19625 15691
rect 19625 15657 19659 15691
rect 19659 15657 19668 15691
rect 19616 15648 19668 15657
rect 19984 15580 20036 15632
rect 5724 15444 5776 15496
rect 6552 15444 6604 15496
rect 11704 15512 11756 15564
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 15752 15512 15804 15564
rect 5080 15376 5132 15428
rect 11980 15444 12032 15496
rect 6828 15376 6880 15428
rect 8116 15376 8168 15428
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 5448 15308 5500 15360
rect 5540 15308 5592 15360
rect 6368 15308 6420 15360
rect 9220 15376 9272 15428
rect 11704 15376 11756 15428
rect 10416 15308 10468 15360
rect 18604 15444 18656 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 19064 15444 19116 15496
rect 21272 15444 21324 15496
rect 14924 15376 14976 15428
rect 15660 15376 15712 15428
rect 16580 15376 16632 15428
rect 17776 15376 17828 15428
rect 13268 15308 13320 15360
rect 13820 15308 13872 15360
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 14740 15308 14792 15360
rect 16396 15308 16448 15360
rect 20168 15308 20220 15360
rect 21088 15419 21140 15428
rect 21088 15385 21106 15419
rect 21106 15385 21140 15419
rect 21088 15376 21140 15385
rect 22376 15308 22428 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 4804 15104 4856 15156
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 6644 15104 6696 15156
rect 7104 15104 7156 15156
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9036 15104 9088 15113
rect 4528 15036 4580 15088
rect 7564 14968 7616 15020
rect 7932 15036 7984 15088
rect 9588 15104 9640 15156
rect 7380 14900 7432 14952
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5448 14764 5500 14816
rect 8576 14875 8628 14884
rect 8576 14841 8585 14875
rect 8585 14841 8619 14875
rect 8619 14841 8628 14875
rect 8576 14832 8628 14841
rect 9496 14900 9548 14952
rect 10968 15036 11020 15088
rect 11704 15104 11756 15156
rect 11980 15104 12032 15156
rect 14740 15104 14792 15156
rect 14924 15147 14976 15156
rect 14924 15113 14933 15147
rect 14933 15113 14967 15147
rect 14967 15113 14976 15147
rect 14924 15104 14976 15113
rect 16396 15104 16448 15156
rect 17224 15104 17276 15156
rect 18144 15104 18196 15156
rect 18236 15104 18288 15156
rect 19984 15104 20036 15156
rect 12164 15036 12216 15088
rect 13728 15036 13780 15088
rect 15752 15036 15804 15088
rect 16120 15036 16172 15088
rect 9956 15011 10008 15020
rect 9956 14977 9979 15011
rect 9979 14977 10008 15011
rect 9956 14968 10008 14977
rect 10324 14968 10376 15020
rect 13360 14968 13412 15020
rect 13544 14968 13596 15020
rect 16396 14968 16448 15020
rect 18328 15036 18380 15088
rect 19524 15036 19576 15088
rect 17684 14968 17736 15020
rect 18144 14968 18196 15020
rect 11888 14900 11940 14952
rect 14740 14900 14792 14952
rect 19064 14968 19116 15020
rect 19800 14968 19852 15020
rect 12072 14832 12124 14884
rect 12164 14832 12216 14884
rect 12716 14832 12768 14884
rect 13820 14832 13872 14884
rect 11704 14764 11756 14816
rect 14464 14764 14516 14816
rect 17040 14832 17092 14884
rect 17224 14764 17276 14816
rect 19524 14764 19576 14816
rect 21088 14807 21140 14816
rect 21088 14773 21097 14807
rect 21097 14773 21131 14807
rect 21131 14773 21140 14807
rect 21088 14764 21140 14773
rect 22468 14764 22520 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 6920 14603 6972 14612
rect 6920 14569 6929 14603
rect 6929 14569 6963 14603
rect 6963 14569 6972 14603
rect 6920 14560 6972 14569
rect 8576 14560 8628 14612
rect 10324 14560 10376 14612
rect 9588 14492 9640 14544
rect 4896 14424 4948 14476
rect 5264 14424 5316 14476
rect 3976 14356 4028 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4712 14356 4764 14408
rect 4068 14288 4120 14340
rect 11980 14560 12032 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 13268 14535 13320 14544
rect 13268 14501 13277 14535
rect 13277 14501 13311 14535
rect 13311 14501 13320 14535
rect 13268 14492 13320 14501
rect 14832 14560 14884 14612
rect 17960 14560 18012 14612
rect 16120 14424 16172 14476
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 7012 14220 7064 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 9956 14288 10008 14340
rect 12348 14288 12400 14340
rect 14832 14288 14884 14340
rect 12532 14220 12584 14272
rect 12624 14220 12676 14272
rect 12900 14220 12952 14272
rect 15108 14220 15160 14272
rect 15936 14220 15988 14272
rect 16948 14288 17000 14340
rect 19524 14356 19576 14408
rect 19984 14356 20036 14408
rect 21272 14356 21324 14408
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 20996 14288 21048 14340
rect 21548 14288 21600 14340
rect 19248 14220 19300 14272
rect 19800 14220 19852 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 4344 14016 4396 14068
rect 4988 14016 5040 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 10968 14059 11020 14068
rect 10968 14025 10977 14059
rect 10977 14025 11011 14059
rect 11011 14025 11020 14059
rect 10968 14016 11020 14025
rect 11980 14059 12032 14068
rect 11980 14025 11989 14059
rect 11989 14025 12023 14059
rect 12023 14025 12032 14059
rect 11980 14016 12032 14025
rect 13636 14016 13688 14068
rect 15936 14016 15988 14068
rect 16120 14016 16172 14068
rect 18328 14016 18380 14068
rect 4620 13948 4672 14000
rect 5448 13948 5500 14000
rect 11704 13948 11756 14000
rect 12532 13948 12584 14000
rect 12992 13948 13044 14000
rect 13544 13948 13596 14000
rect 5264 13880 5316 13932
rect 10048 13880 10100 13932
rect 10324 13923 10376 13932
rect 10324 13889 10342 13923
rect 10342 13889 10376 13923
rect 10324 13880 10376 13889
rect 10968 13880 11020 13932
rect 11980 13880 12032 13932
rect 4068 13812 4120 13864
rect 6552 13812 6604 13864
rect 11244 13812 11296 13864
rect 13820 13880 13872 13932
rect 17408 13948 17460 14000
rect 17868 13948 17920 14000
rect 20628 14016 20680 14068
rect 20812 14016 20864 14068
rect 21088 14016 21140 14068
rect 15568 13880 15620 13932
rect 16120 13880 16172 13932
rect 9312 13744 9364 13796
rect 18972 13880 19024 13932
rect 19984 13880 20036 13932
rect 21364 13923 21416 13932
rect 21364 13889 21373 13923
rect 21373 13889 21407 13923
rect 21407 13889 21416 13923
rect 21364 13880 21416 13889
rect 22100 13812 22152 13864
rect 5448 13676 5500 13728
rect 9128 13676 9180 13728
rect 9864 13676 9916 13728
rect 10416 13676 10468 13728
rect 13636 13676 13688 13728
rect 14740 13676 14792 13728
rect 15292 13676 15344 13728
rect 16212 13676 16264 13728
rect 19984 13719 20036 13728
rect 19984 13685 19993 13719
rect 19993 13685 20027 13719
rect 20027 13685 20036 13719
rect 19984 13676 20036 13685
rect 21088 13676 21140 13728
rect 22008 13676 22060 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 6828 13472 6880 13524
rect 10784 13472 10836 13524
rect 11704 13472 11756 13524
rect 15292 13472 15344 13524
rect 16028 13472 16080 13524
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 5172 13336 5224 13388
rect 9036 13311 9088 13320
rect 9036 13277 9045 13311
rect 9045 13277 9079 13311
rect 9079 13277 9088 13311
rect 9036 13268 9088 13277
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 16120 13404 16172 13456
rect 19064 13472 19116 13524
rect 18420 13404 18472 13456
rect 20260 13472 20312 13524
rect 21364 13472 21416 13524
rect 21272 13336 21324 13388
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 5724 13132 5776 13141
rect 7656 13200 7708 13252
rect 9312 13243 9364 13252
rect 9312 13209 9346 13243
rect 9346 13209 9364 13243
rect 11980 13268 12032 13320
rect 9312 13200 9364 13209
rect 12624 13200 12676 13252
rect 7380 13132 7432 13184
rect 9864 13132 9916 13184
rect 9956 13132 10008 13184
rect 11980 13132 12032 13184
rect 12164 13132 12216 13184
rect 16764 13268 16816 13320
rect 17684 13268 17736 13320
rect 20536 13268 20588 13320
rect 20996 13268 21048 13320
rect 14740 13200 14792 13252
rect 17868 13200 17920 13252
rect 19984 13200 20036 13252
rect 20260 13200 20312 13252
rect 14464 13132 14516 13184
rect 15568 13132 15620 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 5724 12928 5776 12980
rect 10140 12928 10192 12980
rect 10508 12928 10560 12980
rect 5540 12860 5592 12912
rect 6552 12792 6604 12844
rect 9036 12860 9088 12912
rect 11612 12903 11664 12912
rect 9220 12792 9272 12844
rect 11612 12869 11621 12903
rect 11621 12869 11655 12903
rect 11655 12869 11664 12903
rect 11612 12860 11664 12869
rect 13728 12860 13780 12912
rect 5448 12724 5500 12776
rect 12072 12792 12124 12844
rect 5724 12699 5776 12708
rect 5724 12665 5733 12699
rect 5733 12665 5767 12699
rect 5767 12665 5776 12699
rect 5724 12656 5776 12665
rect 11980 12724 12032 12776
rect 8484 12588 8536 12640
rect 9956 12588 10008 12640
rect 10048 12588 10100 12640
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 14464 12724 14516 12776
rect 16120 12928 16172 12980
rect 14740 12860 14792 12912
rect 18144 12860 18196 12912
rect 19064 12860 19116 12912
rect 20628 12860 20680 12912
rect 22928 12860 22980 12912
rect 15384 12792 15436 12844
rect 16120 12792 16172 12844
rect 18236 12792 18288 12844
rect 18420 12792 18472 12844
rect 19800 12792 19852 12844
rect 21272 12792 21324 12844
rect 20168 12656 20220 12708
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 6552 12316 6604 12368
rect 7840 12384 7892 12436
rect 7932 12384 7984 12436
rect 8300 12384 8352 12436
rect 10324 12384 10376 12436
rect 8208 12316 8260 12368
rect 8484 12316 8536 12368
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 13268 12316 13320 12368
rect 13544 12316 13596 12368
rect 14740 12384 14792 12436
rect 16120 12384 16172 12436
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10508 12248 10560 12300
rect 11152 12248 11204 12300
rect 10600 12180 10652 12232
rect 15568 12248 15620 12300
rect 16120 12248 16172 12300
rect 18420 12384 18472 12436
rect 19524 12427 19576 12436
rect 16856 12223 16908 12232
rect 6000 12044 6052 12096
rect 7380 12044 7432 12096
rect 9864 12112 9916 12164
rect 10784 12112 10836 12164
rect 16856 12189 16874 12223
rect 16874 12189 16908 12223
rect 16856 12180 16908 12189
rect 11612 12112 11664 12164
rect 12164 12112 12216 12164
rect 13176 12112 13228 12164
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 10048 12044 10100 12096
rect 11060 12044 11112 12096
rect 11152 12044 11204 12096
rect 11980 12044 12032 12096
rect 12532 12044 12584 12096
rect 14740 12044 14792 12096
rect 15108 12044 15160 12096
rect 16120 12044 16172 12096
rect 21272 12180 21324 12232
rect 18420 12112 18472 12164
rect 22376 12112 22428 12164
rect 17960 12044 18012 12096
rect 18328 12044 18380 12096
rect 18972 12044 19024 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 6736 11840 6788 11892
rect 7472 11840 7524 11892
rect 7748 11840 7800 11892
rect 8024 11840 8076 11892
rect 5540 11772 5592 11824
rect 11520 11840 11572 11892
rect 12164 11840 12216 11892
rect 12900 11883 12952 11892
rect 12900 11849 12909 11883
rect 12909 11849 12943 11883
rect 12943 11849 12952 11883
rect 12900 11840 12952 11849
rect 14372 11883 14424 11892
rect 14372 11849 14381 11883
rect 14381 11849 14415 11883
rect 14415 11849 14424 11883
rect 14372 11840 14424 11849
rect 14648 11840 14700 11892
rect 15292 11840 15344 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 15844 11840 15896 11892
rect 17684 11883 17736 11892
rect 17684 11849 17693 11883
rect 17693 11849 17727 11883
rect 17727 11849 17736 11883
rect 17684 11840 17736 11849
rect 18052 11840 18104 11892
rect 18236 11840 18288 11892
rect 19340 11840 19392 11892
rect 21364 11840 21416 11892
rect 7840 11704 7892 11756
rect 8024 11704 8076 11756
rect 9864 11704 9916 11756
rect 10324 11747 10376 11756
rect 10324 11713 10353 11747
rect 10353 11713 10376 11747
rect 10324 11704 10376 11713
rect 10784 11704 10836 11756
rect 4528 11568 4580 11620
rect 7196 11636 7248 11688
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8392 11636 8444 11688
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 6920 11500 6972 11552
rect 9312 11500 9364 11552
rect 11060 11704 11112 11756
rect 11428 11704 11480 11756
rect 11980 11704 12032 11756
rect 14372 11704 14424 11756
rect 15200 11704 15252 11756
rect 16396 11704 16448 11756
rect 17132 11704 17184 11756
rect 17500 11747 17552 11756
rect 12164 11636 12216 11688
rect 11060 11568 11112 11620
rect 13728 11636 13780 11688
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 17960 11747 18012 11756
rect 17960 11713 17969 11747
rect 17969 11713 18003 11747
rect 18003 11713 18012 11747
rect 18236 11747 18288 11756
rect 17960 11704 18012 11713
rect 18236 11713 18270 11747
rect 18270 11713 18288 11747
rect 18236 11704 18288 11713
rect 20168 11772 20220 11824
rect 21272 11704 21324 11756
rect 9680 11500 9732 11552
rect 10876 11500 10928 11552
rect 11612 11500 11664 11552
rect 12440 11500 12492 11552
rect 14188 11568 14240 11620
rect 15384 11568 15436 11620
rect 15568 11568 15620 11620
rect 17132 11568 17184 11620
rect 13452 11500 13504 11552
rect 15016 11500 15068 11552
rect 15292 11500 15344 11552
rect 16212 11500 16264 11552
rect 17776 11636 17828 11688
rect 17776 11500 17828 11552
rect 18236 11500 18288 11552
rect 19984 11568 20036 11620
rect 19800 11500 19852 11552
rect 22744 11568 22796 11620
rect 21548 11500 21600 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 7288 11296 7340 11348
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 8024 11228 8076 11280
rect 6000 11160 6052 11212
rect 11612 11296 11664 11348
rect 8208 11160 8260 11212
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7380 11092 7432 11144
rect 7564 11092 7616 11144
rect 7656 11092 7708 11144
rect 9036 11092 9088 11144
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 11520 11160 11572 11212
rect 13452 11296 13504 11348
rect 14832 11296 14884 11348
rect 15200 11339 15252 11348
rect 15200 11305 15209 11339
rect 15209 11305 15243 11339
rect 15243 11305 15252 11339
rect 15200 11296 15252 11305
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 11980 11228 12032 11280
rect 12164 11271 12216 11280
rect 12164 11237 12173 11271
rect 12173 11237 12207 11271
rect 12207 11237 12216 11271
rect 12164 11228 12216 11237
rect 12624 11228 12676 11280
rect 17960 11296 18012 11348
rect 15752 11203 15804 11212
rect 10876 11092 10928 11101
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 6920 11024 6972 11076
rect 7380 10956 7432 11008
rect 8024 10956 8076 11008
rect 9128 10956 9180 11008
rect 9404 10956 9456 11008
rect 11428 11024 11480 11076
rect 12624 11092 12676 11144
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 18328 11228 18380 11280
rect 21088 11228 21140 11280
rect 17960 11092 18012 11144
rect 11520 10956 11572 11008
rect 15844 11024 15896 11076
rect 12164 10956 12216 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 13452 10999 13504 11008
rect 12440 10956 12492 10965
rect 13452 10965 13461 10999
rect 13461 10965 13495 10999
rect 13495 10965 13504 10999
rect 13452 10956 13504 10965
rect 14832 10956 14884 11008
rect 15752 10956 15804 11008
rect 16304 10956 16356 11008
rect 17684 10999 17736 11008
rect 17684 10965 17693 10999
rect 17693 10965 17727 10999
rect 17727 10965 17736 10999
rect 17684 10956 17736 10965
rect 19524 11092 19576 11144
rect 20444 11160 20496 11212
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 20996 11092 21048 11144
rect 18696 11024 18748 11076
rect 20352 11024 20404 11076
rect 21364 11024 21416 11076
rect 22560 11024 22612 11076
rect 18328 10999 18380 11008
rect 18328 10965 18337 10999
rect 18337 10965 18371 10999
rect 18371 10965 18380 10999
rect 18328 10956 18380 10965
rect 19984 10956 20036 11008
rect 20628 10999 20680 11008
rect 20628 10965 20637 10999
rect 20637 10965 20671 10999
rect 20671 10965 20680 10999
rect 20628 10956 20680 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 5724 10752 5776 10804
rect 6460 10752 6512 10804
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 8576 10752 8628 10804
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 10140 10752 10192 10804
rect 10692 10752 10744 10804
rect 11244 10752 11296 10804
rect 12348 10795 12400 10804
rect 12348 10761 12357 10795
rect 12357 10761 12391 10795
rect 12391 10761 12400 10795
rect 12348 10752 12400 10761
rect 12440 10752 12492 10804
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 7932 10684 7984 10736
rect 10324 10684 10376 10736
rect 10876 10684 10928 10736
rect 11980 10727 12032 10736
rect 11980 10693 11989 10727
rect 11989 10693 12023 10727
rect 12023 10693 12032 10727
rect 11980 10684 12032 10693
rect 13084 10684 13136 10736
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 9680 10616 9732 10668
rect 10416 10616 10468 10668
rect 12348 10616 12400 10668
rect 15292 10684 15344 10736
rect 16212 10684 16264 10736
rect 16948 10752 17000 10804
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 18696 10795 18748 10804
rect 18696 10761 18705 10795
rect 18705 10761 18739 10795
rect 18739 10761 18748 10795
rect 18696 10752 18748 10761
rect 21088 10752 21140 10804
rect 22100 10752 22152 10804
rect 16672 10659 16724 10668
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 7748 10548 7800 10600
rect 9036 10548 9088 10600
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 10968 10548 11020 10600
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 13820 10548 13872 10600
rect 14372 10548 14424 10600
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 16948 10616 17000 10668
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 18696 10616 18748 10668
rect 18972 10616 19024 10668
rect 19984 10684 20036 10736
rect 19800 10616 19852 10668
rect 16120 10523 16172 10532
rect 5724 10412 5776 10464
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 16120 10489 16129 10523
rect 16129 10489 16163 10523
rect 16163 10489 16172 10523
rect 16120 10480 16172 10489
rect 13544 10412 13596 10464
rect 15200 10412 15252 10464
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 19708 10548 19760 10600
rect 20076 10548 20128 10600
rect 18788 10480 18840 10532
rect 20444 10480 20496 10532
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18328 10412 18380 10464
rect 20076 10412 20128 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 5356 10072 5408 10124
rect 6828 10208 6880 10260
rect 5540 10140 5592 10192
rect 6460 10140 6512 10192
rect 10048 10208 10100 10260
rect 13360 10208 13412 10260
rect 9680 10140 9732 10192
rect 10140 10140 10192 10192
rect 14004 10208 14056 10260
rect 14464 10208 14516 10260
rect 14924 10208 14976 10260
rect 15016 10208 15068 10260
rect 16672 10208 16724 10260
rect 17592 10208 17644 10260
rect 20812 10251 20864 10260
rect 20812 10217 20821 10251
rect 20821 10217 20855 10251
rect 20855 10217 20864 10251
rect 20812 10208 20864 10217
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 16948 10140 17000 10192
rect 21364 10140 21416 10192
rect 4988 10004 5040 10056
rect 8300 10072 8352 10124
rect 9312 10072 9364 10124
rect 10508 10072 10560 10124
rect 6460 10004 6512 10056
rect 7840 10004 7892 10056
rect 3884 9936 3936 9988
rect 5172 9936 5224 9988
rect 7748 9979 7800 9988
rect 7748 9945 7757 9979
rect 7757 9945 7791 9979
rect 7791 9945 7800 9979
rect 7748 9936 7800 9945
rect 9772 9936 9824 9988
rect 13636 10072 13688 10124
rect 14372 10072 14424 10124
rect 15200 10072 15252 10124
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 17960 10072 18012 10124
rect 18052 10072 18104 10124
rect 18512 10072 18564 10124
rect 13452 10004 13504 10056
rect 13728 10004 13780 10056
rect 15108 10004 15160 10056
rect 16212 10004 16264 10056
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 15016 9936 15068 9988
rect 18696 10004 18748 10056
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 19616 10004 19668 10056
rect 20628 10072 20680 10124
rect 5264 9868 5316 9920
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6000 9868 6052 9920
rect 7564 9868 7616 9920
rect 9680 9868 9732 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 11888 9868 11940 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13544 9868 13596 9920
rect 14096 9868 14148 9920
rect 15108 9911 15160 9920
rect 15108 9877 15117 9911
rect 15117 9877 15151 9911
rect 15151 9877 15160 9911
rect 15108 9868 15160 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 16304 9868 16356 9920
rect 19156 9936 19208 9988
rect 20812 9936 20864 9988
rect 21088 9936 21140 9988
rect 17040 9868 17092 9920
rect 17592 9868 17644 9920
rect 19616 9868 19668 9920
rect 19708 9868 19760 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 6000 9664 6052 9716
rect 9864 9664 9916 9716
rect 10416 9664 10468 9716
rect 5908 9596 5960 9648
rect 5724 9528 5776 9580
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 4804 9392 4856 9444
rect 5264 9392 5316 9444
rect 6276 9460 6328 9512
rect 7288 9460 7340 9512
rect 7196 9324 7248 9376
rect 8116 9596 8168 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 11244 9596 11296 9648
rect 11704 9596 11756 9648
rect 13912 9664 13964 9716
rect 14648 9664 14700 9716
rect 15108 9664 15160 9716
rect 15568 9664 15620 9716
rect 16672 9664 16724 9716
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 17960 9664 18012 9716
rect 18696 9707 18748 9716
rect 18696 9673 18705 9707
rect 18705 9673 18739 9707
rect 18739 9673 18748 9707
rect 18696 9664 18748 9673
rect 19892 9707 19944 9716
rect 13636 9639 13688 9648
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8300 9460 8352 9512
rect 8392 9392 8444 9444
rect 9220 9528 9272 9580
rect 13636 9605 13645 9639
rect 13645 9605 13679 9639
rect 13679 9605 13688 9639
rect 13636 9596 13688 9605
rect 14096 9596 14148 9648
rect 14464 9596 14516 9648
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 12164 9435 12216 9444
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 9680 9324 9732 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 12900 9460 12952 9512
rect 13268 9528 13320 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 14372 9460 14424 9512
rect 14004 9392 14056 9444
rect 14832 9528 14884 9580
rect 15660 9571 15712 9580
rect 14924 9503 14976 9512
rect 14924 9469 14933 9503
rect 14933 9469 14967 9503
rect 14967 9469 14976 9503
rect 14924 9460 14976 9469
rect 15108 9460 15160 9512
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 14832 9392 14884 9444
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 17132 9392 17184 9444
rect 16120 9324 16172 9376
rect 16672 9324 16724 9376
rect 17040 9324 17092 9376
rect 18972 9596 19024 9648
rect 19892 9673 19901 9707
rect 19901 9673 19935 9707
rect 19935 9673 19944 9707
rect 19892 9664 19944 9673
rect 21088 9664 21140 9716
rect 22100 9664 22152 9716
rect 22284 9664 22336 9716
rect 20260 9596 20312 9648
rect 22560 9596 22612 9648
rect 17960 9392 18012 9444
rect 18420 9392 18472 9444
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 19064 9392 19116 9444
rect 19708 9392 19760 9444
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 20260 9460 20312 9512
rect 21180 9435 21232 9444
rect 21180 9401 21189 9435
rect 21189 9401 21223 9435
rect 21223 9401 21232 9435
rect 21180 9392 21232 9401
rect 19156 9324 19208 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 6644 9120 6696 9172
rect 7104 9120 7156 9172
rect 7288 9120 7340 9172
rect 9312 9120 9364 9172
rect 10508 9120 10560 9172
rect 11980 9120 12032 9172
rect 14372 9120 14424 9172
rect 14924 9120 14976 9172
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 15660 9120 15712 9172
rect 18420 9163 18472 9172
rect 6000 8984 6052 9036
rect 7380 9052 7432 9104
rect 10600 9052 10652 9104
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 4712 8848 4764 8900
rect 7012 8984 7064 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 9588 8984 9640 9036
rect 9864 8984 9916 9036
rect 10140 8984 10192 9036
rect 10508 8984 10560 9036
rect 10784 8984 10836 9036
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 16764 8984 16816 9036
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 7380 8780 7432 8832
rect 9680 8916 9732 8968
rect 17408 9052 17460 9104
rect 10140 8848 10192 8900
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 10048 8780 10100 8832
rect 11704 8848 11756 8900
rect 12716 8848 12768 8900
rect 10416 8780 10468 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 11980 8780 12032 8832
rect 14648 8780 14700 8832
rect 14924 8848 14976 8900
rect 17776 8984 17828 9036
rect 17960 9052 18012 9104
rect 18144 9052 18196 9104
rect 18420 9129 18429 9163
rect 18429 9129 18463 9163
rect 18463 9129 18472 9163
rect 18420 9120 18472 9129
rect 18788 9120 18840 9172
rect 19432 9052 19484 9104
rect 18420 8984 18472 9036
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 20352 9120 20404 9172
rect 20720 9052 20772 9104
rect 17408 8916 17460 8968
rect 19616 8916 19668 8968
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 16948 8780 17000 8832
rect 17500 8780 17552 8832
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 18236 8780 18288 8832
rect 18972 8780 19024 8832
rect 20628 8848 20680 8900
rect 20720 8780 20772 8832
rect 20996 8780 21048 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 7288 8619 7340 8628
rect 7288 8585 7297 8619
rect 7297 8585 7331 8619
rect 7331 8585 7340 8619
rect 7288 8576 7340 8585
rect 7932 8576 7984 8628
rect 9496 8576 9548 8628
rect 9588 8576 9640 8628
rect 10416 8576 10468 8628
rect 8300 8508 8352 8560
rect 8208 8440 8260 8492
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 5264 8372 5316 8381
rect 5540 8372 5592 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7932 8372 7984 8424
rect 9128 8372 9180 8424
rect 6644 8304 6696 8356
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 10232 8440 10284 8492
rect 11704 8576 11756 8628
rect 12256 8619 12308 8628
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 13728 8576 13780 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17408 8619 17460 8628
rect 17040 8576 17092 8585
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17592 8576 17644 8628
rect 18144 8619 18196 8628
rect 14464 8508 14516 8560
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 20628 8619 20680 8628
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 12992 8440 13044 8492
rect 11060 8372 11112 8424
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 15108 8440 15160 8492
rect 17592 8440 17644 8492
rect 14280 8372 14332 8424
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14924 8372 14976 8424
rect 17224 8372 17276 8424
rect 17408 8372 17460 8424
rect 17960 8440 18012 8492
rect 20260 8508 20312 8560
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 21088 8551 21140 8560
rect 21088 8517 21097 8551
rect 21097 8517 21131 8551
rect 21131 8517 21140 8551
rect 21088 8508 21140 8517
rect 19064 8440 19116 8492
rect 18420 8372 18472 8424
rect 7380 8236 7432 8288
rect 8208 8236 8260 8288
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9496 8236 9548 8288
rect 10048 8304 10100 8356
rect 12440 8304 12492 8356
rect 15016 8304 15068 8356
rect 11336 8236 11388 8288
rect 11428 8236 11480 8288
rect 11888 8236 11940 8288
rect 13728 8236 13780 8288
rect 14372 8236 14424 8288
rect 16120 8236 16172 8288
rect 19984 8440 20036 8492
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 21456 8372 21508 8424
rect 19800 8304 19852 8356
rect 22652 8304 22704 8356
rect 19432 8236 19484 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 6736 8032 6788 8084
rect 7748 8032 7800 8084
rect 10048 8075 10100 8084
rect 4988 7964 5040 8016
rect 7932 7964 7984 8016
rect 8208 7964 8260 8016
rect 9312 7964 9364 8016
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10324 8032 10376 8084
rect 12624 8032 12676 8084
rect 12992 8032 13044 8084
rect 5356 7896 5408 7948
rect 6000 7896 6052 7948
rect 6644 7896 6696 7948
rect 9128 7896 9180 7948
rect 11428 7964 11480 8016
rect 14556 8032 14608 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 15752 8032 15804 8084
rect 15936 8032 15988 8084
rect 17592 8032 17644 8084
rect 19892 8075 19944 8084
rect 19892 8041 19901 8075
rect 19901 8041 19935 8075
rect 19935 8041 19944 8075
rect 19892 8032 19944 8041
rect 20260 8032 20312 8084
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 13728 7964 13780 8016
rect 18420 7964 18472 8016
rect 18512 7964 18564 8016
rect 12624 7896 12676 7948
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 5540 7828 5592 7880
rect 11060 7828 11112 7880
rect 11980 7828 12032 7880
rect 12440 7828 12492 7880
rect 16120 7896 16172 7948
rect 16212 7896 16264 7948
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 4620 7692 4672 7744
rect 5172 7692 5224 7744
rect 14280 7760 14332 7812
rect 20076 7871 20128 7880
rect 20076 7837 20085 7871
rect 20085 7837 20119 7871
rect 20119 7837 20128 7871
rect 20076 7828 20128 7837
rect 21640 7964 21692 8016
rect 20720 7828 20772 7880
rect 14556 7760 14608 7812
rect 5908 7692 5960 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 10968 7692 11020 7744
rect 11704 7692 11756 7744
rect 12716 7692 12768 7744
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 15292 7760 15344 7812
rect 14464 7692 14516 7701
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 16120 7692 16172 7744
rect 17132 7760 17184 7812
rect 18236 7760 18288 7812
rect 17408 7692 17460 7744
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 18788 7692 18840 7744
rect 22468 7692 22520 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 5908 7488 5960 7540
rect 7104 7488 7156 7540
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 9220 7488 9272 7540
rect 10600 7488 10652 7540
rect 10692 7488 10744 7540
rect 11888 7488 11940 7540
rect 12348 7488 12400 7540
rect 13452 7488 13504 7540
rect 13636 7488 13688 7540
rect 13820 7488 13872 7540
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 15016 7488 15068 7540
rect 16120 7488 16172 7540
rect 16948 7488 17000 7540
rect 17592 7488 17644 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 18420 7488 18472 7540
rect 6092 7420 6144 7472
rect 6828 7420 6880 7472
rect 9588 7420 9640 7472
rect 11704 7420 11756 7472
rect 14372 7420 14424 7472
rect 15108 7420 15160 7472
rect 18052 7420 18104 7472
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 10232 7352 10284 7404
rect 10784 7352 10836 7404
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12716 7352 12768 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16120 7352 16172 7404
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 4896 7148 4948 7200
rect 5448 7284 5500 7336
rect 9864 7284 9916 7336
rect 11520 7284 11572 7336
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 8300 7216 8352 7268
rect 12348 7216 12400 7268
rect 13268 7327 13320 7336
rect 13268 7293 13277 7327
rect 13277 7293 13311 7327
rect 13311 7293 13320 7327
rect 13452 7327 13504 7336
rect 13268 7284 13320 7293
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 15200 7284 15252 7336
rect 15936 7284 15988 7336
rect 17684 7352 17736 7404
rect 18788 7352 18840 7404
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 18604 7284 18656 7336
rect 19524 7488 19576 7540
rect 20444 7488 20496 7540
rect 20904 7531 20956 7540
rect 20904 7497 20913 7531
rect 20913 7497 20947 7531
rect 20947 7497 20956 7531
rect 20904 7488 20956 7497
rect 18972 7420 19024 7472
rect 19340 7395 19392 7404
rect 9772 7148 9824 7200
rect 10416 7148 10468 7200
rect 11980 7148 12032 7200
rect 12256 7148 12308 7200
rect 12992 7148 13044 7200
rect 14556 7148 14608 7200
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 22284 7352 22336 7404
rect 20720 7148 20772 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 6828 6944 6880 6996
rect 10784 6944 10836 6996
rect 11520 6944 11572 6996
rect 13452 6944 13504 6996
rect 13820 6944 13872 6996
rect 14372 6944 14424 6996
rect 15568 6987 15620 6996
rect 15568 6953 15577 6987
rect 15577 6953 15611 6987
rect 15611 6953 15620 6987
rect 15568 6944 15620 6953
rect 16948 6944 17000 6996
rect 17408 6944 17460 6996
rect 10508 6876 10560 6928
rect 10692 6919 10744 6928
rect 10692 6885 10701 6919
rect 10701 6885 10735 6919
rect 10735 6885 10744 6919
rect 10692 6876 10744 6885
rect 11060 6876 11112 6928
rect 12348 6876 12400 6928
rect 12532 6876 12584 6928
rect 12900 6876 12952 6928
rect 12992 6876 13044 6928
rect 18512 6944 18564 6996
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 6828 6740 6880 6792
rect 10968 6808 11020 6860
rect 14832 6808 14884 6860
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9864 6740 9916 6792
rect 13728 6740 13780 6792
rect 10876 6672 10928 6724
rect 11980 6672 12032 6724
rect 12624 6672 12676 6724
rect 12900 6672 12952 6724
rect 16028 6740 16080 6792
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 17316 6808 17368 6860
rect 17776 6740 17828 6792
rect 19156 6876 19208 6928
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18788 6740 18840 6792
rect 15016 6672 15068 6724
rect 20996 6808 21048 6860
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10784 6604 10836 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 13452 6604 13504 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14832 6604 14884 6656
rect 15844 6604 15896 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18052 6604 18104 6656
rect 18236 6604 18288 6656
rect 19064 6604 19116 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20812 6740 20864 6792
rect 21364 6783 21416 6792
rect 21364 6749 21373 6783
rect 21373 6749 21407 6783
rect 21407 6749 21416 6783
rect 21364 6740 21416 6749
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 7932 6400 7984 6452
rect 11980 6400 12032 6452
rect 13544 6400 13596 6452
rect 17592 6400 17644 6452
rect 17960 6400 18012 6452
rect 19064 6400 19116 6452
rect 20352 6400 20404 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 21088 6443 21140 6452
rect 21088 6409 21097 6443
rect 21097 6409 21131 6443
rect 21131 6409 21140 6443
rect 21088 6400 21140 6409
rect 10600 6332 10652 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 7656 6196 7708 6248
rect 8208 6196 8260 6248
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 1584 6171 1636 6180
rect 1584 6137 1593 6171
rect 1593 6137 1627 6171
rect 1627 6137 1636 6171
rect 1584 6128 1636 6137
rect 12164 6264 12216 6316
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13452 6332 13504 6384
rect 15108 6332 15160 6384
rect 19248 6332 19300 6384
rect 15936 6264 15988 6316
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 18420 6264 18472 6316
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19524 6264 19576 6316
rect 20444 6264 20496 6316
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 10692 6060 10744 6112
rect 12348 6128 12400 6180
rect 12624 6128 12676 6180
rect 12808 6171 12860 6180
rect 12808 6137 12817 6171
rect 12817 6137 12851 6171
rect 12851 6137 12860 6171
rect 12808 6128 12860 6137
rect 12900 6060 12952 6112
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13544 6196 13596 6248
rect 14096 6196 14148 6248
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 16948 6196 17000 6248
rect 14832 6128 14884 6180
rect 17408 6196 17460 6248
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 13820 6060 13872 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 16028 6060 16080 6112
rect 17224 6128 17276 6180
rect 21088 6196 21140 6248
rect 22744 6196 22796 6248
rect 16488 6060 16540 6112
rect 18604 6060 18656 6112
rect 18972 6060 19024 6112
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8668 5856 8720 5908
rect 10140 5856 10192 5908
rect 10692 5856 10744 5908
rect 11244 5856 11296 5908
rect 11704 5856 11756 5908
rect 11980 5856 12032 5908
rect 15936 5899 15988 5908
rect 4068 5788 4120 5840
rect 8208 5720 8260 5772
rect 5080 5652 5132 5704
rect 9496 5652 9548 5704
rect 9680 5652 9732 5704
rect 12808 5788 12860 5840
rect 12900 5831 12952 5840
rect 12900 5797 12909 5831
rect 12909 5797 12943 5831
rect 12943 5797 12952 5831
rect 12900 5788 12952 5797
rect 11152 5720 11204 5772
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 13728 5788 13780 5840
rect 16304 5788 16356 5840
rect 13544 5720 13596 5772
rect 12532 5652 12584 5704
rect 13728 5652 13780 5704
rect 8576 5584 8628 5636
rect 10876 5584 10928 5636
rect 11704 5584 11756 5636
rect 13452 5584 13504 5636
rect 15752 5720 15804 5772
rect 16396 5763 16448 5772
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 17684 5720 17736 5772
rect 15108 5652 15160 5704
rect 4252 5516 4304 5568
rect 8392 5516 8444 5568
rect 9772 5516 9824 5568
rect 11244 5516 11296 5568
rect 17224 5652 17276 5704
rect 18880 5788 18932 5840
rect 19892 5788 19944 5840
rect 20168 5720 20220 5772
rect 18144 5584 18196 5636
rect 18420 5627 18472 5636
rect 18420 5593 18429 5627
rect 18429 5593 18463 5627
rect 18463 5593 18472 5627
rect 18420 5584 18472 5593
rect 19616 5584 19668 5636
rect 20628 5652 20680 5704
rect 21180 5652 21232 5704
rect 20720 5584 20772 5636
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 15568 5516 15620 5568
rect 16120 5516 16172 5568
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20536 5559 20588 5568
rect 20536 5525 20545 5559
rect 20545 5525 20579 5559
rect 20579 5525 20588 5559
rect 20536 5516 20588 5525
rect 20628 5516 20680 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 8668 5312 8720 5364
rect 9680 5312 9732 5364
rect 10048 5244 10100 5296
rect 6736 5040 6788 5092
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10692 5312 10744 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 13820 5312 13872 5364
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 15016 5312 15068 5364
rect 16120 5312 16172 5364
rect 16672 5312 16724 5364
rect 18880 5312 18932 5364
rect 19984 5312 20036 5364
rect 20536 5312 20588 5364
rect 16396 5244 16448 5296
rect 12164 5151 12216 5160
rect 10140 5108 10192 5117
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 13360 5176 13412 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 12992 5108 13044 5160
rect 13268 5151 13320 5160
rect 13268 5117 13277 5151
rect 13277 5117 13311 5151
rect 13311 5117 13320 5151
rect 13268 5108 13320 5117
rect 12256 5040 12308 5092
rect 13820 5040 13872 5092
rect 15200 5108 15252 5160
rect 15384 5108 15436 5160
rect 14280 4972 14332 5024
rect 15200 4972 15252 5024
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16304 5176 16356 5228
rect 16396 5040 16448 5092
rect 16028 4972 16080 5024
rect 19800 5244 19852 5296
rect 20260 5244 20312 5296
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 18144 5040 18196 5092
rect 18972 5151 19024 5160
rect 18972 5117 18981 5151
rect 18981 5117 19015 5151
rect 19015 5117 19024 5151
rect 19800 5151 19852 5160
rect 18972 5108 19024 5117
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 21548 5108 21600 5160
rect 22928 5040 22980 5092
rect 16948 4972 17000 5024
rect 17592 4972 17644 5024
rect 18880 4972 18932 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 9128 4768 9180 4820
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 10784 4768 10836 4820
rect 13452 4768 13504 4820
rect 13544 4768 13596 4820
rect 14280 4768 14332 4820
rect 15108 4700 15160 4752
rect 15936 4768 15988 4820
rect 17592 4768 17644 4820
rect 17684 4768 17736 4820
rect 18788 4768 18840 4820
rect 19524 4700 19576 4752
rect 19800 4700 19852 4752
rect 7932 4632 7984 4684
rect 9404 4564 9456 4616
rect 9680 4632 9732 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 11796 4632 11848 4684
rect 12900 4632 12952 4684
rect 13544 4632 13596 4684
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 15292 4632 15344 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 15844 4632 15896 4684
rect 18328 4675 18380 4684
rect 9312 4496 9364 4548
rect 9496 4428 9548 4480
rect 10968 4564 11020 4616
rect 12716 4564 12768 4616
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 13452 4564 13504 4616
rect 15476 4607 15528 4616
rect 10876 4496 10928 4548
rect 11152 4428 11204 4480
rect 11704 4428 11756 4480
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 16948 4564 17000 4616
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 18972 4632 19024 4684
rect 20628 4632 20680 4684
rect 19156 4564 19208 4616
rect 20720 4564 20772 4616
rect 13820 4428 13872 4480
rect 14188 4428 14240 4480
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 17960 4496 18012 4548
rect 19248 4496 19300 4548
rect 14556 4428 14608 4437
rect 15292 4428 15344 4480
rect 15752 4428 15804 4480
rect 16948 4428 17000 4480
rect 17132 4428 17184 4480
rect 17592 4428 17644 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 11060 4224 11112 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 9404 4156 9456 4208
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 10784 4156 10836 4208
rect 12164 4224 12216 4276
rect 12716 4224 12768 4276
rect 14188 4267 14240 4276
rect 14188 4233 14197 4267
rect 14197 4233 14231 4267
rect 14231 4233 14240 4267
rect 14188 4224 14240 4233
rect 14372 4224 14424 4276
rect 15292 4224 15344 4276
rect 15476 4224 15528 4276
rect 16948 4224 17000 4276
rect 18236 4267 18288 4276
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 9772 4020 9824 4072
rect 10968 4020 11020 4072
rect 11980 4020 12032 4072
rect 12624 4088 12676 4140
rect 13084 4088 13136 4140
rect 14924 4156 14976 4208
rect 16580 4156 16632 4208
rect 18236 4233 18245 4267
rect 18245 4233 18279 4267
rect 18279 4233 18288 4267
rect 18236 4224 18288 4233
rect 18420 4156 18472 4208
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13820 4088 13872 4140
rect 14648 4088 14700 4140
rect 15936 4088 15988 4140
rect 16396 4088 16448 4140
rect 13544 4020 13596 4029
rect 15384 4020 15436 4072
rect 15660 4063 15712 4072
rect 15660 4029 15669 4063
rect 15669 4029 15703 4063
rect 15703 4029 15712 4063
rect 15660 4020 15712 4029
rect 17684 4088 17736 4140
rect 20444 4156 20496 4208
rect 18972 4088 19024 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 20628 4088 20680 4140
rect 20352 4020 20404 4072
rect 12624 3952 12676 4004
rect 14832 3952 14884 4004
rect 17224 3952 17276 4004
rect 17776 3952 17828 4004
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8024 3884 8076 3936
rect 8576 3884 8628 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 15936 3884 15988 3936
rect 16672 3884 16724 3936
rect 17684 3884 17736 3936
rect 19064 3884 19116 3936
rect 22468 3952 22520 4004
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 6828 3680 6880 3732
rect 8208 3612 8260 3664
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 9956 3612 10008 3664
rect 10508 3655 10560 3664
rect 10508 3621 10517 3655
rect 10517 3621 10551 3655
rect 10551 3621 10560 3655
rect 10508 3612 10560 3621
rect 10968 3655 11020 3664
rect 10968 3621 10977 3655
rect 10977 3621 11011 3655
rect 11011 3621 11020 3655
rect 10968 3612 11020 3621
rect 12992 3612 13044 3664
rect 15568 3612 15620 3664
rect 18972 3680 19024 3732
rect 940 3476 992 3528
rect 5724 3476 5776 3528
rect 1492 3408 1544 3460
rect 8300 3408 8352 3460
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 4896 3340 4948 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5908 3340 5960 3392
rect 8392 3340 8444 3392
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 9956 3408 10008 3460
rect 11244 3340 11296 3392
rect 12532 3476 12584 3528
rect 14924 3544 14976 3596
rect 15384 3544 15436 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 18604 3612 18656 3664
rect 18696 3612 18748 3664
rect 19156 3612 19208 3664
rect 21548 3612 21600 3664
rect 17316 3544 17368 3596
rect 16580 3519 16632 3528
rect 12348 3408 12400 3460
rect 12072 3340 12124 3392
rect 12624 3340 12676 3392
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 17408 3476 17460 3528
rect 17960 3544 18012 3596
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20536 3519 20588 3528
rect 14832 3340 14884 3392
rect 15292 3340 15344 3392
rect 15476 3340 15528 3392
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 16304 3340 16356 3392
rect 17316 3340 17368 3392
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 18604 3408 18656 3460
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 20168 3451 20220 3460
rect 20168 3417 20177 3451
rect 20177 3417 20211 3451
rect 20211 3417 20220 3451
rect 20168 3408 20220 3417
rect 18512 3340 18564 3392
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 18788 3340 18840 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 7288 3136 7340 3188
rect 11152 3136 11204 3188
rect 5356 3068 5408 3120
rect 5724 3111 5776 3120
rect 5724 3077 5733 3111
rect 5733 3077 5767 3111
rect 5767 3077 5776 3111
rect 5724 3068 5776 3077
rect 8484 3068 8536 3120
rect 1492 3000 1544 3052
rect 4528 3000 4580 3052
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 8116 3000 8168 3052
rect 9220 3000 9272 3052
rect 9772 3000 9824 3052
rect 10048 3000 10100 3052
rect 11704 3000 11756 3052
rect 13452 3136 13504 3188
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 15292 3179 15344 3188
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 18880 3136 18932 3188
rect 19156 3136 19208 3188
rect 13360 3068 13412 3120
rect 15200 3111 15252 3120
rect 12992 3043 13044 3052
rect 3424 2932 3476 2984
rect 9680 2932 9732 2984
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 15200 3077 15209 3111
rect 15209 3077 15243 3111
rect 15243 3077 15252 3111
rect 15200 3068 15252 3077
rect 15936 3068 15988 3120
rect 17132 3043 17184 3052
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 15568 2932 15620 2984
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 17224 2932 17276 2984
rect 17868 3000 17920 3052
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18512 3000 18564 3052
rect 18880 3000 18932 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 5080 2864 5132 2873
rect 7564 2864 7616 2916
rect 10508 2864 10560 2916
rect 11152 2907 11204 2916
rect 11152 2873 11161 2907
rect 11161 2873 11195 2907
rect 11195 2873 11204 2907
rect 11152 2864 11204 2873
rect 11244 2864 11296 2916
rect 15660 2864 15712 2916
rect 16212 2864 16264 2916
rect 2044 2796 2096 2848
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 3148 2839 3200 2848
rect 2780 2796 2832 2805
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 6552 2796 6604 2848
rect 7012 2796 7064 2848
rect 8484 2796 8536 2848
rect 12348 2796 12400 2848
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 13360 2796 13412 2848
rect 15200 2796 15252 2848
rect 16672 2839 16724 2848
rect 16672 2805 16681 2839
rect 16681 2805 16715 2839
rect 16715 2805 16724 2839
rect 16672 2796 16724 2805
rect 17224 2796 17276 2848
rect 18788 2864 18840 2916
rect 21364 2864 21416 2916
rect 18052 2796 18104 2848
rect 20812 2796 20864 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 5724 2592 5776 2644
rect 7656 2592 7708 2644
rect 7932 2592 7984 2644
rect 10232 2592 10284 2644
rect 14556 2592 14608 2644
rect 14648 2592 14700 2644
rect 4620 2499 4672 2508
rect 388 2388 440 2440
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2780 2388 2832 2440
rect 4252 2388 4304 2440
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 5632 2456 5684 2508
rect 9312 2456 9364 2508
rect 6000 2388 6052 2440
rect 7012 2388 7064 2440
rect 8484 2388 8536 2440
rect 8668 2388 8720 2440
rect 2044 2320 2096 2372
rect 3148 2320 3200 2372
rect 5908 2363 5960 2372
rect 5908 2329 5917 2363
rect 5917 2329 5951 2363
rect 5951 2329 5960 2363
rect 5908 2320 5960 2329
rect 6552 2320 6604 2372
rect 7564 2320 7616 2372
rect 8300 2363 8352 2372
rect 8300 2329 8309 2363
rect 8309 2329 8343 2363
rect 8343 2329 8352 2363
rect 8300 2320 8352 2329
rect 10416 2524 10468 2576
rect 13636 2524 13688 2576
rect 14188 2524 14240 2576
rect 15292 2524 15344 2576
rect 16028 2524 16080 2576
rect 10876 2456 10928 2508
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 11520 2320 11572 2372
rect 6736 2252 6788 2304
rect 12808 2456 12860 2508
rect 12900 2456 12952 2508
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 12716 2388 12768 2440
rect 13360 2388 13412 2440
rect 15108 2388 15160 2440
rect 16672 2431 16724 2440
rect 12348 2320 12400 2372
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 16948 2592 17000 2644
rect 17500 2524 17552 2576
rect 19156 2524 19208 2576
rect 20260 2524 20312 2576
rect 17040 2388 17092 2440
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 16396 2320 16448 2372
rect 17684 2456 17736 2508
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 17868 2388 17920 2440
rect 18696 2456 18748 2508
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 11980 2252 12032 2304
rect 12532 2252 12584 2304
rect 13084 2252 13136 2304
rect 13636 2252 13688 2304
rect 14740 2252 14792 2304
rect 15844 2252 15896 2304
rect 18972 2320 19024 2372
rect 19064 2320 19116 2372
rect 18604 2252 18656 2304
rect 19708 2252 19760 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 8024 2048 8076 2100
rect 16028 2048 16080 2100
rect 7840 1980 7892 2032
rect 14648 1980 14700 2032
rect 19800 2048 19852 2100
rect 9496 1912 9548 1964
rect 17040 1980 17092 2032
rect 20444 1980 20496 2032
rect 14924 1912 14976 1964
rect 22652 1912 22704 1964
rect 1676 1708 1728 1760
rect 13728 1708 13780 1760
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3698 22200 3754 23000
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8312 22222 8616 22250
rect 400 20466 428 22200
rect 388 20460 440 20466
rect 388 20402 440 20408
rect 952 19310 980 22200
rect 1504 19854 1532 22200
rect 2056 19854 2084 22200
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 940 19304 992 19310
rect 940 19246 992 19252
rect 952 18426 980 19246
rect 1504 18426 1532 19790
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 940 18420 992 18426
rect 940 18362 992 18368
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1964 16697 1992 19110
rect 2056 18970 2084 19790
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2042 17776 2098 17785
rect 2042 17711 2044 17720
rect 2096 17711 2098 17720
rect 2044 17682 2096 17688
rect 1950 16688 2006 16697
rect 1950 16623 2006 16632
rect 2148 11257 2176 20334
rect 2240 18426 2268 20402
rect 2332 19310 2360 20742
rect 2608 19854 2636 22200
rect 3160 20482 3188 22200
rect 3056 20460 3108 20466
rect 3160 20454 3280 20482
rect 3712 20466 3740 22200
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3056 20402 3108 20408
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2608 18902 2636 19790
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2792 17105 2820 19722
rect 3068 18426 3096 20402
rect 3252 20398 3280 20454
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3146 19952 3202 19961
rect 3146 19887 3202 19896
rect 3160 19242 3188 19887
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 3160 12753 3188 19178
rect 3252 18358 3280 20334
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3436 20058 3464 20198
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3896 20058 3924 20470
rect 4264 20466 4292 22200
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4158 20088 4214 20097
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3884 20052 3936 20058
rect 4158 20023 4214 20032
rect 3884 19994 3936 20000
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3896 18630 3924 19110
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3146 12744 3202 12753
rect 3146 12679 3202 12688
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 2134 11248 2190 11257
rect 2134 11183 2190 11192
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3896 9994 3924 18566
rect 3988 14414 4016 19926
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4080 14346 4108 19450
rect 4172 19446 4200 20023
rect 4342 19816 4398 19825
rect 4252 19780 4304 19786
rect 4342 19751 4398 19760
rect 4252 19722 4304 19728
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4172 18698 4200 19110
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4172 18426 4200 18634
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4172 17882 4200 18362
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 17218 4200 17478
rect 4264 17338 4292 19722
rect 4356 19718 4384 19751
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4356 19145 4384 19178
rect 4342 19136 4398 19145
rect 4342 19071 4398 19080
rect 4448 18850 4476 20334
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4356 18822 4476 18850
rect 4540 18834 4568 19790
rect 4528 18828 4580 18834
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4172 17190 4292 17218
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16250 4200 16390
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5817 1440 6258
rect 1582 6216 1638 6225
rect 1582 6151 1584 6160
rect 1636 6151 1638 6160
rect 1584 6122 1636 6128
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 4080 5846 4108 13806
rect 4068 5840 4120 5846
rect 1398 5808 1454 5817
rect 4068 5782 4120 5788
rect 1398 5743 1454 5752
rect 4264 5574 4292 17190
rect 4356 14414 4384 18822
rect 4528 18770 4580 18776
rect 4436 18760 4488 18766
rect 4434 18728 4436 18737
rect 4488 18728 4490 18737
rect 4434 18663 4490 18672
rect 4540 18578 4568 18770
rect 4448 18550 4568 18578
rect 4448 14906 4476 18550
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15094 4568 15846
rect 4632 15366 4660 15982
rect 4620 15360 4672 15366
rect 4618 15328 4620 15337
rect 4672 15328 4674 15337
rect 4618 15263 4674 15272
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4448 14878 4568 14906
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 14074 4384 14350
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4540 11626 4568 14878
rect 4724 14414 4752 20266
rect 4816 19378 4844 22200
rect 5368 20466 5396 22200
rect 5722 20496 5778 20505
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5356 20460 5408 20466
rect 5722 20431 5778 20440
rect 5356 20402 5408 20408
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4816 18970 4844 19314
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4908 17202 4936 20198
rect 5000 18358 5028 20402
rect 5092 18902 5120 20402
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 19378 5580 20198
rect 5736 19990 5764 20431
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5920 19854 5948 22200
rect 6472 21298 6500 22200
rect 6472 21270 6592 21298
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6564 20398 6592 21270
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6552 20392 6604 20398
rect 6920 20392 6972 20398
rect 6552 20334 6604 20340
rect 6826 20360 6882 20369
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5540 19372 5592 19378
rect 5460 19332 5540 19360
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4908 16114 4936 16594
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15162 4844 15846
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4908 14906 4936 16050
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 4816 14878 4936 14906
rect 4712 14408 4764 14414
rect 4632 14356 4712 14362
rect 4632 14350 4764 14356
rect 4632 14334 4752 14350
rect 4632 14006 4660 14334
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4632 7834 4660 13942
rect 4724 8906 4752 14214
rect 4816 9450 4844 14878
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4908 11642 4936 14418
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5000 12434 5028 14010
rect 5092 13394 5120 15370
rect 5184 13394 5212 19110
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 18426 5304 18634
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5368 17066 5396 17818
rect 5460 17542 5488 19332
rect 5540 19314 5592 19320
rect 5538 19272 5594 19281
rect 5538 19207 5594 19216
rect 5552 18154 5580 19207
rect 5644 18630 5672 19790
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5736 18154 5764 19314
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16794 5396 17002
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5552 16522 5580 17070
rect 5644 16969 5672 17138
rect 5630 16960 5686 16969
rect 5630 16895 5686 16904
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 15502 5764 16390
rect 5828 16250 5856 19450
rect 5920 18290 5948 19790
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 6012 17814 6040 20334
rect 6920 20334 6972 20340
rect 6826 20295 6882 20304
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6564 18426 6592 19858
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19514 6684 19790
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6656 19417 6684 19450
rect 6642 19408 6698 19417
rect 6642 19343 6698 19352
rect 6748 18902 6776 19722
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5460 14822 5488 15302
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13938 5304 14418
rect 5368 13977 5396 14758
rect 5460 14006 5488 14758
rect 5448 14000 5500 14006
rect 5354 13968 5410 13977
rect 5264 13932 5316 13938
rect 5448 13942 5500 13948
rect 5354 13903 5410 13912
rect 5264 13874 5316 13880
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5000 12406 5120 12434
rect 4908 11614 5028 11642
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4632 7806 4752 7834
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 388 2440 440 2446
rect 388 2382 440 2388
rect 400 800 428 2382
rect 952 800 980 3470
rect 1412 2446 1440 3878
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1504 3058 1532 3402
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1504 800 1532 2994
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 1766 1716 2382
rect 2056 2378 2084 2790
rect 2792 2446 2820 2790
rect 2780 2440 2832 2446
rect 2608 2388 2780 2394
rect 2608 2382 2832 2388
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 2608 2366 2820 2382
rect 3160 2378 3188 2790
rect 3148 2372 3200 2378
rect 1676 1760 1728 1766
rect 1676 1702 1728 1708
rect 2056 800 2084 2314
rect 2608 800 2636 2366
rect 3148 2314 3200 2320
rect 3160 800 3188 2314
rect 386 0 442 800
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3436 762 3464 2926
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 4264 2446 4292 3334
rect 4540 3058 4568 7142
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4632 2514 4660 7686
rect 4724 7313 4752 7806
rect 4710 7304 4766 7313
rect 4710 7239 4766 7248
rect 4908 7206 4936 11494
rect 5000 10062 5028 11614
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 8022 5028 9998
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 5000 7342 5028 7958
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 5092 5710 5120 12406
rect 5276 12220 5304 13874
rect 5460 13852 5488 13942
rect 5368 13824 5488 13852
rect 5368 12628 5396 13824
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5460 12782 5488 13670
rect 5552 12918 5580 15302
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12986 5764 13126
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5722 12744 5778 12753
rect 5722 12679 5724 12688
rect 5776 12679 5778 12688
rect 5724 12650 5776 12656
rect 5368 12600 5580 12628
rect 5552 12322 5580 12600
rect 5828 12434 5856 16050
rect 5736 12406 5856 12434
rect 5552 12294 5672 12322
rect 5276 12192 5488 12220
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5184 7750 5212 9930
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9450 5304 9862
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5368 9217 5396 10066
rect 5460 9518 5488 12192
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5552 11121 5580 11766
rect 5538 11112 5594 11121
rect 5538 11047 5540 11056
rect 5592 11047 5594 11056
rect 5540 11018 5592 11024
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5354 9208 5410 9217
rect 5354 9143 5410 9152
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5276 7546 5304 8366
rect 5368 7954 5396 9143
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5460 7342 5488 9454
rect 5552 8974 5580 10134
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 7886 5580 8366
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5078 4176 5134 4185
rect 5078 4111 5134 4120
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4908 2774 4936 2994
rect 5092 2922 5120 4111
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 3126 5396 3334
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4816 2746 4936 2774
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 3620 870 3740 898
rect 3620 762 3648 870
rect 3712 800 3740 870
rect 4264 800 4292 2382
rect 4816 800 4844 2746
rect 5368 800 5396 3062
rect 5644 2774 5672 12294
rect 5736 10810 5764 12406
rect 5920 12322 5948 17478
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5828 12294 5948 12322
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 9926 5764 10406
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5722 9480 5778 9489
rect 5828 9466 5856 12294
rect 6012 12186 6040 16934
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15473 6408 15846
rect 6552 15496 6604 15502
rect 6366 15464 6422 15473
rect 6552 15438 6604 15444
rect 6366 15399 6422 15408
rect 6380 15366 6408 15399
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6564 15162 6592 15438
rect 6656 15162 6684 18702
rect 6840 18630 6868 20295
rect 6932 19689 6960 20334
rect 7024 20233 7052 22200
rect 7576 20584 7604 22200
rect 7576 20556 7696 20584
rect 7668 20398 7696 20556
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7010 20224 7066 20233
rect 7010 20159 7066 20168
rect 7194 20088 7250 20097
rect 7194 20023 7250 20032
rect 6918 19680 6974 19689
rect 6918 19615 6974 19624
rect 7102 19680 7158 19689
rect 7102 19615 7158 19624
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6918 19348 6974 19357
rect 6918 19283 6974 19292
rect 6932 18902 6960 19283
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6564 13870 6592 13901
rect 6552 13864 6604 13870
rect 6550 13832 6552 13841
rect 6604 13832 6606 13841
rect 6550 13767 6606 13776
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6564 12850 6592 13767
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 5920 12158 6040 12186
rect 5920 9654 5948 12158
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11218 6040 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 10198 6500 10746
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6472 10062 6500 10134
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9722 6040 9862
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 6276 9512 6328 9518
rect 5828 9438 5948 9466
rect 6276 9454 6328 9460
rect 5722 9415 5778 9424
rect 5736 3534 5764 9415
rect 5920 7834 5948 9438
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6012 7954 6040 8978
rect 6288 8838 6316 9454
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5920 7806 6040 7834
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7546 5948 7686
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6012 6769 6040 7806
rect 6564 7732 6592 12310
rect 6748 11898 6776 18226
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16114 6868 16594
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 13682 6868 15370
rect 6932 14618 6960 18702
rect 7024 18426 7052 19450
rect 7116 19446 7144 19615
rect 7208 19514 7236 20023
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7300 19786 7328 19858
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7286 19544 7342 19553
rect 7196 19508 7248 19514
rect 7286 19479 7342 19488
rect 7196 19450 7248 19456
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7194 19408 7250 19417
rect 7194 19343 7250 19352
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 16250 7052 18022
rect 7116 17882 7144 18634
rect 7208 18290 7236 19343
rect 7300 18834 7328 19479
rect 7392 19417 7420 19654
rect 7378 19408 7434 19417
rect 7378 19343 7434 19352
rect 7484 19174 7512 19722
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 16794 7236 17614
rect 7300 17610 7328 18566
rect 7392 18290 7420 18838
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17746 7420 18226
rect 7576 18222 7604 19858
rect 7668 19145 7696 20334
rect 8128 19922 8156 22200
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8312 19802 8340 22222
rect 8588 22114 8616 22222
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11164 22222 11376 22250
rect 8680 22114 8708 22200
rect 8588 22086 8708 22114
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8220 19786 8340 19802
rect 8404 19786 8432 19858
rect 8208 19780 8340 19786
rect 8260 19774 8340 19780
rect 8392 19780 8444 19786
rect 8208 19722 8260 19728
rect 8392 19722 8444 19728
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 8114 19680 8170 19689
rect 7746 19544 7802 19553
rect 7746 19479 7802 19488
rect 7760 19378 7788 19479
rect 7944 19417 7972 19654
rect 8114 19615 8170 19624
rect 8128 19514 8156 19615
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 7930 19408 7986 19417
rect 7748 19372 7800 19378
rect 7930 19343 7986 19352
rect 7748 19314 7800 19320
rect 8404 19310 8432 19722
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 7840 19168 7892 19174
rect 7654 19136 7710 19145
rect 8496 19122 8524 19654
rect 7840 19110 7892 19116
rect 7654 19071 7710 19080
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7300 16046 7328 17546
rect 7668 16130 7696 18566
rect 7852 18426 7880 19110
rect 8404 19094 8524 19122
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 17814 8064 18226
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7748 17672 7800 17678
rect 7746 17640 7748 17649
rect 7800 17640 7802 17649
rect 7746 17575 7802 17584
rect 7760 17338 7788 17575
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7392 16102 7696 16130
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7024 15706 7052 15982
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7116 15162 7144 15574
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6840 13654 6960 13682
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 12306 6868 13466
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6932 12186 6960 13654
rect 6840 12158 6960 12186
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 9178 6684 10542
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6656 7954 6684 8298
rect 6748 8090 6776 10610
rect 6840 10266 6868 12158
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11082 6960 11494
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7024 9042 7052 14214
rect 7208 12434 7236 15914
rect 7392 14958 7420 16102
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7116 12406 7236 12434
rect 7116 9178 7144 12406
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11150 7236 11630
rect 7300 11354 7328 14214
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12434 7420 13126
rect 7392 12406 7512 12434
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7392 11150 7420 12038
rect 7484 11898 7512 12406
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10810 7420 10950
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7208 8974 7236 9318
rect 7300 9178 7328 9454
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7392 8838 7420 9046
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7300 8537 7328 8570
rect 7286 8528 7342 8537
rect 7286 8463 7342 8472
rect 7380 8424 7432 8430
rect 6826 8392 6882 8401
rect 7380 8366 7432 8372
rect 6826 8327 6882 8336
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6564 7704 6776 7732
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 5998 6760 6054 6769
rect 5998 6695 6054 6704
rect 6104 6644 6132 7414
rect 6012 6616 6132 6644
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5722 3224 5778 3233
rect 5722 3159 5778 3168
rect 5736 3126 5764 3159
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5644 2746 5764 2774
rect 5630 2680 5686 2689
rect 5736 2650 5764 2746
rect 5630 2615 5686 2624
rect 5724 2644 5776 2650
rect 5644 2514 5672 2615
rect 5724 2586 5776 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5644 2417 5672 2450
rect 5630 2408 5686 2417
rect 5920 2378 5948 3334
rect 6012 2446 6040 6616
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6748 5098 6776 7704
rect 6840 7478 6868 8327
rect 7392 8294 7420 8366
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7546 7144 7686
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 7002 6868 7414
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6564 2378 6592 2790
rect 5630 2343 5686 2352
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 5920 800 5948 2314
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 1850 6592 2314
rect 6748 2310 6776 5034
rect 6840 3738 6868 6734
rect 7484 6225 7512 11630
rect 7576 11354 7604 14962
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 11150 7696 13194
rect 7852 12442 7880 17750
rect 8220 17678 8248 18906
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8220 16658 8248 17274
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15094 7972 15846
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7576 9926 7604 11086
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7576 6066 7604 9862
rect 7668 6254 7696 11086
rect 7760 10690 7788 11834
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11354 7880 11698
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7944 10742 7972 12378
rect 8036 11898 8064 16390
rect 8128 15434 8156 16390
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8220 12434 8248 15574
rect 8312 12442 8340 15846
rect 8128 12406 8248 12434
rect 8300 12436 8352 12442
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11286 8064 11698
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8022 11112 8078 11121
rect 8022 11047 8078 11056
rect 8036 11014 8064 11047
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7932 10736 7984 10742
rect 7760 10662 7880 10690
rect 7932 10678 7984 10684
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 9994 7788 10542
rect 7852 10062 7880 10662
rect 8036 10470 8064 10950
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8090 7788 9522
rect 7852 9042 7880 9998
rect 7930 9208 7986 9217
rect 8036 9194 8064 10406
rect 8128 9654 8156 12406
rect 8300 12378 8352 12384
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8220 11218 8248 12310
rect 8404 11880 8432 19094
rect 8588 18766 8616 19110
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 17542 8616 18702
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17270 8616 17478
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8588 17066 8616 17206
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16658 8616 17002
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8588 16182 8616 16594
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8588 15706 8616 16118
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8574 14920 8630 14929
rect 8574 14855 8576 14864
rect 8628 14855 8630 14864
rect 8576 14826 8628 14832
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12374 8524 12582
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8312 11852 8432 11880
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8312 10130 8340 11852
rect 8588 11778 8616 14554
rect 8404 11750 8616 11778
rect 8404 11694 8432 11750
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 10810 8616 11630
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8390 10160 8446 10169
rect 8300 10124 8352 10130
rect 8390 10095 8446 10104
rect 8300 10066 8352 10072
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8312 9518 8340 10066
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8404 9450 8432 10095
rect 8680 9654 8708 20198
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 9232 19553 9260 22200
rect 9312 20392 9364 20398
rect 9784 20346 9812 22200
rect 10336 20534 10364 22200
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9312 20334 9364 20340
rect 9218 19544 9274 19553
rect 9324 19514 9352 20334
rect 9600 20318 9812 20346
rect 9494 20088 9550 20097
rect 9494 20023 9550 20032
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9218 19479 9274 19488
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9126 19136 9182 19145
rect 8747 19068 9055 19077
rect 9126 19071 9182 19080
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8956 18698 8984 18838
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8956 18222 8984 18634
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15910 8984 16458
rect 9140 16250 9168 19071
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9232 18358 9260 18906
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9232 16946 9260 18294
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9324 17542 9352 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 9324 17134 9352 17167
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9232 16918 9352 16946
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 15162 9076 15642
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 15337 9260 15370
rect 9218 15328 9274 15337
rect 9218 15263 9274 15272
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 13841 9260 14010
rect 9218 13832 9274 13841
rect 9324 13802 9352 16918
rect 9218 13767 9274 13776
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9036 13320 9088 13326
rect 9140 13308 9168 13670
rect 9088 13280 9168 13308
rect 9036 13262 9088 13268
rect 9048 12918 9076 13262
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9036 12912 9088 12918
rect 9088 12872 9168 12900
rect 9324 12889 9352 13194
rect 9036 12854 9088 12860
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9140 12238 9168 12872
rect 9310 12880 9366 12889
rect 9220 12844 9272 12850
rect 9310 12815 9366 12824
rect 9220 12786 9272 12792
rect 9232 12434 9260 12786
rect 9232 12406 9352 12434
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9324 11558 9352 12406
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 10606 9076 11086
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8036 9166 8156 9194
rect 7930 9143 7986 9152
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7018 7880 8978
rect 7944 8634 7972 9143
rect 8022 9072 8078 9081
rect 8022 9007 8078 9016
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 8022 7972 8366
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 8036 7546 8064 9007
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7852 6990 7972 7018
rect 7838 6896 7894 6905
rect 7838 6831 7840 6840
rect 7892 6831 7894 6840
rect 7840 6802 7892 6808
rect 7944 6458 7972 6990
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7576 6038 7696 6066
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7300 3194 7328 5607
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2446 7052 2790
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6472 1822 6592 1850
rect 6472 800 6500 1822
rect 7024 800 7052 2382
rect 7576 2378 7604 2858
rect 7668 2650 7696 6038
rect 7944 4690 7972 6394
rect 8022 5808 8078 5817
rect 8128 5794 8156 9166
rect 8300 8560 8352 8566
rect 8206 8528 8262 8537
rect 8300 8502 8352 8508
rect 8206 8463 8208 8472
rect 8260 8463 8262 8472
rect 8208 8434 8260 8440
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 8022 8248 8230
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8206 7848 8262 7857
rect 8206 7783 8262 7792
rect 8220 6866 8248 7783
rect 8312 7274 8340 8502
rect 9140 8430 9168 10950
rect 9324 10130 9352 11494
rect 9416 11014 9444 19722
rect 9508 19718 9536 20023
rect 9600 19922 9628 20318
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9508 18850 9536 19450
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9600 18970 9628 19314
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9508 18822 9628 18850
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17542 9536 17750
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9600 15314 9628 18822
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9784 15638 9812 18226
rect 9876 17202 9904 19654
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9968 16561 9996 20402
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10336 19786 10364 20334
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10704 20058 10732 20198
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10324 19780 10376 19786
rect 10324 19722 10376 19728
rect 10336 19446 10364 19722
rect 10888 19718 10916 22200
rect 11164 20466 11192 22222
rect 11348 22114 11376 22222
rect 11426 22200 11482 23000
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13634 22200 13690 23000
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 15290 22200 15346 23000
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21560 22222 21864 22250
rect 11440 22114 11468 22200
rect 11348 22086 11468 22114
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 18290 10732 18702
rect 10796 18426 10824 19178
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10980 18086 11008 19246
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 17082 10180 17138
rect 10060 17054 10180 17082
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9600 15286 9720 15314
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9508 12889 9536 14894
rect 9600 14550 9628 15098
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9692 14396 9720 15286
rect 9968 15026 9996 15846
rect 10060 15706 10088 17054
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16182 10272 16934
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 14906 9996 14962
rect 9600 14368 9720 14396
rect 9784 14878 9996 14906
rect 9494 12880 9550 12889
rect 9494 12815 9550 12824
rect 9600 12730 9628 14368
rect 9508 12702 9628 12730
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9402 10840 9458 10849
rect 9402 10775 9404 10784
rect 9456 10775 9458 10784
rect 9404 10746 9456 10752
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9310 10024 9366 10033
rect 9310 9959 9366 9968
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 9140 7954 9168 8230
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9232 7546 9260 9522
rect 9324 9178 9352 9959
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9324 8022 9352 9114
rect 9508 8786 9536 12702
rect 9784 12458 9812 14878
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13190 9904 13670
rect 9968 13190 9996 14282
rect 10060 13938 10088 15642
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9600 12430 9812 12458
rect 9876 12434 9904 13126
rect 9968 12646 9996 13126
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9600 9042 9628 12430
rect 9876 12406 9996 12434
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9692 11558 9720 12271
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11762 9904 12106
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 10554 9720 10610
rect 9692 10526 9812 10554
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9692 9926 9720 10134
rect 9784 9994 9812 10526
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9692 8974 9720 9318
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9416 8758 9536 8786
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 8574 7440 8630 7449
rect 8574 7375 8630 7384
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8482 6896 8538 6905
rect 8208 6860 8260 6866
rect 8482 6831 8538 6840
rect 8208 6802 8260 6808
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8078 5766 8156 5794
rect 8220 5778 8248 6190
rect 8208 5772 8260 5778
rect 8022 5743 8078 5752
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 8036 4162 8064 5743
rect 8208 5714 8260 5720
rect 8392 5568 8444 5574
rect 8206 5536 8262 5545
rect 8392 5510 8444 5516
rect 8206 5471 8262 5480
rect 7944 4134 8064 4162
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7576 800 7604 2314
rect 7852 2038 7880 3878
rect 7944 2650 7972 4134
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8036 2106 8064 3878
rect 8220 3670 8248 5471
rect 8404 5370 8432 5510
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8404 5137 8432 5306
rect 8390 5128 8446 5137
rect 8390 5063 8446 5072
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8312 3097 8340 3402
rect 8404 3398 8432 5063
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8496 3126 8524 6831
rect 8588 5914 8616 7375
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9128 6792 9180 6798
rect 8666 6760 8722 6769
rect 8666 6695 8722 6704
rect 9126 6760 9128 6769
rect 9180 6760 9182 6769
rect 9126 6695 9182 6704
rect 8680 6497 8708 6695
rect 8666 6488 8722 6497
rect 8666 6423 8722 6432
rect 8680 5914 8708 6423
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 4146 8616 5578
rect 8680 5370 8708 5850
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9140 4826 9168 6258
rect 9218 4856 9274 4865
rect 9128 4820 9180 4826
rect 9218 4791 9274 4800
rect 9128 4762 9180 4768
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8852 4072 8904 4078
rect 8850 4040 8852 4049
rect 8904 4040 8906 4049
rect 8850 3975 8906 3984
rect 9232 3942 9260 4791
rect 9416 4622 9444 8758
rect 9600 8634 9628 8774
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9508 8514 9536 8570
rect 9508 8486 9720 8514
rect 9692 8430 9720 8486
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 6798 9536 8230
rect 9600 7478 9628 8366
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9784 7206 9812 9930
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9722 9904 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 7342 9904 8978
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9876 6882 9904 7278
rect 9692 6854 9904 6882
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9692 5794 9720 6854
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9600 5766 9720 5794
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9404 4616 9456 4622
rect 9310 4584 9366 4593
rect 9404 4558 9456 4564
rect 9508 4570 9536 5646
rect 9600 5250 9628 5766
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 5370 9720 5646
rect 9784 5574 9812 6598
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9600 5222 9720 5250
rect 9692 4690 9720 5222
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9310 4519 9312 4528
rect 9364 4519 9366 4528
rect 9312 4490 9364 4496
rect 9416 4214 9444 4558
rect 9508 4542 9628 4570
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 8576 3936 8628 3942
rect 8574 3904 8576 3913
rect 9220 3936 9272 3942
rect 8628 3904 8630 3913
rect 9220 3878 9272 3884
rect 8574 3839 8630 3848
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8484 3120 8536 3126
rect 8298 3088 8354 3097
rect 8116 3052 8168 3058
rect 8484 3062 8536 3068
rect 8298 3023 8354 3032
rect 9220 3052 9272 3058
rect 8116 2994 8168 3000
rect 9220 2994 9272 3000
rect 8128 2360 8156 2994
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2446 8524 2790
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8300 2372 8352 2378
rect 8128 2332 8300 2360
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 8128 800 8156 2332
rect 8300 2314 8352 2320
rect 8680 800 8708 2382
rect 9232 800 9260 2994
rect 9310 2544 9366 2553
rect 9310 2479 9312 2488
rect 9364 2479 9366 2488
rect 9312 2450 9364 2456
rect 9508 1970 9536 4422
rect 9600 3074 9628 4542
rect 9772 4072 9824 4078
rect 9876 4049 9904 6734
rect 9968 6254 9996 12406
rect 10060 12102 10088 12582
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 10606 10088 12038
rect 10152 11393 10180 12922
rect 10138 11384 10194 11393
rect 10138 11319 10194 11328
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10060 9738 10088 10202
rect 10152 10198 10180 10746
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10060 9710 10180 9738
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10060 9518 10088 9551
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10152 9042 10180 9710
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10140 8900 10192 8906
rect 10244 8888 10272 16118
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10336 14618 10364 14962
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10336 12442 10364 13874
rect 10428 13734 10456 15302
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10324 12436 10376 12442
rect 10520 12434 10548 12922
rect 10324 12378 10376 12384
rect 10428 12406 10548 12434
rect 10612 12434 10640 18022
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 16114 10732 16526
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10704 15910 10732 16050
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10796 13530 10824 17546
rect 10888 17542 10916 17750
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 15094 11008 17478
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10980 13938 11008 14010
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10612 12406 10732 12434
rect 10428 12322 10456 12406
rect 10336 12294 10456 12322
rect 10508 12300 10560 12306
rect 10336 11762 10364 12294
rect 10508 12242 10560 12248
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10192 8860 10272 8888
rect 10140 8842 10192 8848
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 8514 10088 8774
rect 10060 8486 10180 8514
rect 10244 8498 10272 8860
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10060 8090 10088 8298
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7410 10088 8026
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10152 6474 10180 8486
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 8090 10364 10678
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10428 9722 10456 10610
rect 10520 10606 10548 12242
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10520 9178 10548 10066
rect 10612 9761 10640 12174
rect 10704 10810 10732 12406
rect 10796 12170 10824 13466
rect 11072 12209 11100 20334
rect 11164 19938 11192 20402
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11164 19910 11284 19938
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11164 18154 11192 19722
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11150 17776 11206 17785
rect 11150 17711 11206 17720
rect 11164 13297 11192 17711
rect 11256 17241 11284 19910
rect 11532 19718 11560 20334
rect 11624 20058 11652 20334
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11348 19145 11376 19450
rect 11518 19408 11574 19417
rect 11518 19343 11520 19352
rect 11572 19343 11574 19352
rect 11520 19314 11572 19320
rect 11334 19136 11390 19145
rect 11334 19071 11390 19080
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11242 17232 11298 17241
rect 11242 17167 11298 17176
rect 11716 16674 11744 20470
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11900 19922 11928 20266
rect 11992 20058 12020 22200
rect 12544 20602 12572 22200
rect 13096 20602 13124 22200
rect 13648 20618 13676 22200
rect 13648 20602 13860 20618
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 13084 20596 13136 20602
rect 13648 20596 13872 20602
rect 13648 20590 13820 20596
rect 13084 20538 13136 20544
rect 13820 20538 13872 20544
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12084 19666 12112 20334
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 11808 19638 12112 19666
rect 11808 17814 11836 19638
rect 12176 19514 12204 19926
rect 12544 19854 12572 20266
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11900 17678 11928 19450
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 18290 12296 18566
rect 12452 18426 12480 19314
rect 12530 19136 12586 19145
rect 12530 19071 12586 19080
rect 12544 18766 12572 19071
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12636 18426 12664 19654
rect 12992 19440 13044 19446
rect 12898 19408 12954 19417
rect 12992 19382 13044 19388
rect 12898 19343 12954 19352
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12162 17912 12218 17921
rect 12162 17847 12164 17856
rect 12216 17847 12218 17856
rect 12164 17818 12216 17824
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17338 12204 17546
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11716 16646 11836 16674
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15570 11744 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15434 11744 15506
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 15162 11744 15370
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11716 14006 11744 14758
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11150 13288 11206 13297
rect 11150 13223 11206 13232
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12306 11192 12582
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11058 12200 11114 12209
rect 10784 12164 10836 12170
rect 11058 12135 11114 12144
rect 10784 12106 10836 12112
rect 10796 11880 10824 12106
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10796 11852 11008 11880
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10598 9752 10654 9761
rect 10598 9687 10654 9696
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10612 9110 10640 9318
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8634 10456 8774
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 7970 10456 8570
rect 10336 7942 10456 7970
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10060 6446 10180 6474
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10060 5302 10088 6446
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5914 10180 6258
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10244 5545 10272 7346
rect 10230 5536 10286 5545
rect 10230 5471 10286 5480
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 4014 9824 4020
rect 9862 4040 9918 4049
rect 9784 3505 9812 4014
rect 9862 3975 9918 3984
rect 9876 3670 9904 3975
rect 9968 3670 9996 4626
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9770 3496 9826 3505
rect 9770 3431 9826 3440
rect 9956 3460 10008 3466
rect 9600 3046 9720 3074
rect 9784 3058 9812 3431
rect 9956 3402 10008 3408
rect 9692 2990 9720 3046
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9968 2446 9996 3402
rect 10060 3058 10088 5238
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10152 4690 10180 5102
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10336 2774 10364 7942
rect 10416 7200 10468 7206
rect 10414 7168 10416 7177
rect 10468 7168 10470 7177
rect 10414 7103 10470 7112
rect 10244 2746 10364 2774
rect 10244 2650 10272 2746
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10428 2582 10456 7103
rect 10520 7041 10548 8978
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10612 7546 10640 8366
rect 10704 7546 10732 10542
rect 10796 9042 10824 11698
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11150 10916 11494
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10742 10916 11086
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10980 10606 11008 11852
rect 11072 11762 11100 12038
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11072 11626 11100 11698
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11058 11520 11114 11529
rect 11058 11455 11114 11464
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11072 9674 11100 11455
rect 10888 9646 11100 9674
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10888 7936 10916 9646
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 11072 8430 11100 8599
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 7970 11100 8366
rect 10796 7908 10916 7936
rect 10980 7942 11100 7970
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10796 7410 10824 7908
rect 10980 7868 11008 7942
rect 10888 7840 11008 7868
rect 11060 7880 11112 7886
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10690 7304 10746 7313
rect 10690 7239 10746 7248
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10520 6934 10548 6967
rect 10704 6934 10732 7239
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5817 10548 6054
rect 10506 5808 10562 5817
rect 10506 5743 10562 5752
rect 10612 4826 10640 6326
rect 10704 6118 10732 6870
rect 10796 6662 10824 6938
rect 10888 6730 10916 7840
rect 11060 7822 11112 7828
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 6866 11008 7686
rect 11072 7313 11100 7822
rect 11058 7304 11114 7313
rect 11058 7239 11114 7248
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5370 10732 5850
rect 10888 5642 10916 6666
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10796 4214 10824 4762
rect 10968 4616 11020 4622
rect 11072 4604 11100 6870
rect 11164 5778 11192 12038
rect 11256 10810 11284 13806
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11624 12170 11652 12854
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11257 11468 11698
rect 11426 11248 11482 11257
rect 11532 11218 11560 11834
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11354 11652 11494
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11426 11183 11482 11192
rect 11520 11212 11572 11218
rect 11440 11082 11468 11183
rect 11520 11154 11572 11160
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11520 11008 11572 11014
rect 11716 10996 11744 13466
rect 11572 10968 11744 10996
rect 11520 10950 11572 10956
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11716 9654 11744 10968
rect 11808 10305 11836 16646
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15502 12020 15846
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11794 10296 11850 10305
rect 11794 10231 11850 10240
rect 11900 10180 11928 14894
rect 11992 14618 12020 15098
rect 12084 14890 12112 16390
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 12176 14890 12204 15030
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 14074 12020 14554
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11992 13938 12020 14010
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11992 13326 12020 13874
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12162 13288 12218 13297
rect 12162 13223 12218 13232
rect 12176 13190 12204 13223
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11992 12782 12020 13126
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12102 12020 12718
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 11286 12020 11698
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11808 10152 11928 10180
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11256 5914 11284 9590
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11716 8906 11744 9415
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11716 8634 11744 8842
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11348 7954 11376 8230
rect 11440 8022 11468 8230
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11716 7478 11744 7686
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11532 7002 11560 7278
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11702 6216 11758 6225
rect 11702 6151 11758 6160
rect 11716 5914 11744 6151
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11020 4576 11100 4604
rect 10968 4558 11020 4564
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 4298 10916 4490
rect 10966 4312 11022 4321
rect 10888 4270 10966 4298
rect 11072 4282 11100 4576
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4282 11192 4422
rect 10966 4247 11022 4256
rect 11060 4276 11112 4282
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10980 4078 11008 4247
rect 11060 4218 11112 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11150 4176 11206 4185
rect 11150 4111 11206 4120
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3670 11008 4014
rect 10508 3664 10560 3670
rect 10506 3632 10508 3641
rect 10968 3664 11020 3670
rect 10560 3632 10562 3641
rect 10968 3606 11020 3612
rect 10506 3567 10562 3576
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10520 2446 10548 2858
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 9956 2440 10008 2446
rect 9784 2400 9956 2428
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9784 800 9812 2400
rect 10508 2440 10560 2446
rect 9956 2382 10008 2388
rect 10336 2400 10508 2428
rect 10336 800 10364 2400
rect 10508 2382 10560 2388
rect 10888 800 10916 2450
rect 10980 2446 11008 3470
rect 11164 3194 11192 4111
rect 11256 3534 11284 5510
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11716 5370 11744 5578
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11808 4690 11836 10152
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11900 8838 11928 9862
rect 11992 9178 12020 10678
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8401 12020 8774
rect 11978 8392 12034 8401
rect 11978 8327 12034 8336
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7546 11928 8230
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11150 2952 11206 2961
rect 11256 2922 11284 3334
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11716 3058 11744 4422
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11150 2887 11152 2896
rect 11204 2887 11206 2896
rect 11244 2916 11296 2922
rect 11152 2858 11204 2864
rect 11244 2858 11296 2864
rect 10968 2440 11020 2446
rect 11020 2400 11100 2428
rect 10968 2382 11020 2388
rect 3436 734 3648 762
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11072 762 11100 2400
rect 11520 2372 11572 2378
rect 11900 2360 11928 7346
rect 11992 7206 12020 7822
rect 12084 7342 12112 12786
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11898 12204 12106
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11286 12204 11630
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10441 12204 10950
rect 12268 10656 12296 18226
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12452 17542 12480 17818
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12348 16652 12400 16658
rect 12452 16640 12480 16934
rect 12400 16612 12480 16640
rect 12348 16594 12400 16600
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12360 10810 12388 14282
rect 12452 11558 12480 16612
rect 12544 14278 12572 17478
rect 12636 15910 12664 18362
rect 12716 18352 12768 18358
rect 12714 18320 12716 18329
rect 12768 18320 12770 18329
rect 12714 18255 12770 18264
rect 12820 17921 12848 18838
rect 12806 17912 12862 17921
rect 12806 17847 12862 17856
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12728 14890 12756 16050
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12544 12102 12572 13942
rect 12636 13705 12664 14214
rect 12820 13954 12848 16390
rect 12912 14278 12940 19343
rect 13004 19174 13032 19382
rect 13280 19242 13308 20402
rect 13544 20392 13596 20398
rect 13542 20360 13544 20369
rect 13596 20360 13598 20369
rect 14200 20330 14228 22200
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 13542 20295 13598 20304
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13726 20088 13782 20097
rect 13945 20091 14253 20100
rect 13726 20023 13782 20032
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13464 18970 13492 19790
rect 13740 19446 13768 20023
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 13004 18601 13032 18634
rect 12990 18592 13046 18601
rect 12990 18527 13046 18536
rect 13096 16590 13124 18770
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13556 18426 13584 18702
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13372 18290 13400 18362
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16697 13308 17138
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13266 16688 13322 16697
rect 13266 16623 13322 16632
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13266 15464 13322 15473
rect 13266 15399 13322 15408
rect 13280 15366 13308 15399
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 14550 13308 15302
rect 13372 15026 13400 16458
rect 13464 16114 13492 16594
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15570 13492 16050
rect 13556 15706 13584 16730
rect 13648 16182 13676 18702
rect 13740 18630 13768 19110
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13832 17882 13860 19314
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 18601 14228 18702
rect 14186 18592 14242 18601
rect 14186 18527 14242 18536
rect 14200 18290 14228 18527
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14292 18272 14320 19654
rect 14384 19530 14412 19858
rect 14476 19718 14504 19926
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14384 19502 14504 19530
rect 14568 19514 14596 20810
rect 14752 20602 14780 22200
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 19666 15148 19722
rect 14752 19638 15148 19666
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18766 14412 19246
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14372 18284 14424 18290
rect 14292 18244 14372 18272
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13832 15366 13860 16050
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13820 15360 13872 15366
rect 14188 15360 14240 15366
rect 13820 15302 13872 15308
rect 14186 15328 14188 15337
rect 14240 15328 14242 15337
rect 14186 15263 14242 15272
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 13556 14006 13584 14962
rect 13740 14618 13768 15030
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 12992 14000 13044 14006
rect 12728 13926 12848 13954
rect 12912 13948 12992 13954
rect 12912 13942 13044 13948
rect 13544 14000 13596 14006
rect 13648 13977 13676 14010
rect 13544 13942 13596 13948
rect 13634 13968 13690 13977
rect 12912 13926 13032 13942
rect 12622 13696 12678 13705
rect 12622 13631 12678 13640
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10810 12480 10950
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12348 10668 12400 10674
rect 12268 10628 12348 10656
rect 12348 10610 12400 10616
rect 12162 10432 12218 10441
rect 12162 10367 12218 10376
rect 12162 10296 12218 10305
rect 12162 10231 12218 10240
rect 12176 9897 12204 10231
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 12162 9480 12218 9489
rect 12162 9415 12164 9424
rect 12216 9415 12218 9424
rect 12164 9386 12216 9392
rect 12268 9024 12296 9551
rect 12176 8996 12296 9024
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11992 6497 12020 6666
rect 11978 6488 12034 6497
rect 11978 6423 11980 6432
rect 12032 6423 12034 6432
rect 11980 6394 12032 6400
rect 11992 6363 12020 6394
rect 12176 6322 12204 8996
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 12268 8634 12296 8871
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12360 8378 12388 10610
rect 12360 8362 12480 8378
rect 12360 8356 12492 8362
rect 12360 8350 12440 8356
rect 12440 8298 12492 8304
rect 12544 7970 12572 12038
rect 12636 11286 12664 13194
rect 12728 11801 12756 13926
rect 12912 13818 12940 13926
rect 13634 13903 13690 13912
rect 12820 13790 12940 13818
rect 12714 11792 12770 11801
rect 12714 11727 12770 11736
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12714 11248 12770 11257
rect 12714 11183 12770 11192
rect 12624 11144 12676 11150
rect 12622 11112 12624 11121
rect 12676 11112 12678 11121
rect 12622 11047 12678 11056
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 8090 12664 9862
rect 12728 9489 12756 11183
rect 12714 9480 12770 9489
rect 12714 9415 12770 9424
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12544 7954 12664 7970
rect 12544 7948 12676 7954
rect 12544 7942 12624 7948
rect 12624 7890 12676 7896
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12360 7274 12388 7482
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11992 4729 12020 5850
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11978 4720 12034 4729
rect 11978 4655 12034 4664
rect 11992 4078 12020 4655
rect 12176 4282 12204 5102
rect 12268 5098 12296 7142
rect 12360 6934 12388 7210
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12360 3466 12388 6122
rect 12452 5681 12480 7822
rect 12728 7750 12756 8842
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12622 7576 12678 7585
rect 12622 7511 12678 7520
rect 12530 7032 12586 7041
rect 12530 6967 12586 6976
rect 12544 6934 12572 6967
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12636 6730 12664 7511
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5710 12572 6598
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12532 5704 12584 5710
rect 12438 5672 12494 5681
rect 12636 5681 12664 6122
rect 12532 5646 12584 5652
rect 12622 5672 12678 5681
rect 12438 5607 12494 5616
rect 12622 5607 12678 5616
rect 12728 5114 12756 7346
rect 12820 6338 12848 13790
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 12898 12880 12954 12889
rect 12898 12815 12954 12824
rect 12912 11898 12940 12815
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12990 11792 13046 11801
rect 12990 11727 13046 11736
rect 12898 10976 12954 10985
rect 12898 10911 12954 10920
rect 12912 9518 12940 10911
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13004 8498 13032 11727
rect 13082 10840 13138 10849
rect 13082 10775 13138 10784
rect 13096 10742 13124 10775
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13082 7984 13138 7993
rect 13082 7919 13138 7928
rect 13096 7313 13124 7919
rect 13188 7324 13216 12106
rect 13280 9738 13308 12310
rect 13358 11928 13414 11937
rect 13358 11863 13414 11872
rect 13372 10266 13400 11863
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11354 13492 11494
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13464 10062 13492 10950
rect 13556 10606 13584 12310
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13556 9926 13584 10406
rect 13648 10130 13676 13670
rect 13740 13394 13768 14554
rect 13832 13938 13860 14826
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12918 13768 13330
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13740 12442 13768 12854
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 14186 12336 14242 12345
rect 14186 12271 14242 12280
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 10810 13768 11630
rect 14200 11626 14228 12271
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13634 9752 13690 9761
rect 13280 9710 13400 9738
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 9042 13308 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13268 7336 13320 7342
rect 13082 7304 13138 7313
rect 13188 7296 13268 7324
rect 13268 7278 13320 7284
rect 13082 7239 13138 7248
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 6934 13032 7142
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13266 6896 13322 6905
rect 12912 6730 12940 6870
rect 13266 6831 13322 6840
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6440 13032 6598
rect 13004 6412 13216 6440
rect 12820 6310 13032 6338
rect 13188 6322 13216 6412
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5846 12848 6122
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5846 12940 6054
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 13004 5250 13032 6310
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13082 5536 13138 5545
rect 13082 5471 13138 5480
rect 12912 5222 13032 5250
rect 12728 5086 12848 5114
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12728 4282 12756 4558
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 4010 12664 4082
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3534 12572 3878
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12084 2446 12112 3334
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12360 2378 12388 2790
rect 12636 2446 12664 3334
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2446 12756 2790
rect 12820 2514 12848 5086
rect 12912 4690 12940 5222
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 13004 4622 13032 5102
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13096 4146 13124 5471
rect 13280 5166 13308 6831
rect 13372 6254 13400 9710
rect 13634 9687 13690 9696
rect 13648 9654 13676 9687
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13450 8936 13506 8945
rect 13450 8871 13506 8880
rect 13464 7546 13492 8871
rect 13648 7834 13676 9590
rect 13740 8634 13768 9998
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 8294 13768 8434
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13740 7857 13768 7958
rect 13556 7806 13676 7834
rect 13726 7848 13782 7857
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6390 13492 6598
rect 13556 6458 13584 7806
rect 13726 7783 13782 7792
rect 13636 7744 13688 7750
rect 13634 7712 13636 7721
rect 13688 7712 13690 7721
rect 13634 7647 13690 7656
rect 13832 7546 13860 10542
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13910 10024 13966 10033
rect 13910 9959 13966 9968
rect 13924 9722 13952 9959
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14016 9450 14044 10202
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9654 14136 9862
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14292 8430 14320 18244
rect 14372 18226 14424 18232
rect 14476 17678 14504 19502
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14648 19508 14700 19514
rect 14752 19496 14780 19638
rect 14700 19468 14780 19496
rect 14832 19508 14884 19514
rect 14648 19450 14700 19456
rect 14832 19450 14884 19456
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14660 16017 14688 19450
rect 14844 17882 14872 19450
rect 15212 18970 15240 20402
rect 15304 20330 15332 22200
rect 15856 20602 15884 22200
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 15108 18760 15160 18766
rect 14922 18728 14978 18737
rect 14922 18663 14978 18672
rect 15106 18728 15108 18737
rect 15160 18728 15162 18737
rect 15106 18663 15162 18672
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14740 17672 14792 17678
rect 14738 17640 14740 17649
rect 14792 17640 14794 17649
rect 14738 17575 14794 17584
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14646 16008 14702 16017
rect 14646 15943 14702 15952
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14384 11898 14412 15642
rect 14752 15366 14780 17206
rect 14936 15586 14964 18663
rect 15396 17898 15424 20402
rect 15764 19825 15792 20402
rect 16408 20330 16436 22200
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16670 20496 16726 20505
rect 16670 20431 16672 20440
rect 16724 20431 16726 20440
rect 16672 20402 16724 20408
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16028 19848 16080 19854
rect 15750 19816 15806 19825
rect 16028 19790 16080 19796
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 15750 19751 15806 19760
rect 16040 19378 16068 19790
rect 16316 19514 16344 19790
rect 16776 19718 16804 20334
rect 16960 20262 16988 22200
rect 17512 20602 17540 22200
rect 17958 20904 18014 20913
rect 17958 20839 17960 20848
rect 18012 20839 18014 20848
rect 17960 20810 18012 20816
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15580 18154 15608 18362
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15304 17870 15424 17898
rect 15304 17762 15332 17870
rect 15028 17746 15332 17762
rect 15016 17740 15332 17746
rect 15068 17734 15332 17740
rect 15016 17682 15068 17688
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17202 15148 17614
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15212 16590 15240 17546
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16726 15332 17070
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14936 15558 15056 15586
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14936 15162 14964 15370
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14752 14958 14780 15098
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14464 14816 14516 14822
rect 14462 14784 14464 14793
rect 14516 14784 14518 14793
rect 15028 14770 15056 15558
rect 14462 14719 14518 14728
rect 14936 14742 15056 14770
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14844 14346 14872 14554
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13258 14780 13670
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12782 14504 13126
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 12434 14504 12718
rect 14752 12442 14780 12854
rect 14740 12436 14792 12442
rect 14476 12406 14596 12434
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 10810 14412 11698
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10130 14412 10542
rect 14476 10266 14504 11086
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14384 9178 14412 9454
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14476 8566 14504 9590
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14292 7954 14320 8366
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13648 6610 13676 7482
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13740 6798 13768 7239
rect 13818 7168 13874 7177
rect 13818 7103 13874 7112
rect 13832 7002 13860 7103
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 14096 6656 14148 6662
rect 13648 6582 13768 6610
rect 14096 6598 14148 6604
rect 13544 6452 13596 6458
rect 13596 6412 13676 6440
rect 13544 6394 13596 6400
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13360 6248 13412 6254
rect 13544 6248 13596 6254
rect 13360 6190 13412 6196
rect 13464 6208 13544 6236
rect 13372 5234 13400 6190
rect 13464 5642 13492 6208
rect 13544 6190 13596 6196
rect 13542 5808 13598 5817
rect 13542 5743 13544 5752
rect 13596 5743 13598 5752
rect 13544 5714 13596 5720
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13556 4826 13584 5170
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13464 4622 13492 4762
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13556 4078 13584 4626
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 2514 12940 3334
rect 13004 3058 13032 3606
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 3126 13400 3334
rect 13464 3194 13492 4014
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 13372 2446 13400 2790
rect 13648 2582 13676 6412
rect 13740 5846 13768 6582
rect 14108 6254 14136 6598
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5137 13768 5646
rect 13832 5370 13860 6054
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5681 14320 7754
rect 14384 7478 14412 8230
rect 14476 7750 14504 8366
rect 14568 8090 14596 12406
rect 14740 12378 14792 12384
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14660 9722 14688 11834
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14646 9616 14702 9625
rect 14646 9551 14648 9560
rect 14700 9551 14702 9560
rect 14648 9522 14700 9528
rect 14660 8838 14688 9522
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14568 7546 14596 7754
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14372 7472 14424 7478
rect 14660 7426 14688 8774
rect 14372 7414 14424 7420
rect 14476 7398 14688 7426
rect 14370 7168 14426 7177
rect 14370 7103 14426 7112
rect 14384 7002 14412 7103
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14278 5672 14334 5681
rect 14278 5607 14334 5616
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13726 5128 13782 5137
rect 13726 5063 13782 5072
rect 13820 5092 13872 5098
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 11572 2332 11928 2360
rect 12348 2372 12400 2378
rect 11520 2314 11572 2320
rect 12348 2314 12400 2320
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11348 870 11468 898
rect 11348 762 11376 870
rect 11440 800 11468 870
rect 11992 800 12020 2246
rect 12544 800 12572 2246
rect 13096 800 13124 2246
rect 13648 800 13676 2246
rect 13740 1766 13768 5063
rect 13820 5034 13872 5040
rect 13832 4729 13860 5034
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14292 4826 14320 4966
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 13818 4720 13874 4729
rect 13818 4655 13874 4664
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13832 4146 13860 4422
rect 14200 4282 14228 4422
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 4049 13860 4082
rect 13818 4040 13874 4049
rect 13818 3975 13874 3984
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14186 3496 14242 3505
rect 14292 3482 14320 3975
rect 14242 3454 14320 3482
rect 14186 3431 14242 3440
rect 14200 3194 14228 3431
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14384 2990 14412 4218
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14476 2774 14504 7398
rect 14752 7324 14780 12038
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 9586 14872 10950
rect 14936 10266 14964 14742
rect 15304 14362 15332 16662
rect 15028 14334 15332 14362
rect 15028 11558 15056 14334
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15120 12102 15148 14214
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15384 12844 15436 12850
rect 15488 12832 15516 17478
rect 15580 17202 15608 17546
rect 15764 17270 15792 18634
rect 15844 18624 15896 18630
rect 16592 18612 16620 19110
rect 16868 18834 16896 19314
rect 16856 18828 16908 18834
rect 16908 18788 16988 18816
rect 16856 18770 16908 18776
rect 15844 18566 15896 18572
rect 16408 18584 16620 18612
rect 15856 18222 15884 18566
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15580 16561 15608 17138
rect 15764 16658 15792 17206
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15566 16552 15622 16561
rect 15566 16487 15622 16496
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15672 15434 15700 16186
rect 15764 15978 15792 16594
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15764 15570 15792 15914
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 13190 15608 13874
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15436 12804 15516 12832
rect 15384 12786 15436 12792
rect 15396 12434 15424 12786
rect 15580 12753 15608 13126
rect 15566 12744 15622 12753
rect 15566 12679 15622 12688
rect 15672 12434 15700 15370
rect 15764 15094 15792 15506
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15856 14532 15884 18158
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 15745 15976 16390
rect 15934 15736 15990 15745
rect 15934 15671 15990 15680
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 15304 12406 15424 12434
rect 15488 12406 15700 12434
rect 15764 14504 15884 14532
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15304 11898 15332 12406
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 10606 15056 11494
rect 15212 11354 15240 11698
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 10742 15332 11494
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10282 15240 10406
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15120 10254 15240 10282
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14936 9518 14964 10202
rect 15028 9994 15056 10202
rect 15120 10062 15148 10254
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9722 15148 9862
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15106 9616 15162 9625
rect 15106 9551 15162 9560
rect 15120 9518 15148 9551
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14660 7296 14780 7324
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 5545 14596 7142
rect 14660 6254 14688 7296
rect 14844 6866 14872 9386
rect 14936 9178 14964 9454
rect 15120 9178 15148 9454
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8430 14964 8842
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14936 6746 14964 8366
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 7546 15056 8298
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15120 7478 15148 8434
rect 15212 8129 15240 10066
rect 15198 8120 15254 8129
rect 15198 8055 15254 8064
rect 15304 7936 15332 10678
rect 15396 8090 15424 11562
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15304 7908 15424 7936
rect 15198 7848 15254 7857
rect 15198 7783 15254 7792
rect 15292 7812 15344 7818
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15212 7342 15240 7783
rect 15292 7754 15344 7760
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15304 6984 15332 7754
rect 14752 6718 14964 6746
rect 15120 6956 15332 6984
rect 15016 6724 15068 6730
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14554 5536 14610 5545
rect 14554 5471 14610 5480
rect 14660 4690 14688 6190
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14384 2746 14504 2774
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 14200 800 14228 2518
rect 14384 2417 14412 2746
rect 14568 2650 14596 4422
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14660 3505 14688 4082
rect 14752 4049 14780 6718
rect 15016 6666 15068 6672
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6186 14872 6598
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14844 5370 14872 6122
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14936 4214 14964 5510
rect 15028 5370 15056 6666
rect 15120 6390 15148 6956
rect 15198 6896 15254 6905
rect 15198 6831 15200 6840
rect 15252 6831 15254 6840
rect 15200 6802 15252 6808
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15212 6254 15240 6802
rect 15396 6610 15424 7908
rect 15304 6582 15424 6610
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15106 5944 15162 5953
rect 15106 5879 15162 5888
rect 15120 5710 15148 5879
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15198 5672 15254 5681
rect 15198 5607 15254 5616
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15014 5264 15070 5273
rect 15014 5199 15070 5208
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14738 4040 14794 4049
rect 14738 3975 14794 3984
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14844 3913 14872 3946
rect 14830 3904 14886 3913
rect 14830 3839 14886 3848
rect 15028 3777 15056 5199
rect 15212 5166 15240 5607
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4752 15160 4758
rect 15106 4720 15108 4729
rect 15160 4720 15162 4729
rect 15106 4655 15162 4664
rect 15014 3768 15070 3777
rect 15014 3703 15070 3712
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3194 14872 3334
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14370 2408 14426 2417
rect 14370 2343 14426 2352
rect 14660 2038 14688 2586
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14648 2032 14700 2038
rect 14648 1974 14700 1980
rect 14752 800 14780 2246
rect 14936 1970 14964 3538
rect 15212 3126 15240 4966
rect 15304 4690 15332 6582
rect 15382 6488 15438 6497
rect 15382 6423 15438 6432
rect 15396 6089 15424 6423
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 15488 5250 15516 12406
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15580 11898 15608 12242
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 11626 15608 11834
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15764 11218 15792 14504
rect 16132 14482 16160 15030
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 14074 15976 14214
rect 16132 14074 16160 14418
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16132 13938 16160 14010
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15842 12744 15898 12753
rect 15842 12679 15898 12688
rect 15856 12050 15884 12679
rect 15856 12022 15976 12050
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15856 11082 15884 11834
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10554 15792 10950
rect 15672 10526 15792 10554
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9722 15608 9862
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15672 9586 15700 10526
rect 15750 10296 15806 10305
rect 15750 10231 15806 10240
rect 15764 10130 15792 10231
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 8129 15608 9454
rect 15672 9178 15700 9522
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15566 8120 15622 8129
rect 15566 8055 15622 8064
rect 15672 7750 15700 8191
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 7002 15608 7346
rect 15672 7041 15700 7686
rect 15658 7032 15714 7041
rect 15568 6996 15620 7002
rect 15658 6967 15714 6976
rect 15568 6938 15620 6944
rect 15566 6624 15622 6633
rect 15566 6559 15622 6568
rect 15580 5681 15608 6559
rect 15764 5778 15792 8026
rect 15856 6662 15884 11018
rect 15948 8090 15976 12022
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16040 7834 16068 13466
rect 16132 13462 16160 13874
rect 16224 13734 16252 16458
rect 16316 15065 16344 18090
rect 16408 17610 16436 18584
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16960 18426 16988 18788
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16868 18306 16896 18362
rect 16868 18278 16988 18306
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 16794 16712 17138
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16500 15706 16528 16050
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16592 15434 16620 15982
rect 16868 15858 16896 16186
rect 16960 16114 16988 18278
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16960 16017 16988 16050
rect 16946 16008 17002 16017
rect 16946 15943 17002 15952
rect 16868 15830 16988 15858
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15162 16436 15302
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16302 15056 16358 15065
rect 16302 14991 16358 15000
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16120 13456 16172 13462
rect 16120 13398 16172 13404
rect 16132 12986 16160 13398
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 12850 16160 12922
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 12442 16160 12786
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16132 12306 16160 12378
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 10538 16160 12038
rect 16408 11937 16436 14962
rect 16960 14770 16988 15830
rect 17052 14890 17080 19722
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17144 18329 17172 18362
rect 17130 18320 17186 18329
rect 17130 18255 17186 18264
rect 17236 17882 17264 20402
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 16960 14742 17080 14770
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16762 13424 16818 13433
rect 16762 13359 16818 13368
rect 16776 13326 16804 13359
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16856 12232 16908 12238
rect 16854 12200 16856 12209
rect 16908 12200 16910 12209
rect 16854 12135 16910 12144
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16394 11928 16450 11937
rect 16544 11931 16852 11940
rect 16394 11863 16450 11872
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 10742 16252 11494
rect 16408 11354 16436 11698
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10849 16344 10950
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16302 10840 16358 10849
rect 16544 10843 16852 10852
rect 16960 10810 16988 14282
rect 16302 10775 16358 10784
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16212 10736 16264 10742
rect 16212 10678 16264 10684
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16394 10432 16450 10441
rect 16394 10367 16450 10376
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16120 9376 16172 9382
rect 16118 9344 16120 9353
rect 16172 9344 16174 9353
rect 16118 9279 16174 9288
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8673 16160 8774
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7954 16160 8230
rect 16224 8072 16252 9998
rect 16304 9920 16356 9926
rect 16408 9897 16436 10367
rect 16684 10266 16712 10610
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16960 10198 16988 10610
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 17052 10010 17080 14742
rect 17144 11762 17172 17546
rect 17224 17536 17276 17542
rect 17222 17504 17224 17513
rect 17316 17536 17368 17542
rect 17276 17504 17278 17513
rect 17316 17478 17368 17484
rect 17222 17439 17278 17448
rect 17328 17338 17356 17478
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17420 17270 17448 17818
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17236 15162 17264 17138
rect 17328 15910 17356 17138
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17144 10810 17172 11562
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17130 10160 17186 10169
rect 17130 10095 17186 10104
rect 17144 10062 17172 10095
rect 16960 9982 17080 10010
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 16304 9862 16356 9868
rect 16394 9888 16450 9897
rect 16316 8634 16344 9862
rect 16394 9823 16450 9832
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16578 9480 16634 9489
rect 16578 9415 16634 9424
rect 16592 9217 16620 9415
rect 16684 9382 16712 9658
rect 16960 9602 16988 9982
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9722 17080 9862
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16868 9574 16988 9602
rect 16868 9518 16896 9574
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16578 9208 16634 9217
rect 16578 9143 16634 9152
rect 16868 9058 16896 9454
rect 16960 9217 16988 9454
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16946 9208 17002 9217
rect 16946 9143 17002 9152
rect 16776 9042 16896 9058
rect 16764 9036 16896 9042
rect 16816 9030 16896 9036
rect 16764 8978 16816 8984
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8634 16988 8774
rect 17052 8634 17080 9318
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16224 8044 16344 8072
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 15948 7806 16068 7834
rect 15948 7342 15976 7806
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16040 6798 16068 7686
rect 16132 7546 16160 7686
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16132 6746 16160 7346
rect 16224 6866 16252 7890
rect 16316 7426 16344 8044
rect 17144 7818 17172 9386
rect 17236 8430 17264 14758
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 12434 17448 13942
rect 17328 12406 17448 12434
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17236 7857 17264 7890
rect 17222 7848 17278 7857
rect 17132 7812 17184 7818
rect 17222 7783 17278 7792
rect 17132 7754 17184 7760
rect 16946 7712 17002 7721
rect 16544 7644 16852 7653
rect 16946 7647 17002 7656
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16960 7546 16988 7647
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16316 7398 16436 7426
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16132 6718 16252 6746
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 16118 6352 16174 6361
rect 15936 6316 15988 6322
rect 16118 6287 16174 6296
rect 15936 6258 15988 6264
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15566 5672 15622 5681
rect 15566 5607 15622 5616
rect 15580 5574 15608 5607
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15488 5222 15608 5250
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15474 5128 15530 5137
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4282 15332 4422
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15396 4078 15424 5102
rect 15474 5063 15530 5072
rect 15488 4622 15516 5063
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15488 4282 15516 4558
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15396 3602 15424 4014
rect 15580 3670 15608 5222
rect 15764 4690 15792 5714
rect 15856 4690 15884 6054
rect 15948 5914 15976 6258
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15934 5400 15990 5409
rect 16040 5386 16068 6054
rect 16132 5574 16160 6287
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15990 5358 16068 5386
rect 16132 5370 16160 5510
rect 16120 5364 16172 5370
rect 15934 5335 15990 5344
rect 15948 5234 15976 5335
rect 16120 5306 16172 5312
rect 16026 5264 16082 5273
rect 15936 5228 15988 5234
rect 16026 5199 16082 5208
rect 15936 5170 15988 5176
rect 16040 5030 16068 5199
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15764 4486 15792 4626
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15658 4312 15714 4321
rect 15658 4247 15714 4256
rect 15672 4078 15700 4247
rect 15948 4146 15976 4762
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15474 3496 15530 3505
rect 15474 3431 15530 3440
rect 15488 3398 15516 3431
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15304 3194 15332 3334
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15580 2990 15608 3606
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15672 2922 15700 3334
rect 15948 3126 15976 3878
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16224 2922 16252 6718
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16316 5846 16344 6258
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16408 5778 16436 7398
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 7002 16988 7278
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17222 6896 17278 6905
rect 17328 6866 17356 12406
rect 17498 12336 17554 12345
rect 17498 12271 17554 12280
rect 17512 11762 17540 12271
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17604 11336 17632 16526
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16046 17724 16390
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17788 15706 17816 20402
rect 18064 20058 18092 22200
rect 18616 20602 18644 22200
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18234 20496 18290 20505
rect 18234 20431 18290 20440
rect 18512 20460 18564 20466
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17972 19825 18000 19994
rect 18156 19990 18184 20266
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17958 19816 18014 19825
rect 17958 19751 18014 19760
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17972 18714 18000 18906
rect 18064 18873 18092 19858
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18050 18864 18106 18873
rect 18050 18799 18106 18808
rect 17972 18686 18092 18714
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17868 18352 17920 18358
rect 17972 18329 18000 18566
rect 17868 18294 17920 18300
rect 17958 18320 18014 18329
rect 17880 17678 17908 18294
rect 17958 18255 18014 18264
rect 18064 18170 18092 18686
rect 17972 18142 18092 18170
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 16182 17908 17614
rect 17972 16998 18000 18142
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17610 18092 18022
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17696 14793 17724 14962
rect 17682 14784 17738 14793
rect 17682 14719 17738 14728
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 11898 17724 13262
rect 17788 12434 17816 15370
rect 18156 15162 18184 19790
rect 18248 19174 18276 20431
rect 18512 20402 18564 20408
rect 18326 19272 18382 19281
rect 18326 19207 18382 19216
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 15706 18276 18702
rect 18340 18154 18368 19207
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18432 18630 18460 18663
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18418 17640 18474 17649
rect 18418 17575 18474 17584
rect 18432 17338 18460 17575
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18524 17134 18552 20402
rect 19168 20330 19196 22200
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18616 17542 18644 19110
rect 18708 18766 18736 20198
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19614 20088 19670 20097
rect 19614 20023 19670 20032
rect 18878 19952 18934 19961
rect 18878 19887 18934 19896
rect 18892 19854 18920 19887
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 18193 18736 18566
rect 18694 18184 18750 18193
rect 18694 18119 18750 18128
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 16522 18552 16934
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18248 15065 18276 15098
rect 18328 15088 18380 15094
rect 18234 15056 18290 15065
rect 18144 15020 18196 15026
rect 18328 15030 18380 15036
rect 18234 14991 18290 15000
rect 18144 14962 18196 14968
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 14006 17908 14214
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 13161 17908 13194
rect 17866 13152 17922 13161
rect 17866 13087 17922 13096
rect 17972 12753 18000 14554
rect 18156 12918 18184 14962
rect 18340 14521 18368 15030
rect 18326 14512 18382 14521
rect 18326 14447 18382 14456
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13841 18276 14214
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 17958 12744 18014 12753
rect 17958 12679 18014 12688
rect 17788 12406 18000 12434
rect 17774 12336 17830 12345
rect 17774 12271 17830 12280
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17788 11694 17816 12271
rect 17972 12102 18000 12406
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 18248 11898 18276 12786
rect 18340 12186 18368 14010
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 18432 13297 18460 13398
rect 18418 13288 18474 13297
rect 18418 13223 18474 13232
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 12442 18460 12786
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18340 12170 18460 12186
rect 18340 12164 18472 12170
rect 18340 12158 18420 12164
rect 18420 12106 18472 12112
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18064 11801 18092 11834
rect 18050 11792 18106 11801
rect 17960 11756 18012 11762
rect 18050 11727 18106 11736
rect 18236 11756 18288 11762
rect 17960 11698 18012 11704
rect 18236 11698 18288 11704
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17420 11308 17632 11336
rect 17420 9110 17448 11308
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17512 10674 17540 11183
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17590 10704 17646 10713
rect 17500 10668 17552 10674
rect 17590 10639 17646 10648
rect 17500 10610 17552 10616
rect 17498 10296 17554 10305
rect 17604 10266 17632 10639
rect 17696 10470 17724 10950
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17498 10231 17554 10240
rect 17592 10260 17644 10266
rect 17512 9466 17540 10231
rect 17592 10202 17644 10208
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 9625 17632 9862
rect 17590 9616 17646 9625
rect 17590 9551 17646 9560
rect 17512 9438 17632 9466
rect 17498 9208 17554 9217
rect 17498 9143 17554 9152
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8634 17448 8910
rect 17512 8838 17540 9143
rect 17604 9092 17632 9438
rect 17788 9364 17816 11494
rect 17972 11354 18000 11698
rect 18248 11558 18276 11698
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18340 11286 18368 12038
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 10713 18000 11086
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18234 10840 18290 10849
rect 18340 10810 18368 10950
rect 18234 10775 18290 10784
rect 18328 10804 18380 10810
rect 17958 10704 18014 10713
rect 17958 10639 18014 10648
rect 17972 10130 18000 10639
rect 18248 10606 18276 10775
rect 18328 10746 18380 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 10010 18092 10066
rect 17972 9982 18092 10010
rect 17972 9722 18000 9982
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17788 9336 17908 9364
rect 17604 9064 17724 9092
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17420 7750 17448 8366
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17420 7002 17448 7686
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17406 6896 17462 6905
rect 17222 6831 17278 6840
rect 17316 6860 17368 6866
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16762 6352 16818 6361
rect 16960 6338 16988 6598
rect 16762 6287 16818 6296
rect 16868 6310 16988 6338
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16500 5556 16528 6054
rect 16776 5953 16804 6287
rect 16762 5944 16818 5953
rect 16762 5879 16818 5888
rect 16408 5528 16528 5556
rect 16868 5556 16896 6310
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5914 16988 6190
rect 17236 6186 17264 6831
rect 17406 6831 17462 6840
rect 17316 6802 17368 6808
rect 17420 6254 17448 6831
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17236 5710 17264 6122
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 16868 5528 17080 5556
rect 16408 5302 16436 5528
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16684 5234 16712 5306
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16316 3398 16344 5170
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16408 4146 16436 5034
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4622 16988 4966
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16960 4282 16988 4422
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16580 4208 16632 4214
rect 17052 4185 17080 5528
rect 17406 5128 17462 5137
rect 17406 5063 17462 5072
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16580 4150 16632 4156
rect 17038 4176 17094 4185
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16592 3534 16620 4150
rect 17038 4111 17094 4120
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16684 3602 16712 3878
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17144 3058 17172 4422
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2990 17264 3946
rect 17420 3777 17448 5063
rect 17406 3768 17462 3777
rect 17406 3703 17462 3712
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17328 3398 17356 3538
rect 17420 3534 17448 3703
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17316 3392 17368 3398
rect 17512 3380 17540 8774
rect 17590 8664 17646 8673
rect 17590 8599 17592 8608
rect 17644 8599 17646 8608
rect 17592 8570 17644 8576
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17604 8090 17632 8434
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7546 17632 7686
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17696 7410 17724 9064
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 8809 17816 8978
rect 17774 8800 17830 8809
rect 17774 8735 17830 8744
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5030 17632 6394
rect 17682 5944 17738 5953
rect 17682 5879 17738 5888
rect 17696 5778 17724 5879
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4826 17632 4966
rect 17696 4826 17724 5170
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17316 3334 17368 3340
rect 17420 3352 17540 3380
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 15108 2440 15160 2446
rect 15212 2428 15240 2790
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 15160 2400 15240 2428
rect 15108 2382 15160 2388
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 15304 800 15332 2518
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 800 15884 2246
rect 16040 2106 16068 2518
rect 16684 2446 16712 2790
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16028 2100 16080 2106
rect 16028 2042 16080 2048
rect 16408 800 16436 2314
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 800 16988 2586
rect 17236 2446 17264 2790
rect 17420 2553 17448 3352
rect 17604 3058 17632 4422
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 4049 17724 4082
rect 17682 4040 17738 4049
rect 17788 4010 17816 6734
rect 17880 5166 17908 9336
rect 17972 9110 18000 9386
rect 18248 9217 18276 10542
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18234 9208 18290 9217
rect 18234 9143 18290 9152
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 17958 8936 18014 8945
rect 17958 8871 18014 8880
rect 17972 8838 18000 8871
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 18156 8634 18184 9046
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 6458 18000 8434
rect 18142 8392 18198 8401
rect 18142 8327 18198 8336
rect 18050 7712 18106 7721
rect 18050 7647 18106 7656
rect 18064 7478 18092 7647
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6866 18092 7278
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17866 4992 17922 5001
rect 17866 4927 17922 4936
rect 17880 4457 17908 4927
rect 17972 4554 18000 5199
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17866 4448 17922 4457
rect 17866 4383 17922 4392
rect 17682 3975 17738 3984
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17500 2576 17552 2582
rect 17406 2544 17462 2553
rect 17500 2518 17552 2524
rect 17406 2479 17462 2488
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17052 2038 17080 2382
rect 17040 2032 17092 2038
rect 17040 1974 17092 1980
rect 17512 800 17540 2518
rect 17696 2514 17724 3878
rect 17958 3632 18014 3641
rect 17958 3567 17960 3576
rect 18012 3567 18014 3576
rect 17960 3538 18012 3544
rect 18064 3505 18092 6598
rect 18156 5642 18184 8327
rect 18248 8265 18276 8774
rect 18234 8256 18290 8265
rect 18234 8191 18290 8200
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18248 7546 18276 7754
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6361 18276 6598
rect 18234 6352 18290 6361
rect 18234 6287 18290 6296
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18248 5817 18276 6190
rect 18234 5808 18290 5817
rect 18234 5743 18290 5752
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18050 3496 18106 3505
rect 18050 3431 18106 3440
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17788 2446 17816 3334
rect 18156 3058 18184 5034
rect 18340 4690 18368 10406
rect 18432 10305 18460 12106
rect 18418 10296 18474 10305
rect 18418 10231 18474 10240
rect 18524 10130 18552 16458
rect 18616 15706 18644 17138
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18510 10024 18566 10033
rect 18510 9959 18566 9968
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18432 9178 18460 9386
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8430 18460 8978
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18524 8022 18552 9959
rect 18420 8016 18472 8022
rect 18512 8016 18564 8022
rect 18420 7958 18472 7964
rect 18510 7984 18512 7993
rect 18564 7984 18566 7993
rect 18432 7857 18460 7958
rect 18510 7919 18566 7928
rect 18418 7848 18474 7857
rect 18418 7783 18474 7792
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18432 7546 18460 7686
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18524 7002 18552 7686
rect 18616 7342 18644 15438
rect 18708 11234 18736 18022
rect 18800 12209 18828 19450
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18984 18086 19012 18226
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 16658 18920 17614
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19260 17241 19288 17478
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 19076 15502 19104 17002
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16794 19564 17478
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18892 15337 18920 15438
rect 18878 15328 18934 15337
rect 18878 15263 18934 15272
rect 19536 15094 19564 15914
rect 19628 15706 19656 20023
rect 19720 19718 19748 22200
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19708 19440 19760 19446
rect 19708 19382 19760 19388
rect 19720 18630 19748 19382
rect 19812 18698 19840 19722
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18786 12200 18842 12209
rect 18786 12135 18842 12144
rect 18984 12102 19012 13874
rect 19076 13530 19104 14962
rect 19614 14920 19670 14929
rect 19614 14855 19670 14864
rect 19524 14816 19576 14822
rect 19522 14784 19524 14793
rect 19576 14784 19578 14793
rect 19143 14716 19451 14725
rect 19522 14719 19578 14728
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 13977 19288 14214
rect 19246 13968 19302 13977
rect 19246 13903 19302 13912
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11676 19012 12038
rect 18892 11648 19012 11676
rect 18708 11206 18828 11234
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 10810 18736 11018
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 10062 18736 10610
rect 18800 10538 18828 11206
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18708 9625 18736 9658
rect 18694 9616 18750 9625
rect 18694 9551 18750 9560
rect 18800 9178 18828 10474
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18786 8800 18842 8809
rect 18786 8735 18842 8744
rect 18694 7984 18750 7993
rect 18694 7919 18696 7928
rect 18748 7919 18750 7928
rect 18696 7890 18748 7896
rect 18800 7834 18828 8735
rect 18708 7806 18828 7834
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 5817 18460 6258
rect 18604 6112 18656 6118
rect 18510 6080 18566 6089
rect 18604 6054 18656 6060
rect 18510 6015 18566 6024
rect 18418 5808 18474 5817
rect 18418 5743 18474 5752
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4282 18276 4422
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18432 4214 18460 5578
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18524 3534 18552 6015
rect 18616 5681 18644 6054
rect 18602 5672 18658 5681
rect 18602 5607 18658 5616
rect 18708 3670 18736 7806
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7410 18828 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 4826 18828 6734
rect 18892 5846 18920 11648
rect 18970 11520 19026 11529
rect 18970 11455 19026 11464
rect 18984 10674 19012 11455
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18984 8922 19012 9590
rect 19076 9450 19104 12854
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19536 12442 19564 14350
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19338 11928 19394 11937
rect 19338 11863 19340 11872
rect 19392 11863 19394 11872
rect 19340 11834 19392 11840
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19168 9382 19196 9930
rect 19260 9489 19288 9998
rect 19246 9480 19302 9489
rect 19246 9415 19302 9424
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18984 8894 19104 8922
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 7478 19012 8774
rect 19076 8673 19104 8894
rect 19062 8664 19118 8673
rect 19062 8599 19118 8608
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18970 6760 19026 6769
rect 18970 6695 19026 6704
rect 18984 6322 19012 6695
rect 19076 6662 19104 8434
rect 19444 8294 19472 9046
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19536 7546 19564 11086
rect 19628 10062 19656 14855
rect 19720 10606 19748 18566
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 15026 19840 15846
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 13433 19840 14214
rect 19798 13424 19854 13433
rect 19798 13359 19854 13368
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19812 11558 19840 12786
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19628 8974 19656 9862
rect 19720 9586 19748 9862
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19720 9042 19748 9386
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19812 8514 19840 10610
rect 19904 9722 19932 16050
rect 19996 15638 20024 19722
rect 20088 16182 20116 20402
rect 20272 20398 20300 22200
rect 20350 21312 20406 21321
rect 20350 21247 20406 21256
rect 20364 20806 20392 21247
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20364 19378 20392 20742
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19854 20760 20198
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 20180 15366 20208 19314
rect 20456 18698 20484 19450
rect 20732 19310 20760 19790
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 18834 20760 19246
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20364 16454 20392 17138
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20168 15360 20220 15366
rect 20166 15328 20168 15337
rect 20220 15328 20222 15337
rect 20166 15263 20222 15272
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19996 14414 20024 15098
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19996 13938 20024 14350
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13258 20024 13670
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20272 13258 20300 13466
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20364 13138 20392 16390
rect 20272 13110 20392 13138
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 11626 20024 12582
rect 20180 11830 20208 12650
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10742 20024 10950
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 20076 10600 20128 10606
rect 20074 10568 20076 10577
rect 20128 10568 20130 10577
rect 20074 10503 20130 10512
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19982 9480 20038 9489
rect 19982 9415 20038 9424
rect 19720 8486 19840 8514
rect 19996 8498 20024 9415
rect 19984 8492 20036 8498
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19338 7440 19394 7449
rect 19536 7426 19564 7482
rect 19536 7398 19656 7426
rect 19338 7375 19340 7384
rect 19392 7375 19394 7384
rect 19340 7346 19392 7352
rect 19522 7304 19578 7313
rect 19522 7239 19578 7248
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19536 7041 19564 7239
rect 19522 7032 19578 7041
rect 19522 6967 19578 6976
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6458 19104 6598
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19168 6338 19196 6870
rect 19536 6798 19564 6967
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19246 6624 19302 6633
rect 19246 6559 19302 6568
rect 19260 6390 19288 6559
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19076 6310 19196 6338
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19524 6316 19576 6322
rect 18984 6225 19012 6258
rect 18970 6216 19026 6225
rect 18970 6151 19026 6160
rect 18972 6112 19024 6118
rect 18970 6080 18972 6089
rect 19024 6080 19026 6089
rect 18970 6015 19026 6024
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 5370 18920 5510
rect 19076 5409 19104 6310
rect 19524 6258 19576 6264
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19062 5400 19118 5409
rect 18880 5364 18932 5370
rect 19062 5335 19118 5344
rect 18880 5306 18932 5312
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18616 3466 18644 3606
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18524 3058 18552 3334
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 17880 2446 17908 2994
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18064 800 18092 2790
rect 18708 2514 18736 3334
rect 18800 2922 18828 3334
rect 18892 3194 18920 4966
rect 18984 4690 19012 5102
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19536 4758 19564 6258
rect 19628 5642 19656 7398
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19614 5400 19670 5409
rect 19614 5335 19670 5344
rect 19628 5001 19656 5335
rect 19614 4992 19670 5001
rect 19614 4927 19670 4936
rect 19720 4842 19748 8486
rect 19984 8434 20036 8440
rect 19890 8392 19946 8401
rect 19800 8356 19852 8362
rect 19890 8327 19946 8336
rect 19800 8298 19852 8304
rect 19812 6798 19840 8298
rect 19904 8090 19932 8327
rect 19982 8256 20038 8265
rect 19982 8191 20038 8200
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19996 7410 20024 8191
rect 20088 7886 20116 10406
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19996 6662 20024 6695
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19812 5302 19840 5510
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19904 5166 19932 5782
rect 20180 5778 20208 11766
rect 20272 9654 20300 13110
rect 20456 11218 20484 18634
rect 20824 17270 20852 22200
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19417 20944 19790
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20902 19408 20958 19417
rect 20902 19343 20958 19352
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16697 20576 17138
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20534 16688 20590 16697
rect 20534 16623 20590 16632
rect 20640 16561 20668 16934
rect 20812 16584 20864 16590
rect 20626 16552 20682 16561
rect 20812 16526 20864 16532
rect 20626 16487 20682 16496
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15609 20760 15846
rect 20718 15600 20774 15609
rect 20718 15535 20774 15544
rect 20824 14498 20852 16526
rect 20732 14470 20852 14498
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20272 9518 20300 9590
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 20364 9178 20392 11018
rect 20456 10538 20484 11154
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20548 9738 20576 13262
rect 20640 12918 20668 14010
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10130 20668 10950
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20456 9710 20576 9738
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20272 8090 20300 8502
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20258 7848 20314 7857
rect 20258 7783 20314 7792
rect 20272 6798 20300 7783
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20364 6458 20392 8434
rect 20456 7546 20484 9710
rect 20732 9110 20760 14470
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20824 10266 20852 14010
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9761 20852 9930
rect 20810 9752 20866 9761
rect 20810 9687 20866 9696
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20640 8634 20668 8842
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20732 7886 20760 8774
rect 20810 8528 20866 8537
rect 20810 8463 20866 8472
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20442 7440 20498 7449
rect 20442 7375 20498 7384
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 6322 20484 7375
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20640 5710 20668 6054
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20732 5642 20760 7142
rect 20824 6798 20852 8463
rect 20916 7546 20944 18702
rect 21008 18358 21036 19654
rect 21376 18970 21404 22200
rect 21560 19174 21588 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21284 18290 21312 18770
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21100 17610 21128 18022
rect 21284 17678 21312 18226
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 21008 14498 21036 17546
rect 21284 17134 21312 17614
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21100 14822 21128 15370
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21008 14470 21128 14498
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21008 13326 21036 14282
rect 21100 14074 21128 14470
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21100 11286 21128 13670
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 21008 8838 21036 11086
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21100 9994 21128 10746
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 21086 9888 21142 9897
rect 21086 9823 21142 9832
rect 21100 9722 21128 9823
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21192 9450 21220 16050
rect 21284 15502 21312 17070
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16017 21404 16934
rect 21468 16833 21496 18566
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21454 16824 21510 16833
rect 21454 16759 21510 16768
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21362 16008 21418 16017
rect 21362 15943 21418 15952
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 14414 21312 15438
rect 21272 14408 21324 14414
rect 21376 14385 21404 15846
rect 21468 15065 21496 16390
rect 21454 15056 21510 15065
rect 21454 14991 21510 15000
rect 21560 14906 21588 18294
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21468 14878 21588 14906
rect 21272 14350 21324 14356
rect 21362 14376 21418 14385
rect 21284 13818 21312 14350
rect 21362 14311 21418 14320
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21376 13818 21404 13874
rect 21284 13790 21404 13818
rect 21284 13394 21312 13790
rect 21362 13560 21418 13569
rect 21362 13495 21364 13504
rect 21416 13495 21418 13504
rect 21364 13466 21416 13472
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21284 12850 21312 13330
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 12238 21312 12786
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11762 21312 12174
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 11218 21312 11698
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21284 10266 21312 11154
rect 21376 11082 21404 11834
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20996 8832 21048 8838
rect 21048 8792 21220 8820
rect 20996 8774 21048 8780
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21008 6866 21036 8434
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 21008 6458 21036 6802
rect 21100 6458 21128 8502
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20628 5568 20680 5574
rect 21100 5545 21128 6190
rect 21192 5710 21220 8792
rect 21284 8090 21312 10202
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21376 9586 21404 10134
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21362 9072 21418 9081
rect 21362 9007 21418 9016
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21376 6798 21404 9007
rect 21468 8430 21496 14878
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 11558 21588 14282
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20628 5510 20680 5516
rect 21086 5536 21142 5545
rect 19982 5400 20038 5409
rect 19982 5335 19984 5344
rect 20036 5335 20038 5344
rect 19984 5306 20036 5312
rect 20272 5302 20300 5510
rect 20548 5370 20576 5510
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 19800 5160 19852 5166
rect 19798 5128 19800 5137
rect 19892 5160 19944 5166
rect 19852 5128 19854 5137
rect 19892 5102 19944 5108
rect 19798 5063 19854 5072
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 19720 4814 19840 4842
rect 19812 4758 19840 4814
rect 19524 4752 19576 4758
rect 19154 4720 19210 4729
rect 18972 4684 19024 4690
rect 19524 4694 19576 4700
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19154 4655 19210 4664
rect 18972 4626 19024 4632
rect 19168 4622 19196 4655
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19246 4584 19302 4593
rect 19246 4519 19248 4528
rect 19300 4519 19302 4528
rect 19248 4490 19300 4496
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3738 19012 4082
rect 20364 4078 20392 4966
rect 20640 4690 20668 5510
rect 21086 5471 21142 5480
rect 21560 5166 21588 11494
rect 21652 8022 21680 17138
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 22112 14056 22140 17546
rect 22020 14028 22140 14056
rect 22020 13734 22048 14028
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 22112 10810 22140 13806
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22006 10296 22062 10305
rect 22062 10254 22140 10282
rect 22006 10231 22062 10240
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 22112 9722 22140 10254
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22006 9616 22062 9625
rect 22204 9602 22232 18362
rect 22480 17882 22508 22200
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22388 12170 22416 15302
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22062 9574 22232 9602
rect 22006 9551 22062 9560
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 22296 7410 22324 9658
rect 22388 7562 22416 12106
rect 22480 7750 22508 14758
rect 22572 12434 22600 18634
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22572 12406 22692 12434
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22572 9654 22600 11018
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22664 8362 22692 12406
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22388 7534 22600 7562
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20626 4448 20682 4457
rect 20626 4383 20682 4392
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 800 18644 2246
rect 18892 1737 18920 2994
rect 18970 2544 19026 2553
rect 18970 2479 19026 2488
rect 18984 2378 19012 2479
rect 19076 2378 19104 3878
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19168 3194 19196 3606
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19444 2961 19472 3470
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19156 2576 19208 2582
rect 20180 2553 20208 3402
rect 20260 2576 20312 2582
rect 19156 2518 19208 2524
rect 20166 2544 20222 2553
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 18878 1728 18934 1737
rect 18878 1663 18934 1672
rect 19168 800 19196 2518
rect 20260 2518 20312 2524
rect 20166 2479 20222 2488
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19708 2304 19760 2310
rect 19708 2246 19760 2252
rect 19720 800 19748 2246
rect 19812 2106 19840 2382
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 20272 800 20300 2518
rect 20456 2038 20484 4150
rect 20640 4146 20668 4383
rect 20732 4185 20760 4558
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 20718 4176 20774 4185
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20628 4140 20680 4146
rect 20718 4111 20774 4120
rect 20628 4082 20680 4088
rect 20548 4049 20576 4082
rect 20534 4040 20590 4049
rect 20534 3975 20590 3984
rect 22468 4004 22520 4010
rect 20548 3777 20576 3975
rect 22468 3946 22520 3952
rect 20534 3768 20590 3777
rect 20534 3703 20590 3712
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 20536 3528 20588 3534
rect 20534 3496 20536 3505
rect 20588 3496 20590 3505
rect 20534 3431 20590 3440
rect 20534 3088 20590 3097
rect 20534 3023 20536 3032
rect 20588 3023 20590 3032
rect 20536 2994 20588 3000
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20444 2032 20496 2038
rect 20442 2000 20444 2009
rect 20496 2000 20498 2009
rect 20442 1935 20498 1944
rect 20456 1909 20484 1935
rect 20824 800 20852 2790
rect 21376 800 21404 2858
rect 11072 734 11376 762
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21560 762 21588 3606
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21836 870 21956 898
rect 21836 762 21864 870
rect 21928 800 21956 870
rect 22480 800 22508 3946
rect 22572 2774 22600 7534
rect 22756 6254 22784 11562
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22940 5098 22968 12854
rect 22928 5092 22980 5098
rect 22928 5034 22980 5040
rect 22572 2746 22692 2774
rect 22664 1970 22692 2746
rect 22652 1964 22704 1970
rect 22652 1906 22704 1912
rect 21560 734 21864 762
rect 21914 0 21970 800
rect 22466 0 22522 800
<< via2 >>
rect 1490 17176 1546 17232
rect 2042 17740 2098 17776
rect 2042 17720 2044 17740
rect 2044 17720 2096 17740
rect 2096 17720 2098 17740
rect 1950 16632 2006 16688
rect 3146 19896 3202 19952
rect 2778 17040 2834 17096
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 4158 20032 4214 20088
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3146 12688 3202 12744
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 2134 11192 2190 11248
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 4342 19760 4398 19816
rect 4342 19080 4398 19136
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 1582 6180 1638 6216
rect 1582 6160 1584 6180
rect 1584 6160 1636 6180
rect 1636 6160 1638 6180
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 1398 5752 1454 5808
rect 4434 18708 4436 18728
rect 4436 18708 4488 18728
rect 4488 18708 4490 18728
rect 4434 18672 4490 18708
rect 4618 15308 4620 15328
rect 4620 15308 4672 15328
rect 4672 15308 4674 15328
rect 4618 15272 4674 15308
rect 5722 20440 5778 20496
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 5538 19216 5594 19272
rect 5630 16904 5686 16960
rect 6826 20304 6882 20360
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6642 19352 6698 19408
rect 5354 13912 5410 13968
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4710 7248 4766 7304
rect 5722 12708 5778 12744
rect 5722 12688 5724 12708
rect 5724 12688 5776 12708
rect 5776 12688 5778 12708
rect 5538 11076 5594 11112
rect 5538 11056 5540 11076
rect 5540 11056 5592 11076
rect 5592 11056 5594 11076
rect 5354 9152 5410 9208
rect 5078 4120 5134 4176
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5722 9424 5778 9480
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6366 15408 6422 15464
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 7010 20168 7066 20224
rect 7194 20032 7250 20088
rect 6918 19624 6974 19680
rect 7102 19624 7158 19680
rect 6918 19292 6974 19348
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6550 13812 6552 13832
rect 6552 13812 6604 13832
rect 6604 13812 6606 13832
rect 6550 13776 6606 13812
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 7286 19488 7342 19544
rect 7194 19352 7250 19408
rect 7378 19352 7434 19408
rect 7746 19488 7802 19544
rect 8114 19624 8170 19680
rect 7930 19352 7986 19408
rect 7654 19080 7710 19136
rect 7746 17620 7748 17640
rect 7748 17620 7800 17640
rect 7800 17620 7802 17640
rect 7746 17584 7802 17620
rect 7286 8472 7342 8528
rect 6826 8336 6882 8392
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5998 6704 6054 6760
rect 5722 3168 5778 3224
rect 5630 2624 5686 2680
rect 5630 2352 5686 2408
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7470 6160 7526 6216
rect 8022 11056 8078 11112
rect 7930 9152 7986 9208
rect 8574 14884 8630 14920
rect 8574 14864 8576 14884
rect 8576 14864 8628 14884
rect 8628 14864 8630 14884
rect 8390 10104 8446 10160
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 9218 19488 9274 19544
rect 9494 20032 9550 20088
rect 9126 19080 9182 19136
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9310 17176 9366 17232
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9218 15272 9274 15328
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9218 13776 9274 13832
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9310 12824 9366 12880
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8022 9016 8078 9072
rect 7838 6860 7894 6896
rect 7838 6840 7840 6860
rect 7840 6840 7892 6860
rect 7892 6840 7894 6860
rect 7286 5616 7342 5672
rect 8022 5752 8078 5808
rect 8206 8492 8262 8528
rect 8206 8472 8208 8492
rect 8208 8472 8260 8492
rect 8260 8472 8262 8492
rect 8206 7792 8262 7848
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 9954 16496 10010 16552
rect 9494 12824 9550 12880
rect 9402 10804 9458 10840
rect 9402 10784 9404 10804
rect 9404 10784 9456 10804
rect 9456 10784 9458 10804
rect 9310 9968 9366 10024
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9678 12280 9734 12336
rect 8574 7384 8630 7440
rect 8482 6840 8538 6896
rect 8206 5480 8262 5536
rect 8390 5072 8446 5128
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8666 6704 8722 6760
rect 9126 6740 9128 6760
rect 9128 6740 9180 6760
rect 9180 6740 9182 6760
rect 9126 6704 9182 6740
rect 8666 6432 8722 6488
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9218 4800 9274 4856
rect 8850 4020 8852 4040
rect 8852 4020 8904 4040
rect 8904 4020 8906 4040
rect 8850 3984 8906 4020
rect 9310 4548 9366 4584
rect 9310 4528 9312 4548
rect 9312 4528 9364 4548
rect 9364 4528 9366 4548
rect 8574 3884 8576 3904
rect 8576 3884 8628 3904
rect 8628 3884 8630 3904
rect 8574 3848 8630 3884
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8298 3032 8354 3088
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9310 2508 9366 2544
rect 9310 2488 9312 2508
rect 9312 2488 9364 2508
rect 9364 2488 9366 2508
rect 10138 11328 10194 11384
rect 10046 9560 10102 9616
rect 11150 17720 11206 17776
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11518 19372 11574 19408
rect 11518 19352 11520 19372
rect 11520 19352 11572 19372
rect 11572 19352 11574 19372
rect 11334 19080 11390 19136
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11242 17176 11298 17232
rect 12530 19080 12586 19136
rect 12898 19352 12954 19408
rect 12162 17876 12218 17912
rect 12162 17856 12164 17876
rect 12164 17856 12216 17876
rect 12216 17856 12218 17876
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11150 13232 11206 13288
rect 11058 12144 11114 12200
rect 10598 9696 10654 9752
rect 10230 5480 10286 5536
rect 9862 3984 9918 4040
rect 9770 3440 9826 3496
rect 10414 7148 10416 7168
rect 10416 7148 10468 7168
rect 10468 7148 10470 7168
rect 10414 7112 10470 7148
rect 11058 11464 11114 11520
rect 11058 8608 11114 8664
rect 10690 7248 10746 7304
rect 10506 6976 10562 7032
rect 10506 5752 10562 5808
rect 11058 7248 11114 7304
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11426 11192 11482 11248
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11794 10240 11850 10296
rect 12162 13232 12218 13288
rect 11702 9424 11758 9480
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11702 6160 11758 6216
rect 10966 4256 11022 4312
rect 11150 4120 11206 4176
rect 10506 3612 10508 3632
rect 10508 3612 10560 3632
rect 10560 3612 10562 3632
rect 10506 3576 10562 3612
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11978 8336 12034 8392
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11150 2916 11206 2952
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11150 2896 11152 2916
rect 11152 2896 11204 2916
rect 11204 2896 11206 2916
rect 12714 18300 12716 18320
rect 12716 18300 12768 18320
rect 12768 18300 12770 18320
rect 12714 18264 12770 18300
rect 12806 17856 12862 17912
rect 13542 20340 13544 20360
rect 13544 20340 13596 20360
rect 13596 20340 13598 20360
rect 13542 20304 13598 20340
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13726 20032 13782 20088
rect 12990 18536 13046 18592
rect 13266 16632 13322 16688
rect 13266 15408 13322 15464
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 14186 18536 14242 18592
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 14186 15308 14188 15328
rect 14188 15308 14240 15328
rect 14240 15308 14242 15328
rect 14186 15272 14242 15308
rect 12622 13640 12678 13696
rect 12162 10376 12218 10432
rect 12162 10240 12218 10296
rect 12162 9832 12218 9888
rect 12254 9560 12310 9616
rect 12162 9444 12218 9480
rect 12162 9424 12164 9444
rect 12164 9424 12216 9444
rect 12216 9424 12218 9444
rect 11978 6452 12034 6488
rect 11978 6432 11980 6452
rect 11980 6432 12032 6452
rect 12032 6432 12034 6452
rect 12254 8880 12310 8936
rect 13634 13912 13690 13968
rect 12714 11736 12770 11792
rect 12714 11192 12770 11248
rect 12622 11092 12624 11112
rect 12624 11092 12676 11112
rect 12676 11092 12678 11112
rect 12622 11056 12678 11092
rect 12714 9424 12770 9480
rect 11978 4664 12034 4720
rect 12622 7520 12678 7576
rect 12530 6976 12586 7032
rect 12438 5616 12494 5672
rect 12622 5616 12678 5672
rect 12898 12824 12954 12880
rect 12990 11736 13046 11792
rect 12898 10920 12954 10976
rect 13082 10784 13138 10840
rect 13082 7928 13138 7984
rect 13358 11872 13414 11928
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14186 12280 14242 12336
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13082 7248 13138 7304
rect 13266 6840 13322 6896
rect 13082 5480 13138 5536
rect 13634 9696 13690 9752
rect 13450 8880 13506 8936
rect 13726 7792 13782 7848
rect 13634 7692 13636 7712
rect 13636 7692 13688 7712
rect 13688 7692 13690 7712
rect 13634 7656 13690 7692
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13910 9968 13966 10024
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14922 18672 14978 18728
rect 15106 18708 15108 18728
rect 15108 18708 15160 18728
rect 15160 18708 15162 18728
rect 15106 18672 15162 18708
rect 14738 17620 14740 17640
rect 14740 17620 14792 17640
rect 14792 17620 14794 17640
rect 14738 17584 14794 17620
rect 14646 15952 14702 16008
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16670 20460 16726 20496
rect 16670 20440 16672 20460
rect 16672 20440 16724 20460
rect 16724 20440 16726 20460
rect 15750 19760 15806 19816
rect 17958 20868 18014 20904
rect 17958 20848 17960 20868
rect 17960 20848 18012 20868
rect 18012 20848 18014 20868
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 14462 14764 14464 14784
rect 14464 14764 14516 14784
rect 14516 14764 14518 14784
rect 14462 14728 14518 14764
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13726 7248 13782 7304
rect 13818 7112 13874 7168
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13542 5772 13598 5808
rect 13542 5752 13544 5772
rect 13544 5752 13596 5772
rect 13596 5752 13598 5772
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14646 9580 14702 9616
rect 14646 9560 14648 9580
rect 14648 9560 14700 9580
rect 14700 9560 14702 9580
rect 14370 7112 14426 7168
rect 14278 5616 14334 5672
rect 13726 5072 13782 5128
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13818 4664 13874 4720
rect 13818 3984 13874 4040
rect 14278 3984 14334 4040
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14186 3440 14242 3496
rect 15566 16496 15622 16552
rect 15566 12688 15622 12744
rect 15934 15680 15990 15736
rect 15106 9560 15162 9616
rect 15198 8064 15254 8120
rect 15198 7792 15254 7848
rect 14554 5480 14610 5536
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15198 6860 15254 6896
rect 15198 6840 15200 6860
rect 15200 6840 15252 6860
rect 15252 6840 15254 6860
rect 15106 5888 15162 5944
rect 15198 5616 15254 5672
rect 15014 5208 15070 5264
rect 14738 3984 14794 4040
rect 14830 3848 14886 3904
rect 15106 4700 15108 4720
rect 15108 4700 15160 4720
rect 15160 4700 15162 4720
rect 15106 4664 15162 4700
rect 15014 3712 15070 3768
rect 14646 3440 14702 3496
rect 14370 2352 14426 2408
rect 15382 6432 15438 6488
rect 15382 6024 15438 6080
rect 15842 12688 15898 12744
rect 15750 10240 15806 10296
rect 15658 8200 15714 8256
rect 15566 8064 15622 8120
rect 15658 6976 15714 7032
rect 15566 6568 15622 6624
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16946 15952 17002 16008
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16302 15000 16358 15056
rect 17130 18264 17186 18320
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16762 13368 16818 13424
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16854 12180 16856 12200
rect 16856 12180 16908 12200
rect 16908 12180 16910 12200
rect 16854 12144 16910 12180
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16394 11872 16450 11928
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16302 10784 16358 10840
rect 16394 10376 16450 10432
rect 16118 9324 16120 9344
rect 16120 9324 16172 9344
rect 16172 9324 16174 9344
rect 16118 9288 16174 9324
rect 16118 8608 16174 8664
rect 17222 17484 17224 17504
rect 17224 17484 17276 17504
rect 17276 17484 17278 17504
rect 17222 17448 17278 17484
rect 17130 10104 17186 10160
rect 16394 9832 16450 9888
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16578 9424 16634 9480
rect 16578 9152 16634 9208
rect 16946 9152 17002 9208
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 17222 7792 17278 7848
rect 16946 7656 17002 7712
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16118 6296 16174 6352
rect 15566 5616 15622 5672
rect 15474 5072 15530 5128
rect 15934 5344 15990 5400
rect 16026 5208 16082 5264
rect 15658 4256 15714 4312
rect 15474 3440 15530 3496
rect 17222 6840 17278 6896
rect 17498 12280 17554 12336
rect 18234 20440 18290 20496
rect 17958 19760 18014 19816
rect 18050 18808 18106 18864
rect 17958 18264 18014 18320
rect 17682 14728 17738 14784
rect 18326 19216 18382 19272
rect 18418 18672 18474 18728
rect 18418 17584 18474 17640
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19614 20032 19670 20088
rect 18878 19896 18934 19952
rect 18694 18128 18750 18184
rect 18234 15000 18290 15056
rect 17866 13096 17922 13152
rect 18326 14456 18382 14512
rect 18234 13776 18290 13832
rect 17958 12688 18014 12744
rect 17774 12280 17830 12336
rect 18418 13232 18474 13288
rect 18050 11736 18106 11792
rect 17498 11192 17554 11248
rect 17590 10648 17646 10704
rect 17498 10240 17554 10296
rect 17590 9560 17646 9616
rect 17498 9152 17554 9208
rect 18234 10784 18290 10840
rect 17958 10648 18014 10704
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16762 6296 16818 6352
rect 16762 5888 16818 5944
rect 17406 6840 17462 6896
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17406 5072 17462 5128
rect 17038 4120 17094 4176
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17406 3712 17462 3768
rect 17590 8628 17646 8664
rect 17590 8608 17592 8628
rect 17592 8608 17644 8628
rect 17644 8608 17646 8628
rect 17774 8744 17830 8800
rect 17682 5888 17738 5944
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17682 3984 17738 4040
rect 18234 9152 18290 9208
rect 17958 8880 18014 8936
rect 18142 8336 18198 8392
rect 18050 7656 18106 7712
rect 17958 5208 18014 5264
rect 17866 4936 17922 4992
rect 17866 4392 17922 4448
rect 17406 2488 17462 2544
rect 17958 3596 18014 3632
rect 17958 3576 17960 3596
rect 17960 3576 18012 3596
rect 18012 3576 18014 3596
rect 18234 8200 18290 8256
rect 18234 6296 18290 6352
rect 18234 5752 18290 5808
rect 18050 3440 18106 3496
rect 18418 10240 18474 10296
rect 18510 9968 18566 10024
rect 18510 7964 18512 7984
rect 18512 7964 18564 7984
rect 18564 7964 18566 7984
rect 18510 7928 18566 7964
rect 18418 7792 18474 7848
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19246 17176 19302 17232
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 18878 15272 18934 15328
rect 18786 12144 18842 12200
rect 19614 14864 19670 14920
rect 19522 14764 19524 14784
rect 19524 14764 19576 14784
rect 19576 14764 19578 14784
rect 19522 14728 19578 14764
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19246 13912 19302 13968
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18694 9560 18750 9616
rect 18786 8744 18842 8800
rect 18694 7948 18750 7984
rect 18694 7928 18696 7948
rect 18696 7928 18748 7948
rect 18748 7928 18750 7948
rect 18510 6024 18566 6080
rect 18418 5752 18474 5808
rect 18602 5616 18658 5672
rect 18970 11464 19026 11520
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19338 11892 19394 11928
rect 19338 11872 19340 11892
rect 19340 11872 19392 11892
rect 19392 11872 19394 11892
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19246 9424 19302 9480
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19062 8608 19118 8664
rect 18970 6704 19026 6760
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19798 13368 19854 13424
rect 20350 21256 20406 21312
rect 20166 15308 20168 15328
rect 20168 15308 20220 15328
rect 20220 15308 20222 15328
rect 20166 15272 20222 15308
rect 20074 10548 20076 10568
rect 20076 10548 20128 10568
rect 20128 10548 20130 10568
rect 20074 10512 20130 10548
rect 19982 9424 20038 9480
rect 19338 7404 19394 7440
rect 19338 7384 19340 7404
rect 19340 7384 19392 7404
rect 19392 7384 19394 7404
rect 19522 7248 19578 7304
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19522 6976 19578 7032
rect 19246 6568 19302 6624
rect 18970 6160 19026 6216
rect 18970 6060 18972 6080
rect 18972 6060 19024 6080
rect 19024 6060 19026 6080
rect 18970 6024 19026 6060
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19062 5344 19118 5400
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19614 5344 19670 5400
rect 19614 4936 19670 4992
rect 19890 8336 19946 8392
rect 19982 8200 20038 8256
rect 19982 6704 20038 6760
rect 20902 19352 20958 19408
rect 20534 16632 20590 16688
rect 20626 16496 20682 16552
rect 20718 15544 20774 15600
rect 20258 7792 20314 7848
rect 20810 9696 20866 9752
rect 20810 8472 20866 8528
rect 20442 7384 20498 7440
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21086 9832 21142 9888
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21454 16768 21510 16824
rect 21362 15952 21418 16008
rect 21454 15000 21510 15056
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21362 14320 21418 14376
rect 21362 13524 21418 13560
rect 21362 13504 21364 13524
rect 21364 13504 21416 13524
rect 21416 13504 21418 13524
rect 21362 9016 21418 9072
rect 19982 5364 20038 5400
rect 19982 5344 19984 5364
rect 19984 5344 20036 5364
rect 20036 5344 20038 5364
rect 19798 5108 19800 5128
rect 19800 5108 19852 5128
rect 19852 5108 19854 5128
rect 19798 5072 19854 5108
rect 19154 4664 19210 4720
rect 19246 4548 19302 4584
rect 19246 4528 19248 4548
rect 19248 4528 19300 4548
rect 19300 4528 19302 4548
rect 21086 5480 21142 5536
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 22006 10240 22062 10296
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 22006 9560 22062 9616
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 20626 4392 20682 4448
rect 18970 2488 19026 2544
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19430 2896 19486 2952
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 18878 1672 18934 1728
rect 20166 2488 20222 2544
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 20718 4120 20774 4176
rect 20534 3984 20590 4040
rect 20534 3712 20590 3768
rect 20534 3476 20536 3496
rect 20536 3476 20588 3496
rect 20588 3476 20590 3496
rect 20534 3440 20590 3476
rect 20534 3052 20590 3088
rect 20534 3032 20536 3052
rect 20536 3032 20588 3052
rect 20588 3032 20590 3052
rect 20442 1980 20444 2000
rect 20444 1980 20496 2000
rect 20496 1980 20498 2000
rect 20442 1944 20498 1980
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 20345 21314 20411 21317
rect 22200 21314 23000 21344
rect 20345 21312 23000 21314
rect 20345 21256 20350 21312
rect 20406 21256 23000 21312
rect 20345 21254 23000 21256
rect 20345 21251 20411 21254
rect 22200 21224 23000 21254
rect 17953 20906 18019 20909
rect 22200 20906 23000 20936
rect 17953 20904 23000 20906
rect 17953 20848 17958 20904
rect 18014 20848 23000 20904
rect 17953 20846 23000 20848
rect 17953 20843 18019 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 5717 20498 5783 20501
rect 16665 20498 16731 20501
rect 5717 20496 16731 20498
rect 5717 20440 5722 20496
rect 5778 20440 16670 20496
rect 16726 20440 16731 20496
rect 5717 20438 16731 20440
rect 5717 20435 5783 20438
rect 16665 20435 16731 20438
rect 18229 20498 18295 20501
rect 22200 20498 23000 20528
rect 18229 20496 23000 20498
rect 18229 20440 18234 20496
rect 18290 20440 23000 20496
rect 18229 20438 23000 20440
rect 18229 20435 18295 20438
rect 22200 20408 23000 20438
rect 6821 20362 6887 20365
rect 13537 20362 13603 20365
rect 6821 20360 13603 20362
rect 6821 20304 6826 20360
rect 6882 20304 13542 20360
rect 13598 20304 13603 20360
rect 6821 20302 13603 20304
rect 6821 20299 6887 20302
rect 13537 20299 13603 20302
rect 7005 20228 7071 20229
rect 7005 20224 7052 20228
rect 7116 20226 7122 20228
rect 7005 20168 7010 20224
rect 7005 20164 7052 20168
rect 7116 20166 7162 20226
rect 7116 20164 7122 20166
rect 7005 20163 7071 20164
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 4153 20090 4219 20093
rect 7189 20090 7255 20093
rect 4153 20088 7255 20090
rect 4153 20032 4158 20088
rect 4214 20032 7194 20088
rect 7250 20032 7255 20088
rect 4153 20030 7255 20032
rect 4153 20027 4219 20030
rect 7189 20027 7255 20030
rect 9489 20090 9555 20093
rect 13721 20090 13787 20093
rect 9489 20088 13787 20090
rect 9489 20032 9494 20088
rect 9550 20032 13726 20088
rect 13782 20032 13787 20088
rect 9489 20030 13787 20032
rect 9489 20027 9555 20030
rect 13721 20027 13787 20030
rect 19609 20090 19675 20093
rect 22200 20090 23000 20120
rect 19609 20088 23000 20090
rect 19609 20032 19614 20088
rect 19670 20032 23000 20088
rect 19609 20030 23000 20032
rect 19609 20027 19675 20030
rect 22200 20000 23000 20030
rect 3141 19954 3207 19957
rect 18873 19954 18939 19957
rect 3141 19952 18939 19954
rect 3141 19896 3146 19952
rect 3202 19896 18878 19952
rect 18934 19896 18939 19952
rect 3141 19894 18939 19896
rect 3141 19891 3207 19894
rect 18873 19891 18939 19894
rect 4337 19818 4403 19821
rect 15745 19818 15811 19821
rect 4337 19816 15811 19818
rect 4337 19760 4342 19816
rect 4398 19760 15750 19816
rect 15806 19760 15811 19816
rect 4337 19758 15811 19760
rect 4337 19755 4403 19758
rect 15745 19755 15811 19758
rect 17953 19818 18019 19821
rect 17953 19816 22202 19818
rect 17953 19760 17958 19816
rect 18014 19760 22202 19816
rect 17953 19758 22202 19760
rect 17953 19755 18019 19758
rect 22142 19712 22202 19758
rect 6913 19682 6979 19685
rect 6870 19680 6979 19682
rect 6870 19624 6918 19680
rect 6974 19624 6979 19680
rect 6870 19619 6979 19624
rect 7097 19682 7163 19685
rect 8109 19682 8175 19685
rect 7097 19680 8175 19682
rect 7097 19624 7102 19680
rect 7158 19624 8114 19680
rect 8170 19624 8175 19680
rect 7097 19622 8175 19624
rect 22142 19622 23000 19712
rect 7097 19619 7163 19622
rect 8109 19619 8175 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 6637 19412 6703 19413
rect 6637 19410 6684 19412
rect 5582 19408 6684 19410
rect 5582 19352 6642 19408
rect 5582 19350 6684 19352
rect 5582 19277 5642 19350
rect 6637 19348 6684 19350
rect 6748 19348 6754 19412
rect 6870 19353 6930 19619
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 7281 19546 7347 19549
rect 7741 19546 7807 19549
rect 9213 19546 9279 19549
rect 7281 19544 9279 19546
rect 7281 19488 7286 19544
rect 7342 19488 7746 19544
rect 7802 19488 9218 19544
rect 9274 19488 9279 19544
rect 7281 19486 9279 19488
rect 7281 19483 7347 19486
rect 7741 19483 7807 19486
rect 9213 19483 9279 19486
rect 6870 19348 6979 19353
rect 7046 19348 7052 19412
rect 7116 19410 7122 19412
rect 7189 19410 7255 19413
rect 7116 19408 7255 19410
rect 7116 19352 7194 19408
rect 7250 19352 7255 19408
rect 7116 19350 7255 19352
rect 7116 19348 7122 19350
rect 6637 19347 6703 19348
rect 6870 19292 6918 19348
rect 6974 19292 6979 19348
rect 7189 19347 7255 19350
rect 7373 19412 7439 19413
rect 7925 19412 7991 19413
rect 7373 19408 7420 19412
rect 7484 19410 7490 19412
rect 7373 19352 7378 19408
rect 7373 19348 7420 19352
rect 7484 19350 7530 19410
rect 7925 19408 7972 19412
rect 8036 19410 8042 19412
rect 7925 19352 7930 19408
rect 7484 19348 7490 19350
rect 7925 19348 7972 19352
rect 8036 19350 8082 19410
rect 8036 19348 8042 19350
rect 10726 19348 10732 19412
rect 10796 19410 10802 19412
rect 11513 19410 11579 19413
rect 10796 19408 11579 19410
rect 10796 19352 11518 19408
rect 11574 19352 11579 19408
rect 10796 19350 11579 19352
rect 10796 19348 10802 19350
rect 7373 19347 7439 19348
rect 7925 19347 7991 19348
rect 11513 19347 11579 19350
rect 12893 19410 12959 19413
rect 20897 19410 20963 19413
rect 12893 19408 20963 19410
rect 12893 19352 12898 19408
rect 12954 19352 20902 19408
rect 20958 19352 20963 19408
rect 12893 19350 20963 19352
rect 12893 19347 12959 19350
rect 20897 19347 20963 19350
rect 6870 19290 6979 19292
rect 6913 19287 6979 19290
rect 5533 19272 5642 19277
rect 5533 19216 5538 19272
rect 5594 19216 5642 19272
rect 5533 19214 5642 19216
rect 18321 19274 18387 19277
rect 22200 19274 23000 19304
rect 18321 19272 23000 19274
rect 18321 19216 18326 19272
rect 18382 19216 23000 19272
rect 18321 19214 23000 19216
rect 5533 19211 5599 19214
rect 18321 19211 18387 19214
rect 22200 19184 23000 19214
rect 4337 19138 4403 19141
rect 7649 19138 7715 19141
rect 4337 19136 7715 19138
rect 4337 19080 4342 19136
rect 4398 19080 7654 19136
rect 7710 19080 7715 19136
rect 4337 19078 7715 19080
rect 4337 19075 4403 19078
rect 7649 19075 7715 19078
rect 9121 19138 9187 19141
rect 11329 19138 11395 19141
rect 12525 19138 12591 19141
rect 9121 19136 12591 19138
rect 9121 19080 9126 19136
rect 9182 19080 11334 19136
rect 11390 19080 12530 19136
rect 12586 19080 12591 19136
rect 9121 19078 12591 19080
rect 9121 19075 9187 19078
rect 11329 19075 11395 19078
rect 12525 19075 12591 19078
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 18045 18866 18111 18869
rect 22200 18866 23000 18896
rect 18045 18864 23000 18866
rect 18045 18808 18050 18864
rect 18106 18808 23000 18864
rect 18045 18806 23000 18808
rect 18045 18803 18111 18806
rect 22200 18776 23000 18806
rect 4429 18730 4495 18733
rect 14917 18730 14983 18733
rect 15101 18730 15167 18733
rect 4429 18728 15167 18730
rect 4429 18672 4434 18728
rect 4490 18672 14922 18728
rect 14978 18672 15106 18728
rect 15162 18672 15167 18728
rect 4429 18670 15167 18672
rect 4429 18667 4495 18670
rect 14917 18667 14983 18670
rect 15101 18667 15167 18670
rect 16062 18668 16068 18732
rect 16132 18730 16138 18732
rect 18413 18730 18479 18733
rect 16132 18728 18479 18730
rect 16132 18672 18418 18728
rect 18474 18672 18479 18728
rect 16132 18670 18479 18672
rect 16132 18668 16138 18670
rect 18413 18667 18479 18670
rect 12985 18594 13051 18597
rect 14181 18594 14247 18597
rect 12985 18592 14247 18594
rect 12985 18536 12990 18592
rect 13046 18536 14186 18592
rect 14242 18536 14247 18592
rect 12985 18534 14247 18536
rect 12985 18531 13051 18534
rect 14181 18531 14247 18534
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 22200 18458 23000 18488
rect 22142 18368 23000 18458
rect 12709 18322 12775 18325
rect 17125 18322 17191 18325
rect 12709 18320 17191 18322
rect 12709 18264 12714 18320
rect 12770 18264 17130 18320
rect 17186 18264 17191 18320
rect 12709 18262 17191 18264
rect 12709 18259 12775 18262
rect 17125 18259 17191 18262
rect 17953 18322 18019 18325
rect 22142 18322 22202 18368
rect 17953 18320 22202 18322
rect 17953 18264 17958 18320
rect 18014 18264 22202 18320
rect 17953 18262 22202 18264
rect 17953 18259 18019 18262
rect 18689 18186 18755 18189
rect 18689 18184 19626 18186
rect 18689 18128 18694 18184
rect 18750 18128 19626 18184
rect 18689 18126 19626 18128
rect 18689 18123 18755 18126
rect 19566 18050 19626 18126
rect 22200 18050 23000 18080
rect 19566 17990 23000 18050
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 12157 17914 12223 17917
rect 12801 17914 12867 17917
rect 12157 17912 12867 17914
rect 12157 17856 12162 17912
rect 12218 17856 12806 17912
rect 12862 17856 12867 17912
rect 12157 17854 12867 17856
rect 12157 17851 12223 17854
rect 12801 17851 12867 17854
rect 2037 17778 2103 17781
rect 11145 17778 11211 17781
rect 2037 17776 11211 17778
rect 2037 17720 2042 17776
rect 2098 17720 11150 17776
rect 11206 17720 11211 17776
rect 2037 17718 11211 17720
rect 2037 17715 2103 17718
rect 11145 17715 11211 17718
rect 7741 17644 7807 17645
rect 7741 17642 7788 17644
rect 7696 17640 7788 17642
rect 7696 17584 7746 17640
rect 7696 17582 7788 17584
rect 7741 17580 7788 17582
rect 7852 17580 7858 17644
rect 14733 17642 14799 17645
rect 18413 17642 18479 17645
rect 22200 17642 23000 17672
rect 14733 17640 17050 17642
rect 14733 17584 14738 17640
rect 14794 17584 17050 17640
rect 14733 17582 17050 17584
rect 7741 17579 7807 17580
rect 14733 17579 14799 17582
rect 16990 17506 17050 17582
rect 18413 17640 23000 17642
rect 18413 17584 18418 17640
rect 18474 17584 23000 17640
rect 18413 17582 23000 17584
rect 18413 17579 18479 17582
rect 22200 17552 23000 17582
rect 17217 17506 17283 17509
rect 17350 17506 17356 17508
rect 16990 17504 17356 17506
rect 16990 17448 17222 17504
rect 17278 17448 17356 17504
rect 16990 17446 17356 17448
rect 17217 17443 17283 17446
rect 17350 17444 17356 17446
rect 17420 17444 17426 17508
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 9305 17234 9371 17237
rect 11237 17234 11303 17237
rect 9305 17232 11303 17234
rect 9305 17176 9310 17232
rect 9366 17176 11242 17232
rect 11298 17176 11303 17232
rect 9305 17174 11303 17176
rect 9305 17171 9371 17174
rect 11237 17171 11303 17174
rect 19241 17234 19307 17237
rect 22200 17234 23000 17264
rect 19241 17232 23000 17234
rect 19241 17176 19246 17232
rect 19302 17176 23000 17232
rect 19241 17174 23000 17176
rect 19241 17171 19307 17174
rect 22200 17144 23000 17174
rect 2773 17098 2839 17101
rect 10910 17098 10916 17100
rect 2773 17096 10916 17098
rect 2773 17040 2778 17096
rect 2834 17040 10916 17096
rect 2773 17038 10916 17040
rect 2773 17035 2839 17038
rect 10910 17036 10916 17038
rect 10980 17036 10986 17100
rect 5390 16900 5396 16964
rect 5460 16962 5466 16964
rect 5625 16962 5691 16965
rect 5460 16960 5691 16962
rect 5460 16904 5630 16960
rect 5686 16904 5691 16960
rect 5460 16902 5691 16904
rect 5460 16900 5466 16902
rect 5625 16899 5691 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 21449 16826 21515 16829
rect 22200 16826 23000 16856
rect 21449 16824 23000 16826
rect 21449 16768 21454 16824
rect 21510 16768 23000 16824
rect 21449 16766 23000 16768
rect 21449 16763 21515 16766
rect 22200 16736 23000 16766
rect 1945 16690 2011 16693
rect 9438 16690 9444 16692
rect 1945 16688 9444 16690
rect 1945 16632 1950 16688
rect 2006 16632 9444 16688
rect 1945 16630 9444 16632
rect 1945 16627 2011 16630
rect 9438 16628 9444 16630
rect 9508 16628 9514 16692
rect 13261 16690 13327 16693
rect 13486 16690 13492 16692
rect 13261 16688 13492 16690
rect 13261 16632 13266 16688
rect 13322 16632 13492 16688
rect 13261 16630 13492 16632
rect 13261 16627 13327 16630
rect 13486 16628 13492 16630
rect 13556 16628 13562 16692
rect 20110 16628 20116 16692
rect 20180 16690 20186 16692
rect 20529 16690 20595 16693
rect 20180 16688 20595 16690
rect 20180 16632 20534 16688
rect 20590 16632 20595 16688
rect 20180 16630 20595 16632
rect 20180 16628 20186 16630
rect 20529 16627 20595 16630
rect 9949 16554 10015 16557
rect 12014 16554 12020 16556
rect 9949 16552 12020 16554
rect 9949 16496 9954 16552
rect 10010 16496 12020 16552
rect 9949 16494 12020 16496
rect 9949 16491 10015 16494
rect 12014 16492 12020 16494
rect 12084 16492 12090 16556
rect 14774 16492 14780 16556
rect 14844 16554 14850 16556
rect 15561 16554 15627 16557
rect 14844 16552 15627 16554
rect 14844 16496 15566 16552
rect 15622 16496 15627 16552
rect 14844 16494 15627 16496
rect 14844 16492 14850 16494
rect 15561 16491 15627 16494
rect 20621 16554 20687 16557
rect 20621 16552 22202 16554
rect 20621 16496 20626 16552
rect 20682 16496 22202 16552
rect 20621 16494 22202 16496
rect 20621 16491 20687 16494
rect 22142 16448 22202 16494
rect 22142 16358 23000 16448
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 10174 15948 10180 16012
rect 10244 16010 10250 16012
rect 14641 16010 14707 16013
rect 16941 16012 17007 16013
rect 16941 16010 16988 16012
rect 10244 16008 14707 16010
rect 10244 15952 14646 16008
rect 14702 15952 14707 16008
rect 10244 15950 14707 15952
rect 16896 16008 16988 16010
rect 16896 15952 16946 16008
rect 16896 15950 16988 15952
rect 10244 15948 10250 15950
rect 14641 15947 14707 15950
rect 16941 15948 16988 15950
rect 17052 15948 17058 16012
rect 21357 16010 21423 16013
rect 22200 16010 23000 16040
rect 21357 16008 23000 16010
rect 21357 15952 21362 16008
rect 21418 15952 23000 16008
rect 21357 15950 23000 15952
rect 16941 15947 17007 15948
rect 21357 15947 21423 15950
rect 22200 15920 23000 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 15929 15740 15995 15741
rect 15878 15738 15884 15740
rect 15838 15678 15884 15738
rect 15948 15736 15995 15740
rect 15990 15680 15995 15736
rect 15878 15676 15884 15678
rect 15948 15676 15995 15680
rect 15929 15675 15995 15676
rect 20713 15602 20779 15605
rect 22200 15602 23000 15632
rect 20713 15600 23000 15602
rect 20713 15544 20718 15600
rect 20774 15544 23000 15600
rect 20713 15542 23000 15544
rect 20713 15539 20779 15542
rect 22200 15512 23000 15542
rect 5758 15404 5764 15468
rect 5828 15466 5834 15468
rect 6361 15466 6427 15469
rect 13261 15466 13327 15469
rect 5828 15464 13327 15466
rect 5828 15408 6366 15464
rect 6422 15408 13266 15464
rect 13322 15408 13327 15464
rect 5828 15406 13327 15408
rect 5828 15404 5834 15406
rect 6361 15403 6427 15406
rect 13261 15403 13327 15406
rect 4102 15268 4108 15332
rect 4172 15330 4178 15332
rect 4613 15330 4679 15333
rect 4172 15328 4679 15330
rect 4172 15272 4618 15328
rect 4674 15272 4679 15328
rect 4172 15270 4679 15272
rect 4172 15268 4178 15270
rect 4613 15267 4679 15270
rect 8518 15268 8524 15332
rect 8588 15330 8594 15332
rect 9213 15330 9279 15333
rect 8588 15328 9279 15330
rect 8588 15272 9218 15328
rect 9274 15272 9279 15328
rect 8588 15270 9279 15272
rect 8588 15268 8594 15270
rect 9213 15267 9279 15270
rect 14181 15330 14247 15333
rect 15326 15330 15332 15332
rect 14181 15328 15332 15330
rect 14181 15272 14186 15328
rect 14242 15272 15332 15328
rect 14181 15270 15332 15272
rect 14181 15267 14247 15270
rect 15326 15268 15332 15270
rect 15396 15268 15402 15332
rect 18873 15330 18939 15333
rect 19742 15330 19748 15332
rect 18873 15328 19748 15330
rect 18873 15272 18878 15328
rect 18934 15272 19748 15328
rect 18873 15270 19748 15272
rect 18873 15267 18939 15270
rect 19742 15268 19748 15270
rect 19812 15268 19818 15332
rect 19926 15268 19932 15332
rect 19996 15330 20002 15332
rect 20161 15330 20227 15333
rect 19996 15328 20227 15330
rect 19996 15272 20166 15328
rect 20222 15272 20227 15328
rect 19996 15270 20227 15272
rect 19996 15268 20002 15270
rect 20161 15267 20227 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 22200 15194 23000 15224
rect 22142 15104 23000 15194
rect 16297 15058 16363 15061
rect 18229 15058 18295 15061
rect 16297 15056 18295 15058
rect 16297 15000 16302 15056
rect 16358 15000 18234 15056
rect 18290 15000 18295 15056
rect 16297 14998 18295 15000
rect 16297 14995 16363 14998
rect 18229 14995 18295 14998
rect 21449 15058 21515 15061
rect 22142 15058 22202 15104
rect 21449 15056 22202 15058
rect 21449 15000 21454 15056
rect 21510 15000 22202 15056
rect 21449 14998 22202 15000
rect 21449 14995 21515 14998
rect 8569 14922 8635 14925
rect 19609 14922 19675 14925
rect 8569 14920 19675 14922
rect 8569 14864 8574 14920
rect 8630 14864 19614 14920
rect 19670 14864 19675 14920
rect 8569 14862 19675 14864
rect 8569 14859 8635 14862
rect 19609 14859 19675 14862
rect 14457 14786 14523 14789
rect 17677 14786 17743 14789
rect 17902 14786 17908 14788
rect 14457 14784 17908 14786
rect 14457 14728 14462 14784
rect 14518 14728 17682 14784
rect 17738 14728 17908 14784
rect 14457 14726 17908 14728
rect 14457 14723 14523 14726
rect 17677 14723 17743 14726
rect 17902 14724 17908 14726
rect 17972 14724 17978 14788
rect 19517 14786 19583 14789
rect 22200 14786 23000 14816
rect 19517 14784 23000 14786
rect 19517 14728 19522 14784
rect 19578 14728 23000 14784
rect 19517 14726 23000 14728
rect 19517 14723 19583 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 18321 14516 18387 14517
rect 18270 14514 18276 14516
rect 18230 14454 18276 14514
rect 18340 14512 18387 14516
rect 18382 14456 18387 14512
rect 18270 14452 18276 14454
rect 18340 14452 18387 14456
rect 18321 14451 18387 14452
rect 21357 14378 21423 14381
rect 22200 14378 23000 14408
rect 21357 14376 23000 14378
rect 21357 14320 21362 14376
rect 21418 14320 23000 14376
rect 21357 14318 23000 14320
rect 21357 14315 21423 14318
rect 22200 14288 23000 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 5349 13970 5415 13973
rect 11830 13970 11836 13972
rect 5349 13968 11836 13970
rect 5349 13912 5354 13968
rect 5410 13912 11836 13968
rect 5349 13910 11836 13912
rect 5349 13907 5415 13910
rect 11830 13908 11836 13910
rect 11900 13908 11906 13972
rect 12934 13908 12940 13972
rect 13004 13970 13010 13972
rect 13629 13970 13695 13973
rect 13004 13968 13695 13970
rect 13004 13912 13634 13968
rect 13690 13912 13695 13968
rect 13004 13910 13695 13912
rect 13004 13908 13010 13910
rect 13629 13907 13695 13910
rect 19241 13970 19307 13973
rect 22200 13970 23000 14000
rect 19241 13968 23000 13970
rect 19241 13912 19246 13968
rect 19302 13912 23000 13968
rect 19241 13910 23000 13912
rect 19241 13907 19307 13910
rect 22200 13880 23000 13910
rect 6545 13834 6611 13837
rect 9213 13834 9279 13837
rect 6545 13832 9279 13834
rect 6545 13776 6550 13832
rect 6606 13776 9218 13832
rect 9274 13776 9279 13832
rect 6545 13774 9279 13776
rect 6545 13771 6611 13774
rect 9213 13771 9279 13774
rect 18086 13772 18092 13836
rect 18156 13834 18162 13836
rect 18229 13834 18295 13837
rect 18156 13832 18295 13834
rect 18156 13776 18234 13832
rect 18290 13776 18295 13832
rect 18156 13774 18295 13776
rect 18156 13772 18162 13774
rect 18229 13771 18295 13774
rect 9438 13636 9444 13700
rect 9508 13698 9514 13700
rect 12617 13698 12683 13701
rect 9508 13696 12683 13698
rect 9508 13640 12622 13696
rect 12678 13640 12683 13696
rect 9508 13638 12683 13640
rect 9508 13636 9514 13638
rect 12617 13635 12683 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 21357 13562 21423 13565
rect 22200 13562 23000 13592
rect 21357 13560 23000 13562
rect 21357 13504 21362 13560
rect 21418 13504 23000 13560
rect 21357 13502 23000 13504
rect 21357 13499 21423 13502
rect 22200 13472 23000 13502
rect 16757 13426 16823 13429
rect 17166 13426 17172 13428
rect 16757 13424 17172 13426
rect 16757 13368 16762 13424
rect 16818 13368 17172 13424
rect 16757 13366 17172 13368
rect 16757 13363 16823 13366
rect 17166 13364 17172 13366
rect 17236 13426 17242 13428
rect 19793 13426 19859 13429
rect 17236 13424 19859 13426
rect 17236 13368 19798 13424
rect 19854 13368 19859 13424
rect 17236 13366 19859 13368
rect 17236 13364 17242 13366
rect 19793 13363 19859 13366
rect 11145 13290 11211 13293
rect 12157 13290 12223 13293
rect 18413 13290 18479 13293
rect 11145 13288 12450 13290
rect 11145 13232 11150 13288
rect 11206 13232 12162 13288
rect 12218 13232 12450 13288
rect 11145 13230 12450 13232
rect 11145 13227 11211 13230
rect 12157 13227 12223 13230
rect 12390 13154 12450 13230
rect 18413 13288 22202 13290
rect 18413 13232 18418 13288
rect 18474 13232 22202 13288
rect 18413 13230 22202 13232
rect 18413 13227 18479 13230
rect 22142 13184 22202 13230
rect 15510 13154 15516 13156
rect 12390 13094 15516 13154
rect 15510 13092 15516 13094
rect 15580 13092 15586 13156
rect 17718 13092 17724 13156
rect 17788 13154 17794 13156
rect 17861 13154 17927 13157
rect 17788 13152 17927 13154
rect 17788 13096 17866 13152
rect 17922 13096 17927 13152
rect 17788 13094 17927 13096
rect 22142 13094 23000 13184
rect 17788 13092 17794 13094
rect 17861 13091 17927 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 9305 12884 9371 12885
rect 9254 12882 9260 12884
rect 9214 12822 9260 12882
rect 9324 12880 9371 12884
rect 9366 12824 9371 12880
rect 9254 12820 9260 12822
rect 9324 12820 9371 12824
rect 9305 12819 9371 12820
rect 9489 12882 9555 12885
rect 12893 12882 12959 12885
rect 9489 12880 12959 12882
rect 9489 12824 9494 12880
rect 9550 12824 12898 12880
rect 12954 12824 12959 12880
rect 9489 12822 12959 12824
rect 9489 12819 9555 12822
rect 12893 12819 12959 12822
rect 3141 12746 3207 12749
rect 5717 12746 5783 12749
rect 15561 12746 15627 12749
rect 15837 12746 15903 12749
rect 3141 12744 5642 12746
rect 3141 12688 3146 12744
rect 3202 12688 5642 12744
rect 3141 12686 5642 12688
rect 3141 12683 3207 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 5582 12474 5642 12686
rect 5717 12744 14474 12746
rect 5717 12688 5722 12744
rect 5778 12688 14474 12744
rect 5717 12686 14474 12688
rect 5717 12683 5783 12686
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 5582 12414 6930 12474
rect 6870 12340 6930 12414
rect 6862 12276 6868 12340
rect 6932 12276 6938 12340
rect 9673 12338 9739 12341
rect 14181 12338 14247 12341
rect 9673 12336 14247 12338
rect 9673 12280 9678 12336
rect 9734 12280 14186 12336
rect 14242 12280 14247 12336
rect 9673 12278 14247 12280
rect 14414 12338 14474 12686
rect 15561 12744 15903 12746
rect 15561 12688 15566 12744
rect 15622 12688 15842 12744
rect 15898 12688 15903 12744
rect 15561 12686 15903 12688
rect 15561 12683 15627 12686
rect 15837 12683 15903 12686
rect 17953 12746 18019 12749
rect 22200 12746 23000 12776
rect 17953 12744 23000 12746
rect 17953 12688 17958 12744
rect 18014 12688 23000 12744
rect 17953 12686 23000 12688
rect 17953 12683 18019 12686
rect 22200 12656 23000 12686
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 17493 12338 17559 12341
rect 14414 12336 17559 12338
rect 14414 12280 17498 12336
rect 17554 12280 17559 12336
rect 14414 12278 17559 12280
rect 9673 12275 9739 12278
rect 14181 12275 14247 12278
rect 17493 12275 17559 12278
rect 17769 12338 17835 12341
rect 22200 12338 23000 12368
rect 17769 12336 23000 12338
rect 17769 12280 17774 12336
rect 17830 12280 23000 12336
rect 17769 12278 23000 12280
rect 17769 12275 17835 12278
rect 22200 12248 23000 12278
rect 11053 12202 11119 12205
rect 16849 12202 16915 12205
rect 17534 12202 17540 12204
rect 11053 12200 11162 12202
rect 11053 12144 11058 12200
rect 11114 12144 11162 12200
rect 11053 12139 11162 12144
rect 16849 12200 17540 12202
rect 16849 12144 16854 12200
rect 16910 12144 17540 12200
rect 16849 12142 17540 12144
rect 16849 12139 16915 12142
rect 17534 12140 17540 12142
rect 17604 12202 17610 12204
rect 18781 12202 18847 12205
rect 17604 12200 18847 12202
rect 17604 12144 18786 12200
rect 18842 12144 18847 12200
rect 17604 12142 18847 12144
rect 17604 12140 17610 12142
rect 18781 12139 18847 12142
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11102 11525 11162 12139
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 13353 11930 13419 11933
rect 16389 11930 16455 11933
rect 19333 11930 19399 11933
rect 22200 11930 23000 11960
rect 13353 11928 16455 11930
rect 13353 11872 13358 11928
rect 13414 11872 16394 11928
rect 16450 11872 16455 11928
rect 13353 11870 16455 11872
rect 13353 11867 13419 11870
rect 16389 11867 16455 11870
rect 16990 11928 19399 11930
rect 16990 11872 19338 11928
rect 19394 11872 19399 11928
rect 16990 11870 19399 11872
rect 12709 11794 12775 11797
rect 12985 11794 13051 11797
rect 16990 11794 17050 11870
rect 19333 11867 19399 11870
rect 22142 11840 23000 11930
rect 12709 11792 17050 11794
rect 12709 11736 12714 11792
rect 12770 11736 12990 11792
rect 13046 11736 17050 11792
rect 12709 11734 17050 11736
rect 18045 11794 18111 11797
rect 22142 11794 22202 11840
rect 18045 11792 22202 11794
rect 18045 11736 18050 11792
rect 18106 11736 22202 11792
rect 18045 11734 22202 11736
rect 12709 11731 12775 11734
rect 12985 11731 13051 11734
rect 18045 11731 18111 11734
rect 18968 11598 19626 11658
rect 18968 11525 19028 11598
rect 11053 11520 11162 11525
rect 11053 11464 11058 11520
rect 11114 11464 11162 11520
rect 11053 11462 11162 11464
rect 18965 11520 19031 11525
rect 18965 11464 18970 11520
rect 19026 11464 19031 11520
rect 11053 11459 11119 11462
rect 18965 11459 19031 11464
rect 19566 11522 19626 11598
rect 22200 11522 23000 11552
rect 19566 11462 23000 11522
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 10133 11386 10199 11389
rect 12382 11386 12388 11388
rect 10133 11384 12388 11386
rect 10133 11328 10138 11384
rect 10194 11328 12388 11384
rect 10133 11326 12388 11328
rect 10133 11323 10199 11326
rect 12382 11324 12388 11326
rect 12452 11324 12458 11388
rect 2129 11250 2195 11253
rect 11421 11250 11487 11253
rect 2129 11248 11487 11250
rect 2129 11192 2134 11248
rect 2190 11192 11426 11248
rect 11482 11192 11487 11248
rect 2129 11190 11487 11192
rect 2129 11187 2195 11190
rect 11421 11187 11487 11190
rect 11830 11188 11836 11252
rect 11900 11250 11906 11252
rect 12198 11250 12204 11252
rect 11900 11190 12204 11250
rect 11900 11188 11906 11190
rect 12198 11188 12204 11190
rect 12268 11250 12274 11252
rect 12709 11250 12775 11253
rect 12268 11248 12775 11250
rect 12268 11192 12714 11248
rect 12770 11192 12775 11248
rect 12268 11190 12775 11192
rect 12268 11188 12274 11190
rect 12709 11187 12775 11190
rect 17493 11250 17559 11253
rect 17493 11248 20178 11250
rect 17493 11192 17498 11248
rect 17554 11192 20178 11248
rect 17493 11190 20178 11192
rect 17493 11187 17559 11190
rect 5533 11116 5599 11117
rect 5533 11114 5580 11116
rect 5488 11112 5580 11114
rect 5488 11056 5538 11112
rect 5488 11054 5580 11056
rect 5533 11052 5580 11054
rect 5644 11052 5650 11116
rect 6862 11052 6868 11116
rect 6932 11114 6938 11116
rect 8017 11114 8083 11117
rect 6932 11112 8083 11114
rect 6932 11056 8022 11112
rect 8078 11056 8083 11112
rect 6932 11054 8083 11056
rect 6932 11052 6938 11054
rect 5533 11051 5599 11052
rect 8017 11051 8083 11054
rect 12617 11114 12683 11117
rect 15142 11114 15148 11116
rect 12617 11112 15148 11114
rect 12617 11056 12622 11112
rect 12678 11056 15148 11112
rect 12617 11054 15148 11056
rect 12617 11051 12683 11054
rect 15142 11052 15148 11054
rect 15212 11052 15218 11116
rect 18822 11052 18828 11116
rect 18892 11114 18898 11116
rect 19926 11114 19932 11116
rect 18892 11054 19932 11114
rect 18892 11052 18898 11054
rect 19926 11052 19932 11054
rect 19996 11052 20002 11116
rect 20118 11114 20178 11190
rect 22200 11114 23000 11144
rect 20118 11054 23000 11114
rect 22200 11024 23000 11054
rect 12893 10978 12959 10981
rect 16062 10978 16068 10980
rect 12893 10976 16068 10978
rect 12893 10920 12898 10976
rect 12954 10920 16068 10976
rect 12893 10918 16068 10920
rect 12893 10915 12959 10918
rect 16062 10916 16068 10918
rect 16132 10916 16138 10980
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 9397 10844 9463 10845
rect 9397 10842 9444 10844
rect 9352 10840 9444 10842
rect 9352 10784 9402 10840
rect 9352 10782 9444 10784
rect 9397 10780 9444 10782
rect 9508 10780 9514 10844
rect 13077 10842 13143 10845
rect 16297 10842 16363 10845
rect 13077 10840 16363 10842
rect 13077 10784 13082 10840
rect 13138 10784 16302 10840
rect 16358 10784 16363 10840
rect 13077 10782 16363 10784
rect 9397 10779 9463 10780
rect 13077 10779 13143 10782
rect 16297 10779 16363 10782
rect 17902 10780 17908 10844
rect 17972 10842 17978 10844
rect 18229 10842 18295 10845
rect 17972 10840 18295 10842
rect 17972 10784 18234 10840
rect 18290 10784 18295 10840
rect 17972 10782 18295 10784
rect 17972 10780 17978 10782
rect 18229 10779 18295 10782
rect 10726 10644 10732 10708
rect 10796 10706 10802 10708
rect 17585 10706 17651 10709
rect 10796 10704 17651 10706
rect 10796 10648 17590 10704
rect 17646 10648 17651 10704
rect 10796 10646 17651 10648
rect 10796 10644 10802 10646
rect 17585 10643 17651 10646
rect 17953 10706 18019 10709
rect 22200 10706 23000 10736
rect 17953 10704 23000 10706
rect 17953 10648 17958 10704
rect 18014 10648 23000 10704
rect 17953 10646 23000 10648
rect 17953 10643 18019 10646
rect 22200 10616 23000 10646
rect 19926 10570 19932 10572
rect 19014 10510 19932 10570
rect 12157 10434 12223 10437
rect 12750 10434 12756 10436
rect 12157 10432 12756 10434
rect 12157 10376 12162 10432
rect 12218 10376 12756 10432
rect 12157 10374 12756 10376
rect 12157 10371 12223 10374
rect 12750 10372 12756 10374
rect 12820 10372 12826 10436
rect 16389 10434 16455 10437
rect 19014 10434 19074 10510
rect 19926 10508 19932 10510
rect 19996 10570 20002 10572
rect 20069 10570 20135 10573
rect 19996 10568 20135 10570
rect 19996 10512 20074 10568
rect 20130 10512 20135 10568
rect 19996 10510 20135 10512
rect 19996 10508 20002 10510
rect 20069 10507 20135 10510
rect 16389 10432 19074 10434
rect 16389 10376 16394 10432
rect 16450 10376 19074 10432
rect 16389 10374 19074 10376
rect 16389 10371 16455 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 11789 10298 11855 10301
rect 12157 10298 12223 10301
rect 11789 10296 12223 10298
rect 11789 10240 11794 10296
rect 11850 10240 12162 10296
rect 12218 10240 12223 10296
rect 11789 10238 12223 10240
rect 11789 10235 11855 10238
rect 12157 10235 12223 10238
rect 15745 10298 15811 10301
rect 15878 10298 15884 10300
rect 15745 10296 15884 10298
rect 15745 10240 15750 10296
rect 15806 10240 15884 10296
rect 15745 10238 15884 10240
rect 15745 10235 15811 10238
rect 15878 10236 15884 10238
rect 15948 10236 15954 10300
rect 17493 10298 17559 10301
rect 18413 10298 18479 10301
rect 17493 10296 18479 10298
rect 17493 10240 17498 10296
rect 17554 10240 18418 10296
rect 18474 10240 18479 10296
rect 17493 10238 18479 10240
rect 17493 10235 17559 10238
rect 18413 10235 18479 10238
rect 22001 10298 22067 10301
rect 22200 10298 23000 10328
rect 22001 10296 23000 10298
rect 22001 10240 22006 10296
rect 22062 10240 23000 10296
rect 22001 10238 23000 10240
rect 22001 10235 22067 10238
rect 22200 10208 23000 10238
rect 8385 10162 8451 10165
rect 17125 10162 17191 10165
rect 8385 10160 17191 10162
rect 8385 10104 8390 10160
rect 8446 10104 17130 10160
rect 17186 10104 17191 10160
rect 8385 10102 17191 10104
rect 8385 10099 8451 10102
rect 17125 10099 17191 10102
rect 8518 9964 8524 10028
rect 8588 10026 8594 10028
rect 9305 10026 9371 10029
rect 8588 10024 9371 10026
rect 8588 9968 9310 10024
rect 9366 9968 9371 10024
rect 8588 9966 9371 9968
rect 8588 9964 8594 9966
rect 9305 9963 9371 9966
rect 13905 10026 13971 10029
rect 18505 10026 18571 10029
rect 13905 10024 18338 10026
rect 13905 9968 13910 10024
rect 13966 9968 18338 10024
rect 13905 9966 18338 9968
rect 13905 9963 13971 9966
rect 12157 9890 12223 9893
rect 16389 9890 16455 9893
rect 11838 9888 16455 9890
rect 11838 9832 12162 9888
rect 12218 9832 16394 9888
rect 16450 9832 16455 9888
rect 11838 9830 16455 9832
rect 18278 9890 18338 9966
rect 18505 10024 22202 10026
rect 18505 9968 18510 10024
rect 18566 9968 22202 10024
rect 18505 9966 22202 9968
rect 18505 9963 18571 9966
rect 22142 9920 22202 9966
rect 21081 9890 21147 9893
rect 18278 9888 21147 9890
rect 18278 9832 21086 9888
rect 21142 9832 21147 9888
rect 18278 9830 21147 9832
rect 22142 9830 23000 9920
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 5390 9692 5396 9756
rect 5460 9754 5466 9756
rect 10593 9754 10659 9757
rect 10726 9754 10732 9756
rect 5460 9694 5780 9754
rect 5460 9692 5466 9694
rect 5720 9485 5780 9694
rect 10593 9752 10732 9754
rect 10593 9696 10598 9752
rect 10654 9696 10732 9752
rect 10593 9694 10732 9696
rect 10593 9691 10659 9694
rect 10726 9692 10732 9694
rect 10796 9692 10802 9756
rect 10041 9618 10107 9621
rect 10174 9618 10180 9620
rect 10041 9616 10180 9618
rect 10041 9560 10046 9616
rect 10102 9560 10180 9616
rect 10041 9558 10180 9560
rect 10041 9555 10107 9558
rect 10174 9556 10180 9558
rect 10244 9556 10250 9620
rect 5717 9480 5783 9485
rect 5717 9424 5722 9480
rect 5778 9424 5783 9480
rect 5717 9419 5783 9424
rect 11697 9482 11763 9485
rect 11838 9482 11898 9830
rect 12157 9827 12223 9830
rect 16389 9827 16455 9830
rect 21081 9827 21147 9830
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 13486 9692 13492 9756
rect 13556 9754 13562 9756
rect 13629 9754 13695 9757
rect 20805 9754 20871 9757
rect 13556 9752 13695 9754
rect 13556 9696 13634 9752
rect 13690 9696 13695 9752
rect 13556 9694 13695 9696
rect 13556 9692 13562 9694
rect 13629 9691 13695 9694
rect 14414 9694 15026 9754
rect 12249 9618 12315 9621
rect 12566 9618 12572 9620
rect 12249 9616 12572 9618
rect 12249 9560 12254 9616
rect 12310 9560 12572 9616
rect 12249 9558 12572 9560
rect 12249 9555 12315 9558
rect 12566 9556 12572 9558
rect 12636 9618 12642 9620
rect 14414 9618 14474 9694
rect 12636 9558 14474 9618
rect 14641 9618 14707 9621
rect 14774 9618 14780 9620
rect 14641 9616 14780 9618
rect 14641 9560 14646 9616
rect 14702 9560 14780 9616
rect 14641 9558 14780 9560
rect 12636 9556 12642 9558
rect 14641 9555 14707 9558
rect 14774 9556 14780 9558
rect 14844 9556 14850 9620
rect 14966 9618 15026 9694
rect 16990 9752 20871 9754
rect 16990 9696 20810 9752
rect 20866 9696 20871 9752
rect 16990 9694 20871 9696
rect 15101 9618 15167 9621
rect 16990 9618 17050 9694
rect 20805 9691 20871 9694
rect 17585 9618 17651 9621
rect 14966 9616 17050 9618
rect 14966 9560 15106 9616
rect 15162 9560 17050 9616
rect 14966 9558 17050 9560
rect 17174 9616 17651 9618
rect 17174 9560 17590 9616
rect 17646 9560 17651 9616
rect 17174 9558 17651 9560
rect 15101 9555 15167 9558
rect 11697 9480 11898 9482
rect 11697 9424 11702 9480
rect 11758 9424 11898 9480
rect 11697 9422 11898 9424
rect 11697 9419 11763 9422
rect 12014 9420 12020 9484
rect 12084 9482 12090 9484
rect 12157 9482 12223 9485
rect 12084 9480 12223 9482
rect 12084 9424 12162 9480
rect 12218 9424 12223 9480
rect 12084 9422 12223 9424
rect 12084 9420 12090 9422
rect 12157 9419 12223 9422
rect 12709 9482 12775 9485
rect 16573 9482 16639 9485
rect 17174 9482 17234 9558
rect 17585 9555 17651 9558
rect 18689 9618 18755 9621
rect 22001 9618 22067 9621
rect 18689 9616 22067 9618
rect 18689 9560 18694 9616
rect 18750 9560 22006 9616
rect 22062 9560 22067 9616
rect 18689 9558 22067 9560
rect 18689 9555 18755 9558
rect 22001 9555 22067 9558
rect 19241 9482 19307 9485
rect 12709 9480 16452 9482
rect 12709 9424 12714 9480
rect 12770 9424 16452 9480
rect 12709 9422 16452 9424
rect 12709 9419 12775 9422
rect 16113 9346 16179 9349
rect 16246 9346 16252 9348
rect 16113 9344 16252 9346
rect 16113 9288 16118 9344
rect 16174 9288 16252 9344
rect 16113 9286 16252 9288
rect 16113 9283 16179 9286
rect 16246 9284 16252 9286
rect 16316 9284 16322 9348
rect 16392 9346 16452 9422
rect 16573 9480 17234 9482
rect 16573 9424 16578 9480
rect 16634 9424 17234 9480
rect 17864 9480 19307 9482
rect 17864 9448 19246 9480
rect 16573 9422 17234 9424
rect 17542 9424 19246 9448
rect 19302 9424 19307 9480
rect 17542 9422 19307 9424
rect 16573 9419 16639 9422
rect 17542 9388 17924 9422
rect 19241 9419 19307 9422
rect 19977 9482 20043 9485
rect 22200 9482 23000 9512
rect 19977 9480 23000 9482
rect 19977 9424 19982 9480
rect 20038 9424 23000 9480
rect 19977 9422 23000 9424
rect 19977 9419 20043 9422
rect 22200 9392 23000 9422
rect 17542 9346 17602 9388
rect 16392 9286 17602 9346
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 5349 9210 5415 9213
rect 7925 9210 7991 9213
rect 5349 9208 7991 9210
rect 5349 9152 5354 9208
rect 5410 9152 7930 9208
rect 7986 9152 7991 9208
rect 5349 9150 7991 9152
rect 5349 9147 5415 9150
rect 7925 9147 7991 9150
rect 15694 9148 15700 9212
rect 15764 9210 15770 9212
rect 16573 9210 16639 9213
rect 15764 9208 16639 9210
rect 15764 9152 16578 9208
rect 16634 9152 16639 9208
rect 15764 9150 16639 9152
rect 15764 9148 15770 9150
rect 16573 9147 16639 9150
rect 16941 9210 17007 9213
rect 17350 9210 17356 9212
rect 16941 9208 17356 9210
rect 16941 9152 16946 9208
rect 17002 9152 17356 9208
rect 16941 9150 17356 9152
rect 16941 9147 17007 9150
rect 17350 9148 17356 9150
rect 17420 9210 17426 9212
rect 17493 9210 17559 9213
rect 17420 9208 17559 9210
rect 17420 9152 17498 9208
rect 17554 9152 17559 9208
rect 17420 9150 17559 9152
rect 17420 9148 17426 9150
rect 17493 9147 17559 9150
rect 17718 9148 17724 9212
rect 17788 9210 17794 9212
rect 18229 9210 18295 9213
rect 17788 9208 18295 9210
rect 17788 9152 18234 9208
rect 18290 9152 18295 9208
rect 17788 9150 18295 9152
rect 17788 9148 17794 9150
rect 18229 9147 18295 9150
rect 8017 9074 8083 9077
rect 21357 9074 21423 9077
rect 22200 9074 23000 9104
rect 8017 9072 23000 9074
rect 8017 9016 8022 9072
rect 8078 9016 21362 9072
rect 21418 9016 23000 9072
rect 8017 9014 23000 9016
rect 8017 9011 8083 9014
rect 21357 9011 21423 9014
rect 22200 8984 23000 9014
rect 12249 8940 12315 8941
rect 12198 8938 12204 8940
rect 12158 8878 12204 8938
rect 12268 8936 12315 8940
rect 12310 8880 12315 8936
rect 12198 8876 12204 8878
rect 12268 8876 12315 8880
rect 12249 8875 12315 8876
rect 13445 8938 13511 8941
rect 17953 8938 18019 8941
rect 18086 8938 18092 8940
rect 13445 8936 18092 8938
rect 13445 8880 13450 8936
rect 13506 8880 17958 8936
rect 18014 8880 18092 8936
rect 13445 8878 18092 8880
rect 13445 8875 13511 8878
rect 17953 8875 18019 8878
rect 18086 8876 18092 8878
rect 18156 8876 18162 8940
rect 17769 8802 17835 8805
rect 18781 8802 18847 8805
rect 17769 8800 18847 8802
rect 17769 8744 17774 8800
rect 17830 8744 18786 8800
rect 18842 8744 18847 8800
rect 17769 8742 18847 8744
rect 17769 8739 17835 8742
rect 18781 8739 18847 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 7414 8604 7420 8668
rect 7484 8666 7490 8668
rect 11053 8666 11119 8669
rect 16113 8668 16179 8669
rect 7484 8664 11119 8666
rect 7484 8608 11058 8664
rect 11114 8608 11119 8664
rect 7484 8606 11119 8608
rect 7484 8604 7490 8606
rect 11053 8603 11119 8606
rect 16062 8604 16068 8668
rect 16132 8666 16179 8668
rect 17585 8666 17651 8669
rect 19057 8666 19123 8669
rect 22200 8666 23000 8696
rect 16132 8664 16224 8666
rect 16174 8608 16224 8664
rect 16132 8606 16224 8608
rect 17585 8664 19123 8666
rect 17585 8608 17590 8664
rect 17646 8608 19062 8664
rect 19118 8608 19123 8664
rect 17585 8606 19123 8608
rect 16132 8604 16179 8606
rect 16113 8603 16179 8604
rect 17585 8603 17651 8606
rect 19057 8603 19123 8606
rect 22142 8576 23000 8666
rect 7281 8530 7347 8533
rect 8201 8530 8267 8533
rect 7281 8528 8267 8530
rect 7281 8472 7286 8528
rect 7342 8472 8206 8528
rect 8262 8472 8267 8528
rect 7281 8470 8267 8472
rect 7281 8467 7347 8470
rect 8201 8467 8267 8470
rect 8334 8468 8340 8532
rect 8404 8530 8410 8532
rect 20805 8530 20871 8533
rect 22142 8530 22202 8576
rect 8404 8528 22202 8530
rect 8404 8472 20810 8528
rect 20866 8472 22202 8528
rect 8404 8470 22202 8472
rect 8404 8468 8410 8470
rect 20805 8467 20871 8470
rect 6821 8394 6887 8397
rect 7782 8394 7788 8396
rect 6821 8392 7788 8394
rect 6821 8336 6826 8392
rect 6882 8336 7788 8392
rect 6821 8334 7788 8336
rect 6821 8331 6887 8334
rect 7782 8332 7788 8334
rect 7852 8332 7858 8396
rect 8518 8332 8524 8396
rect 8588 8394 8594 8396
rect 11973 8394 12039 8397
rect 8588 8392 12039 8394
rect 8588 8336 11978 8392
rect 12034 8336 12039 8392
rect 8588 8334 12039 8336
rect 8588 8332 8594 8334
rect 11973 8331 12039 8334
rect 15142 8332 15148 8396
rect 15212 8394 15218 8396
rect 18137 8394 18203 8397
rect 15212 8392 18203 8394
rect 15212 8336 18142 8392
rect 18198 8336 18203 8392
rect 15212 8334 18203 8336
rect 15212 8332 15218 8334
rect 18137 8331 18203 8334
rect 19742 8332 19748 8396
rect 19812 8394 19818 8396
rect 19885 8394 19951 8397
rect 19812 8392 19951 8394
rect 19812 8336 19890 8392
rect 19946 8336 19951 8392
rect 19812 8334 19951 8336
rect 19812 8332 19818 8334
rect 19885 8331 19951 8334
rect 15653 8258 15719 8261
rect 18229 8258 18295 8261
rect 15653 8256 18295 8258
rect 15653 8200 15658 8256
rect 15714 8200 18234 8256
rect 18290 8200 18295 8256
rect 15653 8198 18295 8200
rect 15653 8195 15719 8198
rect 18229 8195 18295 8198
rect 19977 8258 20043 8261
rect 22200 8258 23000 8288
rect 19977 8256 23000 8258
rect 19977 8200 19982 8256
rect 20038 8200 23000 8256
rect 19977 8198 23000 8200
rect 19977 8195 20043 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 22200 8168 23000 8198
rect 19139 8127 19455 8128
rect 15193 8124 15259 8125
rect 15142 8122 15148 8124
rect 15102 8062 15148 8122
rect 15212 8120 15259 8124
rect 15254 8064 15259 8120
rect 15142 8060 15148 8062
rect 15212 8060 15259 8064
rect 15193 8059 15259 8060
rect 15561 8122 15627 8125
rect 18638 8122 18644 8124
rect 15561 8120 18644 8122
rect 15561 8064 15566 8120
rect 15622 8064 18644 8120
rect 15561 8062 18644 8064
rect 15561 8059 15627 8062
rect 18638 8060 18644 8062
rect 18708 8060 18714 8124
rect 13077 7986 13143 7989
rect 18505 7986 18571 7989
rect 13077 7984 18571 7986
rect 13077 7928 13082 7984
rect 13138 7928 18510 7984
rect 18566 7928 18571 7984
rect 13077 7926 18571 7928
rect 13077 7923 13143 7926
rect 18505 7923 18571 7926
rect 18689 7986 18755 7989
rect 18822 7986 18828 7988
rect 18689 7984 18828 7986
rect 18689 7928 18694 7984
rect 18750 7928 18828 7984
rect 18689 7926 18828 7928
rect 18689 7923 18755 7926
rect 18822 7924 18828 7926
rect 18892 7924 18898 7988
rect 8201 7850 8267 7853
rect 13721 7850 13787 7853
rect 8201 7848 13787 7850
rect 8201 7792 8206 7848
rect 8262 7792 13726 7848
rect 13782 7792 13787 7848
rect 8201 7790 13787 7792
rect 8201 7787 8267 7790
rect 13721 7787 13787 7790
rect 15193 7850 15259 7853
rect 16982 7850 16988 7852
rect 15193 7848 16988 7850
rect 15193 7792 15198 7848
rect 15254 7792 16988 7848
rect 15193 7790 16988 7792
rect 15193 7787 15259 7790
rect 16982 7788 16988 7790
rect 17052 7788 17058 7852
rect 17217 7850 17283 7853
rect 17902 7850 17908 7852
rect 17217 7848 17908 7850
rect 17217 7792 17222 7848
rect 17278 7792 17908 7848
rect 17217 7790 17908 7792
rect 17217 7787 17283 7790
rect 17902 7788 17908 7790
rect 17972 7788 17978 7852
rect 18413 7850 18479 7853
rect 20253 7850 20319 7853
rect 22200 7850 23000 7880
rect 18413 7848 23000 7850
rect 18413 7792 18418 7848
rect 18474 7792 20258 7848
rect 20314 7792 23000 7848
rect 18413 7790 23000 7792
rect 18413 7787 18479 7790
rect 20253 7787 20319 7790
rect 22200 7760 23000 7790
rect 12566 7652 12572 7716
rect 12636 7714 12642 7716
rect 13629 7714 13695 7717
rect 12636 7712 13695 7714
rect 12636 7656 13634 7712
rect 13690 7656 13695 7712
rect 12636 7654 13695 7656
rect 12636 7652 12642 7654
rect 13629 7651 13695 7654
rect 16941 7714 17007 7717
rect 17718 7714 17724 7716
rect 16941 7712 17724 7714
rect 16941 7656 16946 7712
rect 17002 7656 17724 7712
rect 16941 7654 17724 7656
rect 16941 7651 17007 7654
rect 17718 7652 17724 7654
rect 17788 7652 17794 7716
rect 18045 7714 18111 7717
rect 18270 7714 18276 7716
rect 18045 7712 18276 7714
rect 18045 7656 18050 7712
rect 18106 7656 18276 7712
rect 18045 7654 18276 7656
rect 18045 7651 18111 7654
rect 18270 7652 18276 7654
rect 18340 7652 18346 7716
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 12617 7578 12683 7581
rect 15694 7578 15700 7580
rect 12617 7576 15700 7578
rect 12617 7520 12622 7576
rect 12678 7520 15700 7576
rect 12617 7518 15700 7520
rect 12617 7515 12683 7518
rect 15694 7516 15700 7518
rect 15764 7516 15770 7580
rect 17726 7518 19626 7578
rect 8569 7442 8635 7445
rect 17726 7442 17786 7518
rect 8569 7440 17786 7442
rect 8569 7384 8574 7440
rect 8630 7384 17786 7440
rect 8569 7382 17786 7384
rect 8569 7379 8635 7382
rect 17902 7380 17908 7444
rect 17972 7442 17978 7444
rect 19333 7442 19399 7445
rect 17972 7440 19399 7442
rect 17972 7384 19338 7440
rect 19394 7384 19399 7440
rect 17972 7382 19399 7384
rect 19566 7442 19626 7518
rect 20437 7442 20503 7445
rect 22200 7442 23000 7472
rect 19566 7440 23000 7442
rect 19566 7384 20442 7440
rect 20498 7384 23000 7440
rect 19566 7382 23000 7384
rect 17972 7380 17978 7382
rect 19333 7379 19399 7382
rect 20437 7379 20503 7382
rect 22200 7352 23000 7382
rect 4705 7306 4771 7309
rect 10685 7306 10751 7309
rect 4705 7304 10751 7306
rect 4705 7248 4710 7304
rect 4766 7248 10690 7304
rect 10746 7248 10751 7304
rect 4705 7246 10751 7248
rect 4705 7243 4771 7246
rect 10685 7243 10751 7246
rect 11053 7306 11119 7309
rect 13077 7306 13143 7309
rect 11053 7304 13143 7306
rect 11053 7248 11058 7304
rect 11114 7248 13082 7304
rect 13138 7248 13143 7304
rect 11053 7246 13143 7248
rect 11053 7243 11119 7246
rect 13077 7243 13143 7246
rect 13721 7306 13787 7309
rect 19517 7306 19583 7309
rect 13721 7304 19583 7306
rect 13721 7248 13726 7304
rect 13782 7248 19522 7304
rect 19578 7248 19583 7304
rect 13721 7246 19583 7248
rect 13721 7243 13787 7246
rect 19517 7243 19583 7246
rect 10409 7170 10475 7173
rect 13813 7170 13879 7173
rect 10409 7168 13879 7170
rect 10409 7112 10414 7168
rect 10470 7112 13818 7168
rect 13874 7112 13879 7168
rect 10409 7110 13879 7112
rect 10409 7107 10475 7110
rect 13813 7107 13879 7110
rect 14365 7170 14431 7173
rect 18270 7170 18276 7172
rect 14365 7168 18276 7170
rect 14365 7112 14370 7168
rect 14426 7112 18276 7168
rect 14365 7110 18276 7112
rect 14365 7107 14431 7110
rect 18270 7108 18276 7110
rect 18340 7108 18346 7172
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 10501 7034 10567 7037
rect 12525 7034 12591 7037
rect 15653 7034 15719 7037
rect 10501 7032 12591 7034
rect 10501 6976 10506 7032
rect 10562 6976 12530 7032
rect 12586 6976 12591 7032
rect 10501 6974 12591 6976
rect 10501 6971 10567 6974
rect 12525 6971 12591 6974
rect 12758 6974 13554 7034
rect 7833 6898 7899 6901
rect 8334 6898 8340 6900
rect 7833 6896 8340 6898
rect 7833 6840 7838 6896
rect 7894 6840 8340 6896
rect 7833 6838 8340 6840
rect 7833 6835 7899 6838
rect 8334 6836 8340 6838
rect 8404 6836 8410 6900
rect 8477 6898 8543 6901
rect 12758 6898 12818 6974
rect 8477 6896 12818 6898
rect 8477 6840 8482 6896
rect 8538 6840 12818 6896
rect 8477 6838 12818 6840
rect 8477 6835 8543 6838
rect 12934 6836 12940 6900
rect 13004 6898 13010 6900
rect 13261 6898 13327 6901
rect 13004 6896 13327 6898
rect 13004 6840 13266 6896
rect 13322 6840 13327 6896
rect 13004 6838 13327 6840
rect 13494 6898 13554 6974
rect 14966 7032 15719 7034
rect 14966 6976 15658 7032
rect 15714 6976 15719 7032
rect 14966 6974 15719 6976
rect 14966 6898 15026 6974
rect 15653 6971 15719 6974
rect 19517 7034 19583 7037
rect 22200 7034 23000 7064
rect 19517 7032 23000 7034
rect 19517 6976 19522 7032
rect 19578 6976 23000 7032
rect 19517 6974 23000 6976
rect 19517 6971 19583 6974
rect 22200 6944 23000 6974
rect 13494 6838 15026 6898
rect 15193 6898 15259 6901
rect 15510 6898 15516 6900
rect 15193 6896 15516 6898
rect 15193 6840 15198 6896
rect 15254 6840 15516 6896
rect 15193 6838 15516 6840
rect 13004 6836 13010 6838
rect 13261 6835 13327 6838
rect 15193 6835 15259 6838
rect 15510 6836 15516 6838
rect 15580 6836 15586 6900
rect 16246 6836 16252 6900
rect 16316 6898 16322 6900
rect 17217 6898 17283 6901
rect 16316 6896 17283 6898
rect 16316 6840 17222 6896
rect 17278 6840 17283 6896
rect 16316 6838 17283 6840
rect 16316 6836 16322 6838
rect 17217 6835 17283 6838
rect 17401 6898 17467 6901
rect 17534 6898 17540 6900
rect 17401 6896 17540 6898
rect 17401 6840 17406 6896
rect 17462 6840 17540 6896
rect 17401 6838 17540 6840
rect 17401 6835 17467 6838
rect 17534 6836 17540 6838
rect 17604 6836 17610 6900
rect 5993 6762 6059 6765
rect 8661 6762 8727 6765
rect 5993 6760 8727 6762
rect 5993 6704 5998 6760
rect 6054 6704 8666 6760
rect 8722 6704 8727 6760
rect 5993 6702 8727 6704
rect 5993 6699 6059 6702
rect 8661 6699 8727 6702
rect 9121 6762 9187 6765
rect 18965 6762 19031 6765
rect 9121 6760 19031 6762
rect 9121 6704 9126 6760
rect 9182 6704 18970 6760
rect 19026 6704 19031 6760
rect 9121 6702 19031 6704
rect 9121 6699 9187 6702
rect 18965 6699 19031 6702
rect 19977 6762 20043 6765
rect 20110 6762 20116 6764
rect 19977 6760 20116 6762
rect 19977 6704 19982 6760
rect 20038 6704 20116 6760
rect 19977 6702 20116 6704
rect 19977 6699 20043 6702
rect 20110 6700 20116 6702
rect 20180 6700 20186 6764
rect 21590 6702 22202 6762
rect 12750 6564 12756 6628
rect 12820 6626 12826 6628
rect 15561 6626 15627 6629
rect 12820 6624 15627 6626
rect 12820 6568 15566 6624
rect 15622 6568 15627 6624
rect 12820 6566 15627 6568
rect 12820 6564 12826 6566
rect 15561 6563 15627 6566
rect 19241 6626 19307 6629
rect 21590 6626 21650 6702
rect 19241 6624 21650 6626
rect 19241 6568 19246 6624
rect 19302 6568 21650 6624
rect 19241 6566 21650 6568
rect 22142 6656 22202 6702
rect 22142 6566 23000 6656
rect 19241 6563 19307 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 8661 6490 8727 6493
rect 11973 6490 12039 6493
rect 15377 6490 15443 6493
rect 8661 6488 9506 6490
rect 8661 6432 8666 6488
rect 8722 6432 9506 6488
rect 8661 6430 9506 6432
rect 8661 6427 8727 6430
rect 9254 6354 9260 6356
rect 2730 6294 9260 6354
rect 1577 6218 1643 6221
rect 2730 6218 2790 6294
rect 9254 6292 9260 6294
rect 9324 6292 9330 6356
rect 9446 6354 9506 6430
rect 11973 6488 15443 6490
rect 11973 6432 11978 6488
rect 12034 6432 15382 6488
rect 15438 6432 15443 6488
rect 11973 6430 15443 6432
rect 11973 6427 12039 6430
rect 15377 6427 15443 6430
rect 16113 6354 16179 6357
rect 9446 6352 16179 6354
rect 9446 6296 16118 6352
rect 16174 6296 16179 6352
rect 9446 6294 16179 6296
rect 16113 6291 16179 6294
rect 16757 6354 16823 6357
rect 18229 6354 18295 6357
rect 16757 6352 18295 6354
rect 16757 6296 16762 6352
rect 16818 6296 18234 6352
rect 18290 6296 18295 6352
rect 16757 6294 18295 6296
rect 16757 6291 16823 6294
rect 18229 6291 18295 6294
rect 1577 6216 2790 6218
rect 1577 6160 1582 6216
rect 1638 6160 2790 6216
rect 1577 6158 2790 6160
rect 7465 6218 7531 6221
rect 11697 6218 11763 6221
rect 17902 6218 17908 6220
rect 7465 6216 11763 6218
rect 7465 6160 7470 6216
rect 7526 6160 11702 6216
rect 11758 6160 11763 6216
rect 7465 6158 11763 6160
rect 1577 6155 1643 6158
rect 7465 6155 7531 6158
rect 11697 6155 11763 6158
rect 13310 6158 17908 6218
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 12566 5946 12572 5948
rect 9262 5886 12572 5946
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 8017 5810 8083 5813
rect 9262 5810 9322 5886
rect 12566 5884 12572 5886
rect 12636 5884 12642 5948
rect 8017 5808 9322 5810
rect 8017 5752 8022 5808
rect 8078 5752 9322 5808
rect 8017 5750 9322 5752
rect 10501 5810 10567 5813
rect 13310 5810 13370 6158
rect 17902 6156 17908 6158
rect 17972 6156 17978 6220
rect 18965 6218 19031 6221
rect 22200 6218 23000 6248
rect 18965 6216 23000 6218
rect 18965 6160 18970 6216
rect 19026 6160 23000 6216
rect 18965 6158 23000 6160
rect 18965 6155 19031 6158
rect 22200 6128 23000 6158
rect 15377 6082 15443 6085
rect 18505 6082 18571 6085
rect 15377 6080 18571 6082
rect 15377 6024 15382 6080
rect 15438 6024 18510 6080
rect 18566 6024 18571 6080
rect 15377 6022 18571 6024
rect 15377 6019 15443 6022
rect 18505 6019 18571 6022
rect 18638 6020 18644 6084
rect 18708 6082 18714 6084
rect 18965 6082 19031 6085
rect 18708 6080 19031 6082
rect 18708 6024 18970 6080
rect 19026 6024 19031 6080
rect 18708 6022 19031 6024
rect 18708 6020 18714 6022
rect 18965 6019 19031 6022
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 15101 5948 15167 5949
rect 15101 5946 15148 5948
rect 15056 5944 15148 5946
rect 15212 5946 15218 5948
rect 16757 5946 16823 5949
rect 15212 5944 16823 5946
rect 15056 5888 15106 5944
rect 15212 5888 16762 5944
rect 16818 5888 16823 5944
rect 15056 5886 15148 5888
rect 15101 5884 15148 5886
rect 15212 5886 16823 5888
rect 15212 5884 15218 5886
rect 15101 5883 15167 5884
rect 16757 5883 16823 5886
rect 17166 5884 17172 5948
rect 17236 5946 17242 5948
rect 17677 5946 17743 5949
rect 17236 5944 17743 5946
rect 17236 5888 17682 5944
rect 17738 5888 17743 5944
rect 17236 5886 17743 5888
rect 17236 5884 17242 5886
rect 17677 5883 17743 5886
rect 10501 5808 13370 5810
rect 10501 5752 10506 5808
rect 10562 5752 13370 5808
rect 10501 5750 13370 5752
rect 13537 5810 13603 5813
rect 18229 5810 18295 5813
rect 13537 5808 18295 5810
rect 13537 5752 13542 5808
rect 13598 5752 18234 5808
rect 18290 5752 18295 5808
rect 13537 5750 18295 5752
rect 8017 5747 8083 5750
rect 10501 5747 10567 5750
rect 13537 5747 13603 5750
rect 18229 5747 18295 5750
rect 18413 5810 18479 5813
rect 22200 5810 23000 5840
rect 18413 5808 23000 5810
rect 18413 5752 18418 5808
rect 18474 5752 23000 5808
rect 18413 5750 23000 5752
rect 18413 5747 18479 5750
rect 22200 5720 23000 5750
rect 7281 5674 7347 5677
rect 12433 5674 12499 5677
rect 7281 5672 12499 5674
rect 7281 5616 7286 5672
rect 7342 5616 12438 5672
rect 12494 5616 12499 5672
rect 7281 5614 12499 5616
rect 7281 5611 7347 5614
rect 12433 5611 12499 5614
rect 12617 5674 12683 5677
rect 14273 5674 14339 5677
rect 12617 5672 14339 5674
rect 12617 5616 12622 5672
rect 12678 5616 14278 5672
rect 14334 5616 14339 5672
rect 12617 5614 14339 5616
rect 12617 5611 12683 5614
rect 14273 5611 14339 5614
rect 15193 5674 15259 5677
rect 15326 5674 15332 5676
rect 15193 5672 15332 5674
rect 15193 5616 15198 5672
rect 15254 5616 15332 5672
rect 15193 5614 15332 5616
rect 15193 5611 15259 5614
rect 15326 5612 15332 5614
rect 15396 5612 15402 5676
rect 15561 5674 15627 5677
rect 18597 5674 18663 5677
rect 15561 5672 18663 5674
rect 15561 5616 15566 5672
rect 15622 5616 18602 5672
rect 18658 5616 18663 5672
rect 15561 5614 18663 5616
rect 15561 5611 15627 5614
rect 18597 5611 18663 5614
rect 8201 5538 8267 5541
rect 10225 5538 10291 5541
rect 13077 5538 13143 5541
rect 14549 5538 14615 5541
rect 21081 5538 21147 5541
rect 8201 5536 11208 5538
rect 8201 5480 8206 5536
rect 8262 5480 10230 5536
rect 10286 5480 11208 5536
rect 8201 5478 11208 5480
rect 8201 5475 8267 5478
rect 10225 5475 10291 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11148 5266 11208 5478
rect 13077 5536 14615 5538
rect 13077 5480 13082 5536
rect 13138 5480 14554 5536
rect 14610 5480 14615 5536
rect 13077 5478 14615 5480
rect 13077 5475 13143 5478
rect 14549 5475 14615 5478
rect 17542 5536 21147 5538
rect 17542 5480 21086 5536
rect 21142 5480 21147 5536
rect 17542 5478 21147 5480
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 15929 5402 15995 5405
rect 13310 5400 15995 5402
rect 13310 5344 15934 5400
rect 15990 5344 15995 5400
rect 13310 5342 15995 5344
rect 13310 5266 13370 5342
rect 15929 5339 15995 5342
rect 15009 5266 15075 5269
rect 11148 5206 13370 5266
rect 13494 5264 15075 5266
rect 13494 5208 15014 5264
rect 15070 5208 15075 5264
rect 13494 5206 15075 5208
rect 8385 5130 8451 5133
rect 13494 5130 13554 5206
rect 15009 5203 15075 5206
rect 16021 5266 16087 5269
rect 17542 5266 17602 5478
rect 21081 5475 21147 5478
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 19057 5402 19123 5405
rect 19609 5402 19675 5405
rect 19977 5404 20043 5405
rect 19057 5400 19675 5402
rect 19057 5344 19062 5400
rect 19118 5344 19614 5400
rect 19670 5344 19675 5400
rect 19057 5342 19675 5344
rect 19057 5339 19123 5342
rect 19609 5339 19675 5342
rect 19926 5340 19932 5404
rect 19996 5402 20043 5404
rect 22200 5402 23000 5432
rect 19996 5400 20088 5402
rect 20038 5344 20088 5400
rect 19996 5342 20088 5344
rect 19996 5340 20043 5342
rect 19977 5339 20043 5340
rect 22142 5312 23000 5402
rect 16021 5264 17602 5266
rect 16021 5208 16026 5264
rect 16082 5208 17602 5264
rect 16021 5206 17602 5208
rect 17953 5266 18019 5269
rect 22142 5266 22202 5312
rect 17953 5264 22202 5266
rect 17953 5208 17958 5264
rect 18014 5208 22202 5264
rect 17953 5206 22202 5208
rect 16021 5203 16087 5206
rect 17953 5203 18019 5206
rect 8385 5128 13554 5130
rect 8385 5072 8390 5128
rect 8446 5072 13554 5128
rect 8385 5070 13554 5072
rect 13721 5130 13787 5133
rect 15469 5130 15535 5133
rect 13721 5128 15535 5130
rect 13721 5072 13726 5128
rect 13782 5072 15474 5128
rect 15530 5072 15535 5128
rect 13721 5070 15535 5072
rect 8385 5067 8451 5070
rect 13721 5067 13787 5070
rect 15469 5067 15535 5070
rect 17401 5130 17467 5133
rect 19793 5130 19859 5133
rect 17401 5128 19859 5130
rect 17401 5072 17406 5128
rect 17462 5072 19798 5128
rect 19854 5072 19859 5128
rect 17401 5070 19859 5072
rect 17401 5067 17467 5070
rect 19793 5067 19859 5070
rect 16062 4932 16068 4996
rect 16132 4994 16138 4996
rect 17861 4994 17927 4997
rect 16132 4992 17927 4994
rect 16132 4936 17866 4992
rect 17922 4936 17927 4992
rect 16132 4934 17927 4936
rect 16132 4932 16138 4934
rect 17861 4931 17927 4934
rect 19609 4994 19675 4997
rect 22200 4994 23000 5024
rect 19609 4992 23000 4994
rect 19609 4936 19614 4992
rect 19670 4936 23000 4992
rect 19609 4934 23000 4936
rect 19609 4931 19675 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 9213 4858 9279 4861
rect 9213 4856 12450 4858
rect 9213 4800 9218 4856
rect 9274 4800 12450 4856
rect 9213 4798 12450 4800
rect 9213 4795 9279 4798
rect 10726 4660 10732 4724
rect 10796 4722 10802 4724
rect 11973 4722 12039 4725
rect 10796 4720 12039 4722
rect 10796 4664 11978 4720
rect 12034 4664 12039 4720
rect 10796 4662 12039 4664
rect 12390 4722 12450 4798
rect 13813 4722 13879 4725
rect 12390 4720 13879 4722
rect 12390 4664 13818 4720
rect 13874 4664 13879 4720
rect 12390 4662 13879 4664
rect 10796 4660 10802 4662
rect 11973 4659 12039 4662
rect 13813 4659 13879 4662
rect 15101 4722 15167 4725
rect 19149 4722 19215 4725
rect 15101 4720 19215 4722
rect 15101 4664 15106 4720
rect 15162 4664 19154 4720
rect 19210 4664 19215 4720
rect 15101 4662 19215 4664
rect 15101 4659 15167 4662
rect 19149 4659 19215 4662
rect 9305 4586 9371 4589
rect 19241 4586 19307 4589
rect 22200 4586 23000 4616
rect 9305 4584 23000 4586
rect 9305 4528 9310 4584
rect 9366 4528 19246 4584
rect 19302 4528 23000 4584
rect 9305 4526 23000 4528
rect 9305 4523 9371 4526
rect 19241 4523 19307 4526
rect 22200 4496 23000 4526
rect 17861 4450 17927 4453
rect 20621 4450 20687 4453
rect 17861 4448 20687 4450
rect 17861 4392 17866 4448
rect 17922 4392 20626 4448
rect 20682 4392 20687 4448
rect 17861 4390 20687 4392
rect 17861 4387 17927 4390
rect 20621 4387 20687 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 10961 4316 11027 4317
rect 10910 4252 10916 4316
rect 10980 4314 11027 4316
rect 15653 4316 15719 4317
rect 15653 4314 15700 4316
rect 10980 4312 11072 4314
rect 11022 4256 11072 4312
rect 10980 4254 11072 4256
rect 15608 4312 15700 4314
rect 15608 4256 15658 4312
rect 15608 4254 15700 4256
rect 10980 4252 11027 4254
rect 10961 4251 11027 4252
rect 15653 4252 15700 4254
rect 15764 4252 15770 4316
rect 15653 4251 15719 4252
rect 5073 4178 5139 4181
rect 8518 4178 8524 4180
rect 5073 4176 8524 4178
rect 5073 4120 5078 4176
rect 5134 4120 8524 4176
rect 5073 4118 8524 4120
rect 5073 4115 5139 4118
rect 8518 4116 8524 4118
rect 8588 4116 8594 4180
rect 11145 4178 11211 4181
rect 17033 4178 17099 4181
rect 11145 4176 17099 4178
rect 11145 4120 11150 4176
rect 11206 4120 17038 4176
rect 17094 4120 17099 4176
rect 11145 4118 17099 4120
rect 11145 4115 11211 4118
rect 17033 4115 17099 4118
rect 20713 4178 20779 4181
rect 22200 4178 23000 4208
rect 20713 4176 23000 4178
rect 20713 4120 20718 4176
rect 20774 4120 23000 4176
rect 20713 4118 23000 4120
rect 20713 4115 20779 4118
rect 22200 4088 23000 4118
rect 7966 3980 7972 4044
rect 8036 4042 8042 4044
rect 8845 4042 8911 4045
rect 8036 4040 8911 4042
rect 8036 3984 8850 4040
rect 8906 3984 8911 4040
rect 8036 3982 8911 3984
rect 8036 3980 8042 3982
rect 8845 3979 8911 3982
rect 9857 4042 9923 4045
rect 13813 4042 13879 4045
rect 9857 4040 13879 4042
rect 9857 3984 9862 4040
rect 9918 3984 13818 4040
rect 13874 3984 13879 4040
rect 9857 3982 13879 3984
rect 9857 3979 9923 3982
rect 13813 3979 13879 3982
rect 14273 4042 14339 4045
rect 14733 4042 14799 4045
rect 17677 4042 17743 4045
rect 20529 4042 20595 4045
rect 14273 4040 17743 4042
rect 14273 3984 14278 4040
rect 14334 3984 14738 4040
rect 14794 3984 17682 4040
rect 17738 3984 17743 4040
rect 14273 3982 17743 3984
rect 14273 3979 14339 3982
rect 14733 3979 14799 3982
rect 17677 3979 17743 3982
rect 17864 4040 20595 4042
rect 17864 3984 20534 4040
rect 20590 3984 20595 4040
rect 17864 3982 20595 3984
rect 6678 3844 6684 3908
rect 6748 3906 6754 3908
rect 8569 3906 8635 3909
rect 6748 3904 8635 3906
rect 6748 3848 8574 3904
rect 8630 3848 8635 3904
rect 6748 3846 8635 3848
rect 6748 3844 6754 3846
rect 8569 3843 8635 3846
rect 14825 3906 14891 3909
rect 17864 3906 17924 3982
rect 20529 3979 20595 3982
rect 14825 3904 17924 3906
rect 14825 3848 14830 3904
rect 14886 3848 17924 3904
rect 14825 3846 17924 3848
rect 14825 3843 14891 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 15009 3770 15075 3773
rect 17401 3770 17467 3773
rect 15009 3768 17467 3770
rect 15009 3712 15014 3768
rect 15070 3712 17406 3768
rect 17462 3712 17467 3768
rect 15009 3710 17467 3712
rect 15009 3707 15075 3710
rect 17401 3707 17467 3710
rect 20529 3770 20595 3773
rect 22200 3770 23000 3800
rect 20529 3768 23000 3770
rect 20529 3712 20534 3768
rect 20590 3712 23000 3768
rect 20529 3710 23000 3712
rect 20529 3707 20595 3710
rect 22200 3680 23000 3710
rect 10501 3634 10567 3637
rect 17953 3634 18019 3637
rect 10501 3632 18019 3634
rect 10501 3576 10506 3632
rect 10562 3576 17958 3632
rect 18014 3576 18019 3632
rect 10501 3574 18019 3576
rect 10501 3571 10567 3574
rect 17953 3571 18019 3574
rect 9765 3498 9831 3501
rect 14181 3498 14247 3501
rect 9765 3496 14247 3498
rect 9765 3440 9770 3496
rect 9826 3440 14186 3496
rect 14242 3440 14247 3496
rect 9765 3438 14247 3440
rect 9765 3435 9831 3438
rect 14181 3435 14247 3438
rect 14641 3498 14707 3501
rect 15469 3498 15535 3501
rect 18045 3498 18111 3501
rect 14641 3496 18111 3498
rect 14641 3440 14646 3496
rect 14702 3440 15474 3496
rect 15530 3440 18050 3496
rect 18106 3440 18111 3496
rect 14641 3438 18111 3440
rect 14641 3435 14707 3438
rect 15469 3435 15535 3438
rect 18045 3435 18111 3438
rect 20529 3498 20595 3501
rect 20529 3496 22202 3498
rect 20529 3440 20534 3496
rect 20590 3440 22202 3496
rect 20529 3438 22202 3440
rect 20529 3435 20595 3438
rect 22142 3392 22202 3438
rect 22142 3302 23000 3392
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 5717 3228 5783 3229
rect 5717 3226 5764 3228
rect 5672 3224 5764 3226
rect 5672 3168 5722 3224
rect 5672 3166 5764 3168
rect 5717 3164 5764 3166
rect 5828 3164 5834 3228
rect 5717 3163 5783 3164
rect 8293 3090 8359 3093
rect 20529 3090 20595 3093
rect 8293 3088 20730 3090
rect 8293 3032 8298 3088
rect 8354 3032 20534 3088
rect 20590 3032 20730 3088
rect 8293 3030 20730 3032
rect 8293 3027 8359 3030
rect 20529 3027 20595 3030
rect 11145 2954 11211 2957
rect 19425 2954 19491 2957
rect 11145 2952 19491 2954
rect 11145 2896 11150 2952
rect 11206 2896 19430 2952
rect 19486 2896 19491 2952
rect 11145 2894 19491 2896
rect 20670 2954 20730 3030
rect 22200 2954 23000 2984
rect 20670 2894 23000 2954
rect 11145 2891 11211 2894
rect 19425 2891 19491 2894
rect 22200 2864 23000 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 4102 2620 4108 2684
rect 4172 2682 4178 2684
rect 5625 2682 5691 2685
rect 4172 2680 5691 2682
rect 4172 2624 5630 2680
rect 5686 2624 5691 2680
rect 4172 2622 5691 2624
rect 4172 2620 4178 2622
rect 5625 2619 5691 2622
rect 5574 2484 5580 2548
rect 5644 2546 5650 2548
rect 9305 2546 9371 2549
rect 17401 2546 17467 2549
rect 5644 2544 17467 2546
rect 5644 2488 9310 2544
rect 9366 2488 17406 2544
rect 17462 2488 17467 2544
rect 5644 2486 17467 2488
rect 5644 2484 5650 2486
rect 9305 2483 9371 2486
rect 17401 2483 17467 2486
rect 18965 2546 19031 2549
rect 20161 2546 20227 2549
rect 22200 2546 23000 2576
rect 18965 2544 23000 2546
rect 18965 2488 18970 2544
rect 19026 2488 20166 2544
rect 20222 2488 23000 2544
rect 18965 2486 23000 2488
rect 18965 2483 19031 2486
rect 20161 2483 20227 2486
rect 22200 2456 23000 2486
rect 5625 2410 5691 2413
rect 14365 2410 14431 2413
rect 5625 2408 14431 2410
rect 5625 2352 5630 2408
rect 5686 2352 14370 2408
rect 14426 2352 14431 2408
rect 5625 2350 14431 2352
rect 5625 2347 5691 2350
rect 14365 2347 14431 2350
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 22200 2138 23000 2168
rect 22142 2048 23000 2138
rect 20437 2002 20503 2005
rect 22142 2002 22202 2048
rect 20437 2000 22202 2002
rect 20437 1944 20442 2000
rect 20498 1944 22202 2000
rect 20437 1942 22202 1944
rect 20437 1939 20503 1942
rect 18873 1730 18939 1733
rect 22200 1730 23000 1760
rect 18873 1728 23000 1730
rect 18873 1672 18878 1728
rect 18934 1672 23000 1728
rect 18873 1670 23000 1672
rect 18873 1667 18939 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 7052 20224 7116 20228
rect 7052 20168 7066 20224
rect 7066 20168 7116 20224
rect 7052 20164 7116 20168
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 6684 19408 6748 19412
rect 6684 19352 6698 19408
rect 6698 19352 6748 19408
rect 6684 19348 6748 19352
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 7052 19348 7116 19412
rect 7420 19408 7484 19412
rect 7420 19352 7434 19408
rect 7434 19352 7484 19408
rect 7420 19348 7484 19352
rect 7972 19408 8036 19412
rect 7972 19352 7986 19408
rect 7986 19352 8036 19408
rect 7972 19348 8036 19352
rect 10732 19348 10796 19412
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 16068 18668 16132 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 7788 17640 7852 17644
rect 7788 17584 7802 17640
rect 7802 17584 7852 17640
rect 7788 17580 7852 17584
rect 17356 17444 17420 17508
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 10916 17036 10980 17100
rect 5396 16900 5460 16964
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 9444 16628 9508 16692
rect 13492 16628 13556 16692
rect 20116 16628 20180 16692
rect 12020 16492 12084 16556
rect 14780 16492 14844 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 10180 15948 10244 16012
rect 16988 16008 17052 16012
rect 16988 15952 17002 16008
rect 17002 15952 17052 16008
rect 16988 15948 17052 15952
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 15884 15736 15948 15740
rect 15884 15680 15934 15736
rect 15934 15680 15948 15736
rect 15884 15676 15948 15680
rect 5764 15404 5828 15468
rect 4108 15268 4172 15332
rect 8524 15268 8588 15332
rect 15332 15268 15396 15332
rect 19748 15268 19812 15332
rect 19932 15268 19996 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 17908 14724 17972 14788
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 18276 14512 18340 14516
rect 18276 14456 18326 14512
rect 18326 14456 18340 14512
rect 18276 14452 18340 14456
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 11836 13908 11900 13972
rect 12940 13908 13004 13972
rect 18092 13772 18156 13836
rect 9444 13636 9508 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 17172 13364 17236 13428
rect 15516 13092 15580 13156
rect 17724 13092 17788 13156
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 9260 12880 9324 12884
rect 9260 12824 9310 12880
rect 9310 12824 9324 12880
rect 9260 12820 9324 12824
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 6868 12276 6932 12340
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 17540 12140 17604 12204
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 12388 11324 12452 11388
rect 11836 11188 11900 11252
rect 12204 11188 12268 11252
rect 5580 11112 5644 11116
rect 5580 11056 5594 11112
rect 5594 11056 5644 11112
rect 5580 11052 5644 11056
rect 6868 11052 6932 11116
rect 15148 11052 15212 11116
rect 18828 11052 18892 11116
rect 19932 11052 19996 11116
rect 16068 10916 16132 10980
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 9444 10840 9508 10844
rect 9444 10784 9458 10840
rect 9458 10784 9508 10840
rect 9444 10780 9508 10784
rect 17908 10780 17972 10844
rect 10732 10644 10796 10708
rect 12756 10372 12820 10436
rect 19932 10508 19996 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 15884 10236 15948 10300
rect 8524 9964 8588 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 5396 9692 5460 9756
rect 10732 9692 10796 9756
rect 10180 9556 10244 9620
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 13492 9692 13556 9756
rect 12572 9556 12636 9620
rect 14780 9556 14844 9620
rect 12020 9420 12084 9484
rect 16252 9284 16316 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 15700 9148 15764 9212
rect 17356 9148 17420 9212
rect 17724 9148 17788 9212
rect 12204 8936 12268 8940
rect 12204 8880 12254 8936
rect 12254 8880 12268 8936
rect 12204 8876 12268 8880
rect 18092 8876 18156 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 7420 8604 7484 8668
rect 16068 8664 16132 8668
rect 16068 8608 16118 8664
rect 16118 8608 16132 8664
rect 16068 8604 16132 8608
rect 8340 8468 8404 8532
rect 7788 8332 7852 8396
rect 8524 8332 8588 8396
rect 15148 8332 15212 8396
rect 19748 8332 19812 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 15148 8120 15212 8124
rect 15148 8064 15198 8120
rect 15198 8064 15212 8120
rect 15148 8060 15212 8064
rect 18644 8060 18708 8124
rect 18828 7924 18892 7988
rect 16988 7788 17052 7852
rect 17908 7788 17972 7852
rect 12572 7652 12636 7716
rect 17724 7652 17788 7716
rect 18276 7652 18340 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 15700 7516 15764 7580
rect 17908 7380 17972 7444
rect 18276 7108 18340 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 8340 6836 8404 6900
rect 12940 6836 13004 6900
rect 15516 6836 15580 6900
rect 16252 6836 16316 6900
rect 17540 6836 17604 6900
rect 20116 6700 20180 6764
rect 12756 6564 12820 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 9260 6292 9324 6356
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 12572 5884 12636 5948
rect 17908 6156 17972 6220
rect 18644 6020 18708 6084
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 15148 5944 15212 5948
rect 15148 5888 15162 5944
rect 15162 5888 15212 5944
rect 15148 5884 15212 5888
rect 17172 5884 17236 5948
rect 15332 5612 15396 5676
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 19932 5400 19996 5404
rect 19932 5344 19982 5400
rect 19982 5344 19996 5400
rect 19932 5340 19996 5344
rect 16068 4932 16132 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 10732 4660 10796 4724
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 10916 4312 10980 4316
rect 10916 4256 10966 4312
rect 10966 4256 10980 4312
rect 10916 4252 10980 4256
rect 15700 4312 15764 4316
rect 15700 4256 15714 4312
rect 15714 4256 15764 4312
rect 15700 4252 15764 4256
rect 8524 4116 8588 4180
rect 7972 3980 8036 4044
rect 6684 3844 6748 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 5764 3224 5828 3228
rect 5764 3168 5778 3224
rect 5778 3168 5828 3224
rect 5764 3164 5828 3168
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 4108 2620 4172 2684
rect 5580 2484 5644 2548
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 7051 20228 7117 20229
rect 7051 20164 7052 20228
rect 7116 20164 7117 20228
rect 7051 20163 7117 20164
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 7054 19413 7114 20163
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 7051 19412 7117 19413
rect 7051 19348 7052 19412
rect 7116 19348 7117 19412
rect 7051 19347 7117 19348
rect 7419 19412 7485 19413
rect 7419 19348 7420 19412
rect 7484 19348 7485 19412
rect 7419 19347 7485 19348
rect 7971 19412 8037 19413
rect 7971 19348 7972 19412
rect 8036 19348 8037 19412
rect 7971 19347 8037 19348
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5395 16964 5461 16965
rect 5395 16900 5396 16964
rect 5460 16900 5461 16964
rect 5395 16899 5461 16900
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 4110 2685 4170 15267
rect 5398 9757 5458 16899
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 5763 15468 5829 15469
rect 5763 15404 5764 15468
rect 5828 15404 5829 15468
rect 5763 15403 5829 15404
rect 5579 11116 5645 11117
rect 5579 11052 5580 11116
rect 5644 11052 5645 11116
rect 5579 11051 5645 11052
rect 5395 9756 5461 9757
rect 5395 9692 5396 9756
rect 5460 9692 5461 9756
rect 5395 9691 5461 9692
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 5582 2549 5642 11051
rect 5766 3229 5826 15403
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6686 3909 6746 19347
rect 6867 12340 6933 12341
rect 6867 12276 6868 12340
rect 6932 12276 6933 12340
rect 6867 12275 6933 12276
rect 6870 11117 6930 12275
rect 6867 11116 6933 11117
rect 6867 11052 6868 11116
rect 6932 11052 6933 11116
rect 6867 11051 6933 11052
rect 7422 8669 7482 19347
rect 7787 17644 7853 17645
rect 7787 17580 7788 17644
rect 7852 17580 7853 17644
rect 7787 17579 7853 17580
rect 7419 8668 7485 8669
rect 7419 8604 7420 8668
rect 7484 8604 7485 8668
rect 7419 8603 7485 8604
rect 7790 8397 7850 17579
rect 7787 8396 7853 8397
rect 7787 8332 7788 8396
rect 7852 8332 7853 8396
rect 7787 8331 7853 8332
rect 7974 4045 8034 19347
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 10731 19412 10797 19413
rect 10731 19348 10732 19412
rect 10796 19348 10797 19412
rect 10731 19347 10797 19348
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 9443 16692 9509 16693
rect 9443 16628 9444 16692
rect 9508 16628 9509 16692
rect 9443 16627 9509 16628
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8523 15332 8589 15333
rect 8523 15268 8524 15332
rect 8588 15268 8589 15332
rect 8523 15267 8589 15268
rect 8526 10029 8586 15267
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 9446 13701 9506 16627
rect 10179 16012 10245 16013
rect 10179 15948 10180 16012
rect 10244 15948 10245 16012
rect 10179 15947 10245 15948
rect 9443 13700 9509 13701
rect 9443 13636 9444 13700
rect 9508 13636 9509 13700
rect 9443 13635 9509 13636
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 9259 12884 9325 12885
rect 9259 12820 9260 12884
rect 9324 12820 9325 12884
rect 9259 12819 9325 12820
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8523 10028 8589 10029
rect 8523 9964 8524 10028
rect 8588 9964 8589 10028
rect 8523 9963 8589 9964
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8339 8532 8405 8533
rect 8339 8468 8340 8532
rect 8404 8468 8405 8532
rect 8339 8467 8405 8468
rect 8342 6901 8402 8467
rect 8523 8396 8589 8397
rect 8523 8332 8524 8396
rect 8588 8332 8589 8396
rect 8523 8331 8589 8332
rect 8339 6900 8405 6901
rect 8339 6836 8340 6900
rect 8404 6836 8405 6900
rect 8339 6835 8405 6836
rect 8526 4181 8586 8331
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 9262 6357 9322 12819
rect 9446 10845 9506 13635
rect 9443 10844 9509 10845
rect 9443 10780 9444 10844
rect 9508 10780 9509 10844
rect 9443 10779 9509 10780
rect 10182 9621 10242 15947
rect 10734 10709 10794 19347
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 10915 17100 10981 17101
rect 10915 17036 10916 17100
rect 10980 17036 10981 17100
rect 10915 17035 10981 17036
rect 10731 10708 10797 10709
rect 10731 10644 10732 10708
rect 10796 10644 10797 10708
rect 10731 10643 10797 10644
rect 10731 9756 10797 9757
rect 10731 9692 10732 9756
rect 10796 9692 10797 9756
rect 10731 9691 10797 9692
rect 10179 9620 10245 9621
rect 10179 9556 10180 9620
rect 10244 9556 10245 9620
rect 10179 9555 10245 9556
rect 9259 6356 9325 6357
rect 9259 6292 9260 6356
rect 9324 6292 9325 6356
rect 9259 6291 9325 6292
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8523 4180 8589 4181
rect 8523 4116 8524 4180
rect 8588 4116 8589 4180
rect 8523 4115 8589 4116
rect 7971 4044 8037 4045
rect 7971 3980 7972 4044
rect 8036 3980 8037 4044
rect 7971 3979 8037 3980
rect 6683 3908 6749 3909
rect 6683 3844 6684 3908
rect 6748 3844 6749 3908
rect 6683 3843 6749 3844
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5763 3228 5829 3229
rect 5763 3164 5764 3228
rect 5828 3164 5829 3228
rect 5763 3163 5829 3164
rect 5579 2548 5645 2549
rect 5579 2484 5580 2548
rect 5644 2484 5645 2548
rect 5579 2483 5645 2484
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 3840 9061 4864
rect 10734 4725 10794 9691
rect 10731 4724 10797 4725
rect 10731 4660 10732 4724
rect 10796 4660 10797 4724
rect 10731 4659 10797 4660
rect 10918 4317 10978 17035
rect 11340 16352 11660 17376
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16067 18732 16133 18733
rect 16067 18668 16068 18732
rect 16132 18668 16133 18732
rect 16067 18667 16133 18668
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12019 16556 12085 16557
rect 12019 16492 12020 16556
rect 12084 16492 12085 16556
rect 12019 16491 12085 16492
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11835 13972 11901 13973
rect 11835 13908 11836 13972
rect 11900 13908 11901 13972
rect 11835 13907 11901 13908
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11838 11253 11898 13907
rect 11835 11252 11901 11253
rect 11835 11188 11836 11252
rect 11900 11188 11901 11252
rect 11835 11187 11901 11188
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 12022 9485 12082 16491
rect 12939 13972 13005 13973
rect 12939 13908 12940 13972
rect 13004 13908 13005 13972
rect 12939 13907 13005 13908
rect 12387 11388 12453 11389
rect 12387 11324 12388 11388
rect 12452 11324 12453 11388
rect 12387 11323 12453 11324
rect 12203 11252 12269 11253
rect 12203 11188 12204 11252
rect 12268 11188 12269 11252
rect 12390 11250 12450 11323
rect 12390 11190 12634 11250
rect 12203 11187 12269 11188
rect 12019 9484 12085 9485
rect 12019 9420 12020 9484
rect 12084 9420 12085 9484
rect 12019 9419 12085 9420
rect 12206 8941 12266 11187
rect 12574 9621 12634 11190
rect 12755 10436 12821 10437
rect 12755 10372 12756 10436
rect 12820 10372 12821 10436
rect 12755 10371 12821 10372
rect 12571 9620 12637 9621
rect 12571 9556 12572 9620
rect 12636 9556 12637 9620
rect 12571 9555 12637 9556
rect 12203 8940 12269 8941
rect 12203 8876 12204 8940
rect 12268 8876 12269 8940
rect 12203 8875 12269 8876
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 12571 7716 12637 7717
rect 12571 7652 12572 7716
rect 12636 7652 12637 7716
rect 12571 7651 12637 7652
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 12574 5949 12634 7651
rect 12758 6629 12818 10371
rect 12942 6901 13002 13907
rect 13494 9757 13554 16627
rect 13939 15808 14259 16832
rect 14779 16556 14845 16557
rect 14779 16492 14780 16556
rect 14844 16492 14845 16556
rect 14779 16491 14845 16492
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13491 9756 13557 9757
rect 13491 9692 13492 9756
rect 13556 9692 13557 9756
rect 13491 9691 13557 9692
rect 13939 9280 14259 10304
rect 14782 9621 14842 16491
rect 15883 15740 15949 15741
rect 15883 15676 15884 15740
rect 15948 15676 15949 15740
rect 15883 15675 15949 15676
rect 15331 15332 15397 15333
rect 15331 15268 15332 15332
rect 15396 15268 15397 15332
rect 15331 15267 15397 15268
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 14779 9620 14845 9621
rect 14779 9556 14780 9620
rect 14844 9556 14845 9620
rect 14779 9555 14845 9556
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 15150 8397 15210 11051
rect 15147 8396 15213 8397
rect 15147 8332 15148 8396
rect 15212 8332 15213 8396
rect 15147 8331 15213 8332
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 15147 8124 15213 8125
rect 15147 8060 15148 8124
rect 15212 8060 15213 8124
rect 15147 8059 15213 8060
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 12939 6900 13005 6901
rect 12939 6836 12940 6900
rect 13004 6836 13005 6900
rect 12939 6835 13005 6836
rect 12755 6628 12821 6629
rect 12755 6564 12756 6628
rect 12820 6564 12821 6628
rect 12755 6563 12821 6564
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 12571 5948 12637 5949
rect 12571 5884 12572 5948
rect 12636 5884 12637 5948
rect 12571 5883 12637 5884
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 10915 4316 10981 4317
rect 10915 4252 10916 4316
rect 10980 4252 10981 4316
rect 10915 4251 10981 4252
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 4928 14259 5952
rect 15150 5949 15210 8059
rect 15147 5948 15213 5949
rect 15147 5884 15148 5948
rect 15212 5884 15213 5948
rect 15147 5883 15213 5884
rect 15334 5677 15394 15267
rect 15515 13156 15581 13157
rect 15515 13092 15516 13156
rect 15580 13092 15581 13156
rect 15515 13091 15581 13092
rect 15518 6901 15578 13091
rect 15886 10301 15946 15675
rect 16070 10981 16130 18667
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 17355 17508 17421 17509
rect 17355 17444 17356 17508
rect 17420 17444 17421 17508
rect 17355 17443 17421 17444
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16987 16012 17053 16013
rect 16987 15948 16988 16012
rect 17052 15948 17053 16012
rect 16987 15947 17053 15948
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16067 10980 16133 10981
rect 16067 10916 16068 10980
rect 16132 10916 16133 10980
rect 16067 10915 16133 10916
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 15883 10300 15949 10301
rect 15883 10236 15884 10300
rect 15948 10236 15949 10300
rect 15883 10235 15949 10236
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16251 9348 16317 9349
rect 16251 9284 16252 9348
rect 16316 9284 16317 9348
rect 16251 9283 16317 9284
rect 15699 9212 15765 9213
rect 15699 9148 15700 9212
rect 15764 9148 15765 9212
rect 15699 9147 15765 9148
rect 15702 7581 15762 9147
rect 16067 8668 16133 8669
rect 16067 8604 16068 8668
rect 16132 8604 16133 8668
rect 16067 8603 16133 8604
rect 15699 7580 15765 7581
rect 15699 7516 15700 7580
rect 15764 7516 15765 7580
rect 15699 7515 15765 7516
rect 15515 6900 15581 6901
rect 15515 6836 15516 6900
rect 15580 6836 15581 6900
rect 15515 6835 15581 6836
rect 15331 5676 15397 5677
rect 15331 5612 15332 5676
rect 15396 5612 15397 5676
rect 15331 5611 15397 5612
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 15702 4317 15762 7515
rect 16070 4997 16130 8603
rect 16254 6901 16314 9283
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16990 7853 17050 15947
rect 17171 13428 17237 13429
rect 17171 13364 17172 13428
rect 17236 13364 17237 13428
rect 17171 13363 17237 13364
rect 16987 7852 17053 7853
rect 16987 7788 16988 7852
rect 17052 7788 17053 7852
rect 16987 7787 17053 7788
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16251 6900 16317 6901
rect 16251 6836 16252 6900
rect 16316 6836 16317 6900
rect 16251 6835 16317 6836
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 17174 5949 17234 13363
rect 17358 9213 17418 17443
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 20115 16692 20181 16693
rect 20115 16628 20116 16692
rect 20180 16628 20181 16692
rect 20115 16627 20181 16628
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 17907 14788 17973 14789
rect 17907 14724 17908 14788
rect 17972 14724 17973 14788
rect 17907 14723 17973 14724
rect 17723 13156 17789 13157
rect 17723 13092 17724 13156
rect 17788 13092 17789 13156
rect 17723 13091 17789 13092
rect 17539 12204 17605 12205
rect 17539 12140 17540 12204
rect 17604 12140 17605 12204
rect 17539 12139 17605 12140
rect 17355 9212 17421 9213
rect 17355 9148 17356 9212
rect 17420 9148 17421 9212
rect 17355 9147 17421 9148
rect 17542 6901 17602 12139
rect 17726 9346 17786 13091
rect 17910 10845 17970 14723
rect 19137 14720 19457 15744
rect 19747 15332 19813 15333
rect 19747 15268 19748 15332
rect 19812 15268 19813 15332
rect 19747 15267 19813 15268
rect 19931 15332 19997 15333
rect 19931 15268 19932 15332
rect 19996 15268 19997 15332
rect 19931 15267 19997 15268
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 18275 14516 18341 14517
rect 18275 14452 18276 14516
rect 18340 14452 18341 14516
rect 18275 14451 18341 14452
rect 18091 13836 18157 13837
rect 18091 13772 18092 13836
rect 18156 13772 18157 13836
rect 18091 13771 18157 13772
rect 17907 10844 17973 10845
rect 17907 10780 17908 10844
rect 17972 10780 17973 10844
rect 17907 10779 17973 10780
rect 17726 9286 17924 9346
rect 17723 9212 17789 9213
rect 17723 9148 17724 9212
rect 17788 9148 17789 9212
rect 17723 9147 17789 9148
rect 17726 7717 17786 9147
rect 17864 8310 17924 9286
rect 18094 8941 18154 13771
rect 18091 8940 18157 8941
rect 18091 8876 18092 8940
rect 18156 8876 18157 8940
rect 18091 8875 18157 8876
rect 17864 8250 17970 8310
rect 17910 7853 17970 8250
rect 17907 7852 17973 7853
rect 17907 7788 17908 7852
rect 17972 7788 17973 7852
rect 17907 7787 17973 7788
rect 18278 7717 18338 14451
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 18827 11116 18893 11117
rect 18827 11052 18828 11116
rect 18892 11052 18893 11116
rect 18827 11051 18893 11052
rect 18643 8124 18709 8125
rect 18643 8060 18644 8124
rect 18708 8060 18709 8124
rect 18643 8059 18709 8060
rect 17723 7716 17789 7717
rect 17723 7652 17724 7716
rect 17788 7652 17789 7716
rect 17723 7651 17789 7652
rect 18275 7716 18341 7717
rect 18275 7652 18276 7716
rect 18340 7652 18341 7716
rect 18275 7651 18341 7652
rect 17907 7444 17973 7445
rect 17907 7380 17908 7444
rect 17972 7380 17973 7444
rect 17907 7379 17973 7380
rect 17539 6900 17605 6901
rect 17539 6836 17540 6900
rect 17604 6836 17605 6900
rect 17539 6835 17605 6836
rect 17910 6221 17970 7379
rect 18278 7173 18338 7651
rect 18275 7172 18341 7173
rect 18275 7108 18276 7172
rect 18340 7108 18341 7172
rect 18275 7107 18341 7108
rect 17907 6220 17973 6221
rect 17907 6156 17908 6220
rect 17972 6156 17973 6220
rect 17907 6155 17973 6156
rect 18646 6085 18706 8059
rect 18830 7989 18890 11051
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19750 8397 19810 15267
rect 19934 11117 19994 15267
rect 19931 11116 19997 11117
rect 19931 11052 19932 11116
rect 19996 11052 19997 11116
rect 19931 11051 19997 11052
rect 19931 10572 19997 10573
rect 19931 10508 19932 10572
rect 19996 10508 19997 10572
rect 19931 10507 19997 10508
rect 19747 8396 19813 8397
rect 19747 8332 19748 8396
rect 19812 8332 19813 8396
rect 19747 8331 19813 8332
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 18827 7988 18893 7989
rect 18827 7924 18828 7988
rect 18892 7924 18893 7988
rect 18827 7923 18893 7924
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 18643 6084 18709 6085
rect 18643 6020 18644 6084
rect 18708 6020 18709 6084
rect 18643 6019 18709 6020
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 17171 5948 17237 5949
rect 17171 5884 17172 5948
rect 17236 5884 17237 5948
rect 17171 5883 17237 5884
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16067 4996 16133 4997
rect 16067 4932 16068 4996
rect 16132 4932 16133 4996
rect 16067 4931 16133 4932
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 15699 4316 15765 4317
rect 15699 4252 15700 4316
rect 15764 4252 15765 4316
rect 15699 4251 15765 4252
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 4928 19457 5952
rect 19934 5405 19994 10507
rect 20118 6765 20178 16627
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 20115 6764 20181 6765
rect 20115 6700 20116 6764
rect 20180 6700 20181 6764
rect 20115 6699 20181 6700
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 19931 5404 19997 5405
rect 19931 5340 19932 5404
rect 19996 5340 19997 5404
rect 19931 5339 19997 5340
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform -1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform -1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 6624 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform -1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 3128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 9200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 7912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 9200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 9568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 3496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 4968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 3864 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 7728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 1932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 2024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 2300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5060 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9384 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17112 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 2024 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 2392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1649977179
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1649977179
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_12
timestamp 1649977179
transform 1 0 2208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1649977179
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_67
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1649977179
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1649977179
transform 1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1649977179
transform 1 0 13248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1649977179
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_100
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_104
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_114
timestamp 1649977179
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1649977179
transform 1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_17
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_65
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1649977179
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1649977179
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1649977179
transform 1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1649977179
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_148
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_194
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_198
timestamp 1649977179
transform 1 0 19320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1649977179
transform 1 0 7636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1649977179
transform 1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_179
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1649977179
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_124
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1649977179
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1649977179
transform 1 0 14720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_107
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_200
timestamp 1649977179
transform 1 0 19504 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_74
timestamp 1649977179
transform 1 0 7912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_92
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_114
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_150
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_211
timestamp 1649977179
transform 1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_216
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1649977179
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_130
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_191
timestamp 1649977179
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1649977179
transform 1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_129
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_160
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1649977179
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1649977179
transform 1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1649977179
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_60
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_119
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1649977179
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_199
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_210
timestamp 1649977179
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_151
timestamp 1649977179
transform 1 0 14996 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_168
timestamp 1649977179
transform 1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_178
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1649977179
transform 1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1649977179
transform 1 0 7544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1649977179
transform 1 0 7912 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_150
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_200
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1649977179
transform 1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_87
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1649977179
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1649977179
transform 1 0 17296 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1649977179
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_206
timestamp 1649977179
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_73
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_85
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_104
timestamp 1649977179
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_119
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1649977179
transform 1 0 17296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_63
timestamp 1649977179
transform 1 0 6900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_184
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_119
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1649977179
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1649977179
transform 1 0 10672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1649977179
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1649977179
transform 1 0 12696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1649977179
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1649977179
transform 1 0 14628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_35
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_82
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1649977179
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1649977179
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1649977179
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1649977179
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1649977179
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_40
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1649977179
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_63
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_91
timestamp 1649977179
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_86
timestamp 1649977179
transform 1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_55
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_124
timestamp 1649977179
transform 1 0 12512 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1649977179
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1649977179
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_64
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_68
timestamp 1649977179
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_76
timestamp 1649977179
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1649977179
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1649977179
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_117
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1649977179
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_130
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1649977179
transform 1 0 15824 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1649977179
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_34
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_38
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_42
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_46
timestamp 1649977179
transform 1 0 5336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_50
timestamp 1649977179
transform 1 0 5704 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_54
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_58
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_75
timestamp 1649977179
transform 1 0 8004 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_92
timestamp 1649977179
transform 1 0 9568 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_144
timestamp 1649977179
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_202
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_5
timestamp 1649977179
transform 1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_18
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_22
timestamp 1649977179
transform 1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1649977179
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_46
timestamp 1649977179
transform 1 0 5336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_50
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1649977179
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_78
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1649977179
transform 1 0 10488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_117
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_122
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_6
timestamp 1649977179
transform 1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1649977179
transform 1 0 2024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_33
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_45
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1649977179
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1649977179
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_6
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_10
timestamp 1649977179
transform 1 0 2024 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1649977179
transform 1 0 2392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_22
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1649977179
transform 1 0 3496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1649977179
transform 1 0 3864 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_70
timestamp 1649977179
transform 1 0 7544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1649977179
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_8
timestamp 1649977179
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1649977179
transform 1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_63
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1649977179
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_132
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1649977179
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_183
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_216
timestamp 1649977179
transform 1 0 20976 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1649977179
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1649977179
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform -1 0 18952 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform -1 0 18400 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform -1 0 20240 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform -1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform -1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform -1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 18216 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 11868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 12328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 8464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 6072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 8004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 17756 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 14904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform 1 0 17296 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 13800 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 20148 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 4324 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform -1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1649977179
transform -1 0 3496 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 5060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1649977179
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform -1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1649977179
transform -1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform -1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1649977179
transform 1 0 20516 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform -1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15640 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15824 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13524 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11224 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10488 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10856 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13984 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9568 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12880 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16100 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20148 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14812 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14352 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12144 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15180 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18584 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20332 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19504 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_1__155 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11500 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12604 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16100 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_1__158
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_1__160
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_1__161
timestamp 1649977179
transform -1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_1__156
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__157
timestamp 1649977179
transform -1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l1_in_1__159
timestamp 1649977179
transform -1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15916 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__162
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10120 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5796 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform -1 0 9844 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l1_in_3__135
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l1_in_3__145
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5704 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6900 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l1_in_3__146
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5888 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8188 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_1__147
timestamp 1649977179
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_1__163
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_1__164
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5888 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8648 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9200 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_1__165
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9936 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10672 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_1__133
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16560 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l1_in_1__134
timestamp 1649977179
transform -1 0 16928 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18952 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18676 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l1_in_1__136
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20240 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l1_in_1__137
timestamp 1649977179
transform -1 0 20424 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20056 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l2_in_1__138
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17388 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__139
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__140
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__141
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__142
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__143
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__144
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_1__148
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_1__150
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_1__153
timestamp 1649977179
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7636 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_1__154
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6992 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18492 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_1__149
timestamp 1649977179
transform -1 0 19780 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_1__151
timestamp 1649977179
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10212 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l2_in_1__152
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18768 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output72 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 18952 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 18952 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform -1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_1_
port 2 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 5 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 6 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 7 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 8 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 9 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 10 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 11 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 12 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 13 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 14 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 15 nsew signal input
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 16 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 17 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 18 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 19 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 20 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 21 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 22 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 23 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 24 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 25 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 26 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 27 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 28 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 29 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 30 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 31 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 32 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 33 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 34 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 35 nsew signal tristate
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 36 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 37 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 38 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 39 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 40 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 41 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 42 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 43 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 44 nsew signal tristate
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 45 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 46 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 47 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 48 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 49 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 50 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 51 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 52 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 53 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 54 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 55 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 56 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 57 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 58 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 59 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 60 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 61 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 62 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 63 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 64 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 65 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 66 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 67 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 68 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 69 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 70 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 71 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 72 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 73 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 74 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 75 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 76 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 77 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 78 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 79 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 80 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 81 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 82 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 83 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 84 nsew signal tristate
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 85 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 86 nsew signal input
flabel metal2 s 7010 22200 7066 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 87 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 88 nsew signal input
flabel metal2 s 8114 22200 8170 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 89 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 90 nsew signal input
flabel metal2 s 9218 22200 9274 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 91 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 92 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 93 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 94 nsew signal input
flabel metal2 s 11426 22200 11482 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 95 nsew signal input
flabel metal2 s 1490 22200 1546 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 96 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 97 nsew signal input
flabel metal2 s 2594 22200 2650 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 98 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 99 nsew signal input
flabel metal2 s 3698 22200 3754 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 100 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 101 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 102 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 103 nsew signal input
flabel metal2 s 5906 22200 5962 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 104 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 105 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 106 nsew signal tristate
flabel metal2 s 18050 22200 18106 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 107 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 108 nsew signal tristate
flabel metal2 s 19154 22200 19210 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 109 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 110 nsew signal tristate
flabel metal2 s 20258 22200 20314 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 111 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 112 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 113 nsew signal tristate
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 114 nsew signal tristate
flabel metal2 s 22466 22200 22522 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 115 nsew signal tristate
flabel metal2 s 12530 22200 12586 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 116 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 117 nsew signal tristate
flabel metal2 s 13634 22200 13690 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 118 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 119 nsew signal tristate
flabel metal2 s 14738 22200 14794 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 120 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 121 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 122 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 123 nsew signal tristate
flabel metal2 s 16946 22200 17002 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 124 nsew signal tristate
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 125 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 126 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 127 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 128 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 129 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 130 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 131 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 132 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 133 nsew signal input
flabel metal2 s 386 22200 442 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_1_
port 134 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
