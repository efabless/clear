VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_array
  CLASS BLOCK ;
  FOREIGN tie_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 70.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.960 10.640 18.560 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.200 10.640 30.800 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.440 10.640 43.040 57.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.840 10.640 12.440 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.080 10.640 24.680 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.320 10.640 36.920 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.560 10.640 49.160 57.360 ;
    END
  END VPWR
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END x[7]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 57.205 ;
      LAYER met1 ;
        RECT 3.750 10.640 55.590 57.360 ;
      LAYER met2 ;
        RECT 3.780 4.280 55.560 57.305 ;
        RECT 4.330 3.670 10.850 4.280 ;
        RECT 11.690 3.670 18.210 4.280 ;
        RECT 19.050 3.670 25.570 4.280 ;
        RECT 26.410 3.670 32.930 4.280 ;
        RECT 33.770 3.670 40.290 4.280 ;
        RECT 41.130 3.670 47.650 4.280 ;
        RECT 48.490 3.670 55.010 4.280 ;
      LAYER met3 ;
        RECT 10.850 10.715 49.150 57.285 ;
  END
END tie_array
END LIBRARY

