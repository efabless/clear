magic
tech sky130A
magscale 1 2
timestamp 1625784763
<< obsli1 >>
rect 1104 2159 22051 20689
<< obsm1 >>
rect 198 1164 22802 20720
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< obsm2 >>
rect 204 22144 5666 22681
rect 5834 22144 17166 22681
rect 17334 22144 22796 22681
rect 204 856 22796 22144
rect 314 167 514 856
rect 682 167 974 856
rect 1142 167 1434 856
rect 1602 167 1894 856
rect 2062 167 2354 856
rect 2522 167 2814 856
rect 2982 167 3274 856
rect 3442 167 3734 856
rect 3902 167 4194 856
rect 4362 167 4654 856
rect 4822 167 5022 856
rect 5190 167 5482 856
rect 5650 167 5942 856
rect 6110 167 6402 856
rect 6570 167 6862 856
rect 7030 167 7322 856
rect 7490 167 7782 856
rect 7950 167 8242 856
rect 8410 167 8702 856
rect 8870 167 9162 856
rect 9330 167 9530 856
rect 9698 167 9990 856
rect 10158 167 10450 856
rect 10618 167 10910 856
rect 11078 167 11370 856
rect 11538 167 11830 856
rect 11998 167 12290 856
rect 12458 167 12750 856
rect 12918 167 13210 856
rect 13378 167 13670 856
rect 13838 167 14038 856
rect 14206 167 14498 856
rect 14666 167 14958 856
rect 15126 167 15418 856
rect 15586 167 15878 856
rect 16046 167 16338 856
rect 16506 167 16798 856
rect 16966 167 17258 856
rect 17426 167 17718 856
rect 17886 167 18178 856
rect 18346 167 18546 856
rect 18714 167 19006 856
rect 19174 167 19466 856
rect 19634 167 19926 856
rect 20094 167 20386 856
rect 20554 167 20846 856
rect 21014 167 21306 856
rect 21474 167 21766 856
rect 21934 167 22226 856
rect 22394 167 22686 856
<< metal3 >>
rect 0 22584 800 22704
rect 22200 22584 23000 22704
rect 0 22176 800 22296
rect 22200 22176 23000 22296
rect 0 21632 800 21752
rect 22200 21632 23000 21752
rect 0 21224 800 21344
rect 22200 21224 23000 21344
rect 0 20680 800 20800
rect 22200 20680 23000 20800
rect 0 20272 800 20392
rect 22200 20272 23000 20392
rect 0 19728 800 19848
rect 22200 19728 23000 19848
rect 0 19320 800 19440
rect 22200 19320 23000 19440
rect 0 18776 800 18896
rect 22200 18776 23000 18896
rect 0 18368 800 18488
rect 22200 18368 23000 18488
rect 0 17960 800 18080
rect 22200 17960 23000 18080
rect 0 17416 800 17536
rect 22200 17416 23000 17536
rect 0 17008 800 17128
rect 22200 17008 23000 17128
rect 0 16464 800 16584
rect 22200 16464 23000 16584
rect 0 16056 800 16176
rect 22200 16056 23000 16176
rect 0 15512 800 15632
rect 22200 15512 23000 15632
rect 0 15104 800 15224
rect 22200 15104 23000 15224
rect 0 14560 800 14680
rect 22200 14560 23000 14680
rect 0 14152 800 14272
rect 22200 14152 23000 14272
rect 0 13744 800 13864
rect 22200 13744 23000 13864
rect 0 13200 800 13320
rect 22200 13200 23000 13320
rect 0 12792 800 12912
rect 22200 12792 23000 12912
rect 0 12248 800 12368
rect 22200 12248 23000 12368
rect 0 11840 800 11960
rect 22200 11840 23000 11960
rect 0 11296 800 11416
rect 22200 11296 23000 11416
rect 0 10888 800 11008
rect 22200 10888 23000 11008
rect 0 10344 800 10464
rect 22200 10344 23000 10464
rect 0 9936 800 10056
rect 22200 9936 23000 10056
rect 0 9392 800 9512
rect 22200 9392 23000 9512
rect 0 8984 800 9104
rect 22200 8984 23000 9104
rect 0 8576 800 8696
rect 22200 8576 23000 8696
rect 0 8032 800 8152
rect 22200 8032 23000 8152
rect 0 7624 800 7744
rect 22200 7624 23000 7744
rect 0 7080 800 7200
rect 22200 7080 23000 7200
rect 0 6672 800 6792
rect 22200 6672 23000 6792
rect 0 6128 800 6248
rect 22200 6128 23000 6248
rect 0 5720 800 5840
rect 22200 5720 23000 5840
rect 0 5176 800 5296
rect 22200 5176 23000 5296
rect 0 4768 800 4888
rect 22200 4768 23000 4888
rect 0 4360 800 4480
rect 22200 4360 23000 4480
rect 0 3816 800 3936
rect 22200 3816 23000 3936
rect 0 3408 800 3528
rect 22200 3408 23000 3528
rect 0 2864 800 2984
rect 22200 2864 23000 2984
rect 0 2456 800 2576
rect 22200 2456 23000 2576
rect 0 1912 800 2032
rect 22200 1912 23000 2032
rect 0 1504 800 1624
rect 22200 1504 23000 1624
rect 0 960 800 1080
rect 22200 960 23000 1080
rect 0 552 800 672
rect 22200 552 23000 672
rect 0 144 800 264
rect 22200 144 23000 264
<< obsm3 >>
rect 880 22504 22120 22677
rect 800 22376 22200 22504
rect 880 22096 22120 22376
rect 800 21832 22200 22096
rect 880 21552 22120 21832
rect 800 21424 22200 21552
rect 880 21144 22120 21424
rect 800 20880 22200 21144
rect 880 20600 22120 20880
rect 800 20472 22200 20600
rect 880 20192 22120 20472
rect 800 19928 22200 20192
rect 880 19648 22120 19928
rect 800 19520 22200 19648
rect 880 19240 22120 19520
rect 800 18976 22200 19240
rect 880 18696 22120 18976
rect 800 18568 22200 18696
rect 880 18288 22120 18568
rect 800 18160 22200 18288
rect 880 17880 22120 18160
rect 800 17616 22200 17880
rect 880 17336 22120 17616
rect 800 17208 22200 17336
rect 880 16928 22120 17208
rect 800 16664 22200 16928
rect 880 16384 22120 16664
rect 800 16256 22200 16384
rect 880 15976 22120 16256
rect 800 15712 22200 15976
rect 880 15432 22120 15712
rect 800 15304 22200 15432
rect 880 15024 22120 15304
rect 800 14760 22200 15024
rect 880 14480 22120 14760
rect 800 14352 22200 14480
rect 880 14072 22120 14352
rect 800 13944 22200 14072
rect 880 13664 22120 13944
rect 800 13400 22200 13664
rect 880 13120 22120 13400
rect 800 12992 22200 13120
rect 880 12712 22120 12992
rect 800 12448 22200 12712
rect 880 12168 22120 12448
rect 800 12040 22200 12168
rect 880 11760 22120 12040
rect 800 11496 22200 11760
rect 880 11216 22120 11496
rect 800 11088 22200 11216
rect 880 10808 22120 11088
rect 800 10544 22200 10808
rect 880 10264 22120 10544
rect 800 10136 22200 10264
rect 880 9856 22120 10136
rect 800 9592 22200 9856
rect 880 9312 22120 9592
rect 800 9184 22200 9312
rect 880 8904 22120 9184
rect 800 8776 22200 8904
rect 880 8496 22120 8776
rect 800 8232 22200 8496
rect 880 7952 22120 8232
rect 800 7824 22200 7952
rect 880 7544 22120 7824
rect 800 7280 22200 7544
rect 880 7000 22120 7280
rect 800 6872 22200 7000
rect 880 6592 22120 6872
rect 800 6328 22200 6592
rect 880 6048 22120 6328
rect 800 5920 22200 6048
rect 880 5640 22120 5920
rect 800 5376 22200 5640
rect 880 5096 22120 5376
rect 800 4968 22200 5096
rect 880 4688 22120 4968
rect 800 4560 22200 4688
rect 880 4280 22120 4560
rect 800 4016 22200 4280
rect 880 3736 22120 4016
rect 800 3608 22200 3736
rect 880 3328 22120 3608
rect 800 3064 22200 3328
rect 880 2784 22120 3064
rect 800 2656 22200 2784
rect 880 2376 22120 2656
rect 800 2112 22200 2376
rect 880 1832 22120 2112
rect 800 1704 22200 1832
rect 880 1424 22120 1704
rect 800 1160 22200 1424
rect 880 880 22120 1160
rect 800 752 22200 880
rect 880 472 22120 752
rect 800 344 22200 472
rect 880 171 22120 344
<< metal4 >>
rect 4409 2128 4729 20720
rect 7875 2128 8195 20720
rect 11340 2128 11660 20720
rect 14805 2128 15125 20720
rect 18271 2128 18591 20720
<< obsm4 >>
rect 3187 2128 4329 20720
rect 4809 2128 7795 20720
rect 8275 2128 11260 20720
rect 11740 2128 14725 20720
rect 15205 2128 18191 20720
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 2 nsew signal output
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 3 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 4 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 5 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 6 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 7 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 8 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 bottom_left_grid_pin_48_
port 9 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_49_
port 10 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 ccff_head
port 11 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_tail
port 12 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 13 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 14 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 15 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 16 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 17 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 18 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 19 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 20 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 21 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 22 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 24 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 25 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 26 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 27 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 28 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 29 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 30 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 31 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 32 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 33 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 34 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 35 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 36 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 37 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 38 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 39 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 40 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 41 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 42 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 43 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 44 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 45 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 46 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 47 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 48 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 49 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 50 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 51 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 52 nsew signal output
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 53 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 54 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 55 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 56 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 57 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 58 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 59 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 60 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 61 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 62 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 63 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 64 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 65 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 66 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 67 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 68 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 69 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 70 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 71 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 72 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 73 nsew signal output
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 74 nsew signal output
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 75 nsew signal output
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 76 nsew signal output
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 77 nsew signal output
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 78 nsew signal output
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 79 nsew signal output
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 80 nsew signal output
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 81 nsew signal output
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 82 nsew signal output
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 83 nsew signal output
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 84 nsew signal output
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 85 nsew signal output
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 86 nsew signal output
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 87 nsew signal output
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 88 nsew signal output
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 89 nsew signal output
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 90 nsew signal output
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 91 nsew signal output
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 92 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_in[0]
port 93 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[10]
port 94 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[11]
port 95 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[12]
port 96 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[13]
port 97 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[14]
port 98 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[15]
port 99 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[16]
port 100 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 101 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 102 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[19]
port 103 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[1]
port 104 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[2]
port 105 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[3]
port 106 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[4]
port 107 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[5]
port 108 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[6]
port 109 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[7]
port 110 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[8]
port 111 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[9]
port 112 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_out[0]
port 113 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[10]
port 114 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 chany_bottom_out[11]
port 115 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 116 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[13]
port 117 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[14]
port 118 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[15]
port 119 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 chany_bottom_out[16]
port 120 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[17]
port 121 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[18]
port 122 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[19]
port 123 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[1]
port 124 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[2]
port 125 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_out[3]
port 126 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[4]
port 127 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_out[5]
port 128 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[6]
port 129 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 130 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 131 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[9]
port 132 nsew signal output
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 133 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 134 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 135 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 136 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 137 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 138 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 139 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 140 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 141 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 142 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 143 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 144 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 145 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 146 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 147 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 148 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 149 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 150 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 151 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 152 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 153 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 154 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 155 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 156 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 23000 23000
string LEFview TRUE
string GDS_FILE /project/openlane/sb_1__2_/runs/sb_1__2_/results/magic/sb_1__2_.gds
string GDS_END 1572414
string GDS_START 100992
<< end >>

