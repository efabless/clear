* NGSPICE file created from sb_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__1_ VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_
+ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_
+ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ prog_clk_0_N_in top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ top_right_grid_pin_1_
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l1_in_2__S mux_top_track_16.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_44_ bottom_left_grid_pin_42_
+ mux_bottom_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_15.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_35.mux_l1_in_0__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__124__A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_062_ VGND VGND VPWR VPWR _062_/HI _062_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__119__A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
X_114_ _114_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_061_ VGND VGND VPWR VPWR _061_/HI _061_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _070_/A sky130_fd_sc_hd__buf_4
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_113_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.mux_l1_in_3_ _046_/HI left_bottom_grid_pin_41_ mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_15.mux_l3_in_0_ mux_left_track_15.mux_l2_in_1_/X mux_left_track_15.mux_l2_in_0_/X
+ mux_left_track_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_0.mux_l2_in_3_ _048_/HI chanx_left_in[14] mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l2_in_1_ _065_/HI left_bottom_grid_pin_37_ mux_left_track_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l1_in_3__S mux_top_track_24.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_060_ VGND VGND VPWR VPWR _060_/HI _060_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l1_in_3_/X mux_left_track_7.mux_l1_in_2_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
X_112_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.mux_l1_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[7] chanx_left_in[0] mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_15.mux_l2_in_0_ chany_bottom_in[19] mux_left_track_15.mux_l1_in_0_/X
+ mux_left_track_15.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
X_111_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_3.mux_l1_in_3__S mux_left_track_3.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_7.mux_l1_in_1_ left_bottom_grid_pin_35_ chany_bottom_in[6] mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_11.mux_l2_in_0__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[2] top_right_grid_pin_1_ mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _114_/A sky130_fd_sc_hd__buf_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_15.mux_l1_in_0_ chany_bottom_in[12] chany_top_in[12] mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ _110_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l2_in_3_ _061_/HI chanx_left_in[18] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_7.mux_l1_in_0_ chany_bottom_in[3] chany_top_in[6] mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__buf_4
XFILLER_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chany_top_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__091__A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_5__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_3__S mux_bottom_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_39.mux_l2_in_0_ _044_/HI mux_left_track_39.mux_l1_in_0_/X ccff_tail
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__buf_4
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chany_top_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__089__A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 bottom_right_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_1_ _057_/HI mux_bottom_track_25.mux_l1_in_2_/X mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_5__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__097__A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l1_in_2_ chanx_left_in[13] chanx_left_in[6] mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_9.mux_l2_in_1_ bottom_left_grid_pin_49_ bottom_left_grid_pin_45_
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_23.mux_l1_in_0__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_2.mux_l2_in_3__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_15.mux_l1_in_0__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_39.mux_l1_in_0_ left_bottom_grid_pin_41_ chany_top_in[1] mux_left_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_5__A1 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_098_ _098_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_13.mux_l2_in_1__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_43_
+ mux_bottom_track_25.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_track_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_0_ bottom_right_grid_pin_1_ mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_31.mux_l1_in_0__A0 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chany_top_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_3_ _049_/HI chanx_left_in[17] mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_23.mux_l1_in_0__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _068_/A sky130_fd_sc_hd__buf_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_3.mux_l1_in_3_ _039_/HI left_bottom_grid_pin_41_ mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_4.mux_l1_in_5__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l1_in_1__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_4__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_097_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xmux_left_track_11.mux_l3_in_0_ mux_left_track_11.mux_l2_in_1_/X mux_left_track_11.mux_l2_in_0_/X
+ mux_left_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l2_in_1_ mux_top_track_16.mux_l1_in_3_/X mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_2__S mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_31.mux_l1_in_0__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_11.mux_l2_in_1_ _063_/HI left_bottom_grid_pin_35_ mux_left_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_ chanx_left_in[10] chanx_left_in[3] mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_3__A1 chanx_left_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_13.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__100__A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A1 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_5__A1 chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l1_in_6_ chanx_left_in[17] chanx_left_in[10] mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_079_ left_bottom_grid_pin_35_ VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_11.mux_l2_in_0_ chany_bottom_in[11] mux_left_track_11.mux_l1_in_0_/X
+ mux_left_track_11.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[17] chany_bottom_in[8] mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__buf_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__103__A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_33.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_1_ left_bottom_grid_pin_35_ chany_bottom_in[4] mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_095_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__111__A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_6_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_5_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ _078_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ top_left_grid_pin_47_ top_left_grid_pin_43_ mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ chany_bottom_in[9] chany_top_in[9] mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l1_in_1_/X mux_left_track_23.mux_l1_in_0_/X
+ mux_left_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_3_ _060_/HI mux_bottom_track_5.mux_l1_in_6_/X mux_bottom_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__109__A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chany_bottom_in[0] chany_top_in[4] mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_23.mux_l1_in_1_ _036_/HI left_bottom_grid_pin_41_ mux_left_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_094_ _094_/A VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_4_ bottom_left_grid_pin_48_ bottom_left_grid_pin_47_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_4_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__117__A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_29.mux_l1_in_0__A0 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_3__A1 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_3__S mux_top_track_16.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.mux_l2_in_2_ mux_bottom_track_5.mux_l1_in_5_/X mux_bottom_track_5.mux_l1_in_4_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__125__A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_23.mux_l1_in_0_ chany_bottom_in[17] chany_top_in[17] mux_left_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_093_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xmux_left_track_35.mux_l2_in_0_ _042_/HI mux_left_track_35.mux_l1_in_0_/X mux_left_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_3_ bottom_left_grid_pin_46_ bottom_left_grid_pin_45_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_076_ _076_/A VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_37.mux_l1_in_0__A0 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ VGND VGND VPWR VPWR _059_/HI _059_/LO sky130_fd_sc_hd__conb_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_29.mux_l1_in_0__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_092_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_44_ bottom_left_grid_pin_43_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_075_ _075_/A VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_37.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_35.mux_l1_in_0_ left_bottom_grid_pin_39_ chany_top_in[7] mux_left_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_058_ VGND VGND VPWR VPWR _058_/HI _058_/LO sky130_fd_sc_hd__conb_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l2_in_1_ _059_/HI mux_bottom_track_33.mux_l1_in_2_/X mux_bottom_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _066_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_091_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_42_ bottom_right_grid_pin_1_
+ mux_bottom_track_5.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_2_ chanx_left_in[14] chanx_left_in[7] mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_11.mux_l1_in_0__A0 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_074_ _074_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_057_ VGND VGND VPWR VPWR _057_/HI _057_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_right_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_090_ _090_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__buf_4
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_33.mux_l1_in_1_ chanx_left_in[0] bottom_left_grid_pin_48_ mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_11.mux_l1_in_0__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_125_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
X_056_ VGND VGND VPWR VPWR _056_/HI _056_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_3_ _051_/HI chanx_left_in[16] mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_6_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_2.mux_l2_in_3_ _050_/HI chanx_left_in[13] mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_1_ mux_top_track_24.mux_l1_in_3_/X mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_33.mux_l1_in_0_ bottom_left_grid_pin_44_ chany_top_in[10] mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_2_ chanx_left_in[9] chanx_left_in[2] mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
X_107_ _107_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_2.mux_l2_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_1_ _047_/HI left_bottom_grid_pin_34_ mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__079__A left_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_5.mux_l1_in_3__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_4__A0 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_2__S mux_bottom_track_17.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_5 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__092__A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[13] mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0__A0 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_6__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
X_123_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_1_ chany_bottom_in[18] chany_bottom_in[9] mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 top_left_grid_pin_47_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l2_in_3_ _055_/HI chanx_left_in[15] mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1_ _033_/HI left_bottom_grid_pin_38_ mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_106_ _106_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[8] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A1 chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__095__A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_4__A1 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ chany_bottom_in[4] top_left_grid_pin_49_ mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_070_ _070_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l1_in_3__A1 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
X_122_ _122_/A VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_0_ top_left_grid_pin_48_ top_left_grid_pin_44_ mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_2_ chanx_left_in[8] chanx_left_in[1] mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_105_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A0 chanx_left_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chany_bottom_in[13] chany_top_in[13] mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_21.mux_l1_in_1__A1 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.mux_l2_in_0_ _038_/HI mux_left_track_29.mux_l1_in_0_/X mux_left_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_31.mux_l2_in_0_ _040_/HI mux_left_track_31.mux_l1_in_0_/X mux_left_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_9.mux_l1_in_0_ chany_bottom_in[7] chany_top_in[8] mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_4.mux_l1_in_4__A0 chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l2_in_0_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_44_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A0 chanx_left_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_121_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l2_in_1_ bottom_left_grid_pin_49_ mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_104_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A0 chanx_left_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_29.mux_l1_in_0_ left_bottom_grid_pin_36_ chany_top_in[19] mux_left_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_4__A1 top_right_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_45_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_31.mux_l1_in_0_ left_bottom_grid_pin_37_ chany_top_in[15] mux_left_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_5__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_3__S mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
X_120_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_103_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_33.mux_l1_in_1__S mux_bottom_track_33.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_15.mux_l2_in_1__A1 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_43_ bottom_right_grid_pin_1_
+ mux_bottom_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__101__A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X ccff_head VGND VGND
+ VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_16.mux_l1_in_3__A1 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__buf_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ _102_/A VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_2__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__104__A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l1_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__112__A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l1_in_3__S mux_left_track_1.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_3_ _045_/HI left_bottom_grid_pin_40_ mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_13.mux_l3_in_0_ mux_left_track_13.mux_l2_in_1_/X mux_left_track_13.mux_l2_in_0_/X
+ mux_left_track_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__120__A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__buf_4
XANTENNA__115__A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_19.mux_l1_in_1__A1 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.mux_l2_in_1_ _064_/HI left_bottom_grid_pin_36_ mux_left_track_13.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_13.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_7.mux_l1_in_3__A1 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__123__A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_100_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_right_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_3_ _054_/HI chanx_left_in[18] mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_13.mux_l2_in_0_ chany_bottom_in[15] mux_left_track_13.mux_l1_in_0_/X
+ mux_left_track_13.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_32.mux_l2_in_1_ _052_/HI mux_top_track_32.mux_l1_in_2_/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.mux_l1_in_2_ chanx_left_in[15] chanx_left_in[8] mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[5] mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_13.mux_l1_in_0_ chany_bottom_in[10] chany_top_in[10] mux_left_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l1_in_2__S mux_top_track_24.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_1_ chanx_left_in[1] chany_bottom_in[10] mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ chany_bottom_in[1] chany_top_in[5] mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_1_ _037_/HI left_bottom_grid_pin_34_ mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 top_left_grid_pin_46_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_39.mux_l1_in_0__A0 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_32.mux_l1_in_0_ top_left_grid_pin_49_ top_left_grid_pin_45_ mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_25.mux_l1_in_0_ chany_bottom_in[18] chany_top_in[18] mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_088_ _088_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_37.mux_l2_in_0_ _043_/HI mux_left_track_37.mux_l1_in_0_/X mux_left_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A1 chanx_left_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_8.mux_l2_in_0_ top_right_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_39.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_2__S mux_left_track_3.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_43_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _110_/A sky130_fd_sc_hd__buf_4
XFILLER_32_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ _087_/A VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A0 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_37.mux_l1_in_0_ left_bottom_grid_pin_40_ chany_top_in[3] mux_left_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_42_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l1_in_0_ top_left_grid_pin_46_ top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _067_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_069_ _069_/A VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A1 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_4__S mux_bottom_track_5.mux_l1_in_6_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_6_ chanx_left_in[19] chanx_left_in[12] mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__S mux_bottom_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_3__S mux_bottom_track_17.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_3_ _062_/HI left_bottom_grid_pin_40_ mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_1__A1 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_21.mux_l1_in_0__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ _068_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__096__A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_5_ chanx_left_in[5] chany_bottom_in[14] mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_3__A0 top_left_grid_pin_49_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_3_ _053_/HI mux_top_track_4.mux_l1_in_6_/X mux_top_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_6__A0 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_067_ _067_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_15.mux_l2_in_0__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__buf_4
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_4_ chany_bottom_in[5] top_right_grid_pin_1_ mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 top_left_grid_pin_48_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_5.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A0 chanx_left_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l1_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[2] mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l1_in_2__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ _083_/A VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_2_ mux_top_track_4.mux_l1_in_5_/X mux_top_track_4.mux_l1_in_4_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_6__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_066_ _066_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l1_in_1_/X mux_left_track_19.mux_l1_in_0_/X
+ mux_left_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_3_ top_left_grid_pin_49_ top_left_grid_pin_48_ mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
X_118_ _118_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l1_in_1_/X mux_left_track_21.mux_l1_in_0_/X
+ mux_left_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_2__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A1 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_3_ _058_/HI chanx_left_in[16] mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_19.mux_l1_in_1_ _034_/HI left_bottom_grid_pin_39_ mux_left_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[2] chany_top_in[0] mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_2__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_21.mux_l1_in_1_ _035_/HI left_bottom_grid_pin_40_ mux_left_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_23.mux_l1_in_1__A1 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_6__S mux_top_track_4.mux_l1_in_6_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ _082_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _122_/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_065_ VGND VGND VPWR VPWR _065_/HI _065_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_33.mux_l1_in_2__S mux_bottom_track_33.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_6__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_32.mux_l1_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_2_ top_left_grid_pin_47_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_117_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_17.mux_l1_in_3_ _056_/HI chanx_left_in[19] mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_2__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_2_ chanx_left_in[9] chanx_left_in[2] mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_19.mux_l1_in_0_ chany_bottom_in[14] chany_top_in[14] mux_left_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_21.mux_l1_in_0_ chany_bottom_in[16] chany_top_in[16] mux_left_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ _041_/HI mux_left_track_33.mux_l1_in_0_/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_7.mux_l1_in_2__A0 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_081_ _081_/A VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__buf_4
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ VGND VGND VPWR VPWR _064_/HI _064_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_1_ mux_bottom_track_17.mux_l1_in_3_/X mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_4.mux_l1_in_6__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_45_ top_left_grid_pin_44_ mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__105__A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_116_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_17.mux_l1_in_2_ chanx_left_in[12] chanx_left_in[5] mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_1_ bottom_left_grid_pin_48_ bottom_left_grid_pin_46_
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_7.mux_l1_in_2__A1 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__113__A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_35.mux_l1_in_0__A0 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_080_ _080_/A VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_0_ left_bottom_grid_pin_38_ chany_top_in[11] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_063_ VGND VGND VPWR VPWR _063_/HI _063_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_43_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
X_115_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__121__A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_42_
+ mux_bottom_track_17.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__116__A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

