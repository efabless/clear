magic
tech sky130A
magscale 1 2
timestamp 1656406101
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 14 8 22986 21276
<< metal2 >>
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8666 22200 8722 23000
rect 9034 22200 9090 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 21546 22200 21602 23000
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
<< obsm2 >>
rect 20 22144 514 22273
rect 682 22144 882 22273
rect 1050 22144 1250 22273
rect 1418 22144 1618 22273
rect 1786 22144 1986 22273
rect 2154 22144 2354 22273
rect 2522 22144 2722 22273
rect 2890 22144 3090 22273
rect 3258 22144 3458 22273
rect 3626 22144 3826 22273
rect 3994 22144 4194 22273
rect 4362 22144 4562 22273
rect 4730 22144 4930 22273
rect 5098 22144 5298 22273
rect 5466 22144 5666 22273
rect 5834 22144 6034 22273
rect 6202 22144 6402 22273
rect 6570 22144 6770 22273
rect 6938 22144 7138 22273
rect 7306 22144 7506 22273
rect 7674 22144 7874 22273
rect 8042 22144 8242 22273
rect 8410 22144 8610 22273
rect 8778 22144 8978 22273
rect 9146 22144 9346 22273
rect 9514 22144 9714 22273
rect 9882 22144 10082 22273
rect 10250 22144 10450 22273
rect 10618 22144 10818 22273
rect 10986 22144 11186 22273
rect 11354 22144 11554 22273
rect 11722 22144 11922 22273
rect 12090 22144 12290 22273
rect 12458 22144 12658 22273
rect 12826 22144 13026 22273
rect 13194 22144 13394 22273
rect 13562 22144 13762 22273
rect 13930 22144 14130 22273
rect 14298 22144 14498 22273
rect 14666 22144 14866 22273
rect 15034 22144 15234 22273
rect 15402 22144 15602 22273
rect 15770 22144 15970 22273
rect 16138 22144 16338 22273
rect 16506 22144 16706 22273
rect 16874 22144 17074 22273
rect 17242 22144 17442 22273
rect 17610 22144 17810 22273
rect 17978 22144 18178 22273
rect 18346 22144 18546 22273
rect 18714 22144 18914 22273
rect 19082 22144 19282 22273
rect 19450 22144 19650 22273
rect 19818 22144 20018 22273
rect 20186 22144 20386 22273
rect 20554 22144 20754 22273
rect 20922 22144 21122 22273
rect 21290 22144 21490 22273
rect 21658 22144 21858 22273
rect 22026 22144 22226 22273
rect 22394 22144 22980 22273
rect 20 856 22980 22144
rect 20 2 1434 856
rect 1602 2 1802 856
rect 1970 2 2170 856
rect 2338 2 2538 856
rect 2706 2 2906 856
rect 3074 2 3274 856
rect 3442 2 3642 856
rect 3810 2 4010 856
rect 4178 2 4378 856
rect 4546 2 4746 856
rect 4914 2 5114 856
rect 5282 2 5482 856
rect 5650 2 5850 856
rect 6018 2 6218 856
rect 6386 2 6586 856
rect 6754 2 6954 856
rect 7122 2 7322 856
rect 7490 2 7690 856
rect 7858 2 8058 856
rect 8226 2 8426 856
rect 8594 2 8794 856
rect 8962 2 9162 856
rect 9330 2 9530 856
rect 9698 2 9898 856
rect 10066 2 10266 856
rect 10434 2 10634 856
rect 10802 2 11002 856
rect 11170 2 11370 856
rect 11538 2 11738 856
rect 11906 2 12106 856
rect 12274 2 12474 856
rect 12642 2 12842 856
rect 13010 2 13210 856
rect 13378 2 13578 856
rect 13746 2 13946 856
rect 14114 2 14314 856
rect 14482 2 14682 856
rect 14850 2 15050 856
rect 15218 2 15418 856
rect 15586 2 15786 856
rect 15954 2 16154 856
rect 16322 2 16522 856
rect 16690 2 16890 856
rect 17058 2 17258 856
rect 17426 2 17626 856
rect 17794 2 17994 856
rect 18162 2 18362 856
rect 18530 2 18730 856
rect 18898 2 19098 856
rect 19266 2 19466 856
rect 19634 2 19834 856
rect 20002 2 20202 856
rect 20370 2 20570 856
rect 20738 2 20938 856
rect 21106 2 21306 856
rect 21474 2 22980 856
<< metal3 >>
rect 0 22176 800 22296
rect 22200 22176 23000 22296
rect 0 21768 800 21888
rect 22200 21768 23000 21888
rect 0 21360 800 21480
rect 22200 21360 23000 21480
rect 0 20952 800 21072
rect 22200 20952 23000 21072
rect 0 20544 800 20664
rect 22200 20544 23000 20664
rect 0 20136 800 20256
rect 22200 20136 23000 20256
rect 0 19728 800 19848
rect 22200 19728 23000 19848
rect 0 19320 800 19440
rect 22200 19320 23000 19440
rect 0 18912 800 19032
rect 22200 18912 23000 19032
rect 0 18504 800 18624
rect 22200 18504 23000 18624
rect 0 18096 800 18216
rect 22200 18096 23000 18216
rect 0 17688 800 17808
rect 22200 17688 23000 17808
rect 0 17280 800 17400
rect 22200 17280 23000 17400
rect 0 16872 800 16992
rect 22200 16872 23000 16992
rect 0 16464 800 16584
rect 22200 16464 23000 16584
rect 0 16056 800 16176
rect 22200 16056 23000 16176
rect 0 15648 800 15768
rect 22200 15648 23000 15768
rect 0 15240 800 15360
rect 22200 15240 23000 15360
rect 0 14832 800 14952
rect 22200 14832 23000 14952
rect 0 14424 800 14544
rect 22200 14424 23000 14544
rect 0 14016 800 14136
rect 22200 14016 23000 14136
rect 0 13608 800 13728
rect 22200 13608 23000 13728
rect 0 13200 800 13320
rect 22200 13200 23000 13320
rect 0 12792 800 12912
rect 22200 12792 23000 12912
rect 0 12384 800 12504
rect 22200 12384 23000 12504
rect 0 11976 800 12096
rect 22200 11976 23000 12096
rect 0 11568 800 11688
rect 22200 11568 23000 11688
rect 0 11160 800 11280
rect 22200 11160 23000 11280
rect 0 10752 800 10872
rect 22200 10752 23000 10872
rect 0 10344 800 10464
rect 22200 10344 23000 10464
rect 0 9936 800 10056
rect 22200 9936 23000 10056
rect 0 9528 800 9648
rect 22200 9528 23000 9648
rect 0 9120 800 9240
rect 22200 9120 23000 9240
rect 0 8712 800 8832
rect 22200 8712 23000 8832
rect 0 8304 800 8424
rect 22200 8304 23000 8424
rect 0 7896 800 8016
rect 22200 7896 23000 8016
rect 0 7488 800 7608
rect 22200 7488 23000 7608
rect 0 7080 800 7200
rect 22200 7080 23000 7200
rect 0 6672 800 6792
rect 22200 6672 23000 6792
rect 0 6264 800 6384
rect 22200 6264 23000 6384
rect 0 5856 800 5976
rect 22200 5856 23000 5976
rect 0 5448 800 5568
rect 22200 5448 23000 5568
rect 0 5040 800 5160
rect 22200 5040 23000 5160
rect 0 4632 800 4752
rect 22200 4632 23000 4752
rect 0 4224 800 4344
rect 22200 4224 23000 4344
rect 0 3816 800 3936
rect 22200 3816 23000 3936
rect 0 3408 800 3528
rect 22200 3408 23000 3528
rect 0 3000 800 3120
rect 22200 3000 23000 3120
rect 0 2592 800 2712
rect 22200 2592 23000 2712
rect 0 2184 800 2304
rect 22200 2184 23000 2304
rect 0 1776 800 1896
rect 22200 1776 23000 1896
rect 0 1368 800 1488
rect 22200 1368 23000 1488
rect 0 960 800 1080
rect 22200 960 23000 1080
rect 0 552 800 672
rect 22200 552 23000 672
<< obsm3 >>
rect 54 22376 22202 22540
rect 880 22096 22120 22376
rect 54 21968 22202 22096
rect 880 21688 22120 21968
rect 54 21560 22202 21688
rect 880 21280 22120 21560
rect 54 21152 22202 21280
rect 880 20872 22120 21152
rect 54 20744 22202 20872
rect 880 20464 22120 20744
rect 54 20336 22202 20464
rect 880 20056 22120 20336
rect 54 19928 22202 20056
rect 880 19648 22120 19928
rect 54 19520 22202 19648
rect 880 19240 22120 19520
rect 54 19112 22202 19240
rect 880 18832 22120 19112
rect 54 18704 22202 18832
rect 880 18424 22120 18704
rect 54 18296 22202 18424
rect 880 18016 22120 18296
rect 54 17888 22202 18016
rect 880 17608 22120 17888
rect 54 17480 22202 17608
rect 880 17200 22120 17480
rect 54 17072 22202 17200
rect 880 16792 22120 17072
rect 54 16664 22202 16792
rect 880 16384 22120 16664
rect 54 16256 22202 16384
rect 880 15976 22120 16256
rect 54 15848 22202 15976
rect 880 15568 22120 15848
rect 54 15440 22202 15568
rect 880 15160 22120 15440
rect 54 15032 22202 15160
rect 880 14752 22120 15032
rect 54 14624 22202 14752
rect 880 14344 22120 14624
rect 54 14216 22202 14344
rect 880 13936 22120 14216
rect 54 13808 22202 13936
rect 880 13528 22120 13808
rect 54 13400 22202 13528
rect 880 13120 22120 13400
rect 54 12992 22202 13120
rect 880 12712 22120 12992
rect 54 12584 22202 12712
rect 880 12304 22120 12584
rect 54 12176 22202 12304
rect 880 11896 22120 12176
rect 54 11768 22202 11896
rect 880 11488 22120 11768
rect 54 11360 22202 11488
rect 880 11080 22120 11360
rect 54 10952 22202 11080
rect 880 10672 22120 10952
rect 54 10544 22202 10672
rect 880 10264 22120 10544
rect 54 10136 22202 10264
rect 880 9856 22120 10136
rect 54 9728 22202 9856
rect 880 9448 22120 9728
rect 54 9320 22202 9448
rect 880 9040 22120 9320
rect 54 8912 22202 9040
rect 880 8632 22120 8912
rect 54 8504 22202 8632
rect 880 8224 22120 8504
rect 54 8096 22202 8224
rect 880 7816 22120 8096
rect 54 7688 22202 7816
rect 880 7408 22120 7688
rect 54 7280 22202 7408
rect 880 7000 22120 7280
rect 54 6872 22202 7000
rect 880 6592 22120 6872
rect 54 6464 22202 6592
rect 880 6184 22120 6464
rect 54 6056 22202 6184
rect 880 5776 22120 6056
rect 54 5648 22202 5776
rect 880 5368 22120 5648
rect 54 5240 22202 5368
rect 880 4960 22120 5240
rect 54 4832 22202 4960
rect 880 4552 22120 4832
rect 54 4424 22202 4552
rect 880 4144 22120 4424
rect 54 4016 22202 4144
rect 880 3736 22120 4016
rect 54 3608 22202 3736
rect 880 3328 22120 3608
rect 54 3200 22202 3328
rect 880 2920 22120 3200
rect 54 2792 22202 2920
rect 880 2512 22120 2792
rect 54 2384 22202 2512
rect 880 2104 22120 2384
rect 54 1976 22202 2104
rect 880 1696 22120 1976
rect 54 1568 22202 1696
rect 880 1288 22120 1568
rect 54 1160 22202 1288
rect 880 880 22120 1160
rect 54 752 22202 880
rect 880 472 22120 752
rect 54 35 22202 472
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 59 20800 21653 22541
rect 59 2048 3463 20800
rect 3943 2048 6062 20800
rect 6542 2048 8661 20800
rect 9141 2048 11260 20800
rect 11740 2048 13859 20800
rect 14339 2048 16458 20800
rect 16938 2048 19057 20800
rect 19537 2048 21653 20800
rect 59 35 21653 2048
<< labels >>
rlabel metal2 s 18234 22200 18290 23000 6 Test_en_N_out
port 1 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 Test_en_S_in
port 2 nsew signal input
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_42_
port 5 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 bottom_left_grid_pin_43_
port 6 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_44_
port 7 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 bottom_left_grid_pin_45_
port 8 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_46_
port 9 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_47_
port 10 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 bottom_left_grid_pin_48_
port 11 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 bottom_left_grid_pin_49_
port 12 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 ccff_head
port 13 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 ccff_tail
port 14 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 15 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 chanx_left_in[10]
port 16 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[11]
port 17 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[12]
port 18 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[13]
port 19 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 chanx_left_in[14]
port 20 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[15]
port 21 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[16]
port 22 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[17]
port 23 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[18]
port 24 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[19]
port 25 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 chanx_left_in[1]
port 26 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 chanx_left_in[2]
port 27 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 chanx_left_in[3]
port 28 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 chanx_left_in[4]
port 29 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[5]
port 30 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[6]
port 31 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[7]
port 32 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[8]
port 33 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[9]
port 34 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_out[0]
port 35 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[10]
port 36 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[11]
port 37 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[12]
port 38 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[13]
port 39 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 chanx_left_out[14]
port 40 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 chanx_left_out[15]
port 41 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 chanx_left_out[16]
port 42 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 chanx_left_out[17]
port 43 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[18]
port 44 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[19]
port 45 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 chanx_left_out[1]
port 46 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 chanx_left_out[2]
port 47 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[3]
port 48 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[4]
port 49 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[5]
port 50 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[6]
port 51 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 chanx_left_out[7]
port 52 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 chanx_left_out[8]
port 53 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 chanx_left_out[9]
port 54 nsew signal output
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 55 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[10]
port 56 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[11]
port 57 nsew signal input
rlabel metal3 s 22200 8712 23000 8832 6 chanx_right_in[12]
port 58 nsew signal input
rlabel metal3 s 22200 9120 23000 9240 6 chanx_right_in[13]
port 59 nsew signal input
rlabel metal3 s 22200 9528 23000 9648 6 chanx_right_in[14]
port 60 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[15]
port 61 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[16]
port 62 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[17]
port 63 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[18]
port 64 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[19]
port 65 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[1]
port 66 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[2]
port 67 nsew signal input
rlabel metal3 s 22200 5040 23000 5160 6 chanx_right_in[3]
port 68 nsew signal input
rlabel metal3 s 22200 5448 23000 5568 6 chanx_right_in[4]
port 69 nsew signal input
rlabel metal3 s 22200 5856 23000 5976 6 chanx_right_in[5]
port 70 nsew signal input
rlabel metal3 s 22200 6264 23000 6384 6 chanx_right_in[6]
port 71 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[7]
port 72 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[8]
port 73 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[9]
port 74 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_out[0]
port 75 nsew signal output
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[10]
port 76 nsew signal output
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[11]
port 77 nsew signal output
rlabel metal3 s 22200 16872 23000 16992 6 chanx_right_out[12]
port 78 nsew signal output
rlabel metal3 s 22200 17280 23000 17400 6 chanx_right_out[13]
port 79 nsew signal output
rlabel metal3 s 22200 17688 23000 17808 6 chanx_right_out[14]
port 80 nsew signal output
rlabel metal3 s 22200 18096 23000 18216 6 chanx_right_out[15]
port 81 nsew signal output
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[16]
port 82 nsew signal output
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[17]
port 83 nsew signal output
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[18]
port 84 nsew signal output
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[19]
port 85 nsew signal output
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_out[1]
port 86 nsew signal output
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_out[2]
port 87 nsew signal output
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[3]
port 88 nsew signal output
rlabel metal3 s 22200 13608 23000 13728 6 chanx_right_out[4]
port 89 nsew signal output
rlabel metal3 s 22200 14016 23000 14136 6 chanx_right_out[5]
port 90 nsew signal output
rlabel metal3 s 22200 14424 23000 14544 6 chanx_right_out[6]
port 91 nsew signal output
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[7]
port 92 nsew signal output
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[8]
port 93 nsew signal output
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[9]
port 94 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[0]
port 95 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[10]
port 96 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[11]
port 97 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 98 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[13]
port 99 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[14]
port 100 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[15]
port 101 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[16]
port 102 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 103 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[18]
port 104 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[19]
port 105 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[1]
port 106 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[2]
port 107 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[3]
port 108 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[4]
port 109 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[5]
port 110 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[6]
port 111 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[7]
port 112 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[8]
port 113 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[9]
port 114 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[0]
port 115 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_out[10]
port 116 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[11]
port 117 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[12]
port 118 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[13]
port 119 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[14]
port 120 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[15]
port 121 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[16]
port 122 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[17]
port 123 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[18]
port 124 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[19]
port 125 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_out[1]
port 126 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[2]
port 127 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[3]
port 128 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[4]
port 129 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[5]
port 130 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[6]
port 131 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[7]
port 132 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[8]
port 133 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[9]
port 134 nsew signal output
rlabel metal2 s 3514 22200 3570 23000 6 chany_top_in[0]
port 135 nsew signal input
rlabel metal2 s 7194 22200 7250 23000 6 chany_top_in[10]
port 136 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[11]
port 137 nsew signal input
rlabel metal2 s 7930 22200 7986 23000 6 chany_top_in[12]
port 138 nsew signal input
rlabel metal2 s 8298 22200 8354 23000 6 chany_top_in[13]
port 139 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 140 nsew signal input
rlabel metal2 s 9034 22200 9090 23000 6 chany_top_in[15]
port 141 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[16]
port 142 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[17]
port 143 nsew signal input
rlabel metal2 s 10138 22200 10194 23000 6 chany_top_in[18]
port 144 nsew signal input
rlabel metal2 s 10506 22200 10562 23000 6 chany_top_in[19]
port 145 nsew signal input
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[1]
port 146 nsew signal input
rlabel metal2 s 4250 22200 4306 23000 6 chany_top_in[2]
port 147 nsew signal input
rlabel metal2 s 4618 22200 4674 23000 6 chany_top_in[3]
port 148 nsew signal input
rlabel metal2 s 4986 22200 5042 23000 6 chany_top_in[4]
port 149 nsew signal input
rlabel metal2 s 5354 22200 5410 23000 6 chany_top_in[5]
port 150 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[6]
port 151 nsew signal input
rlabel metal2 s 6090 22200 6146 23000 6 chany_top_in[7]
port 152 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[8]
port 153 nsew signal input
rlabel metal2 s 6826 22200 6882 23000 6 chany_top_in[9]
port 154 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_out[0]
port 155 nsew signal output
rlabel metal2 s 14554 22200 14610 23000 6 chany_top_out[10]
port 156 nsew signal output
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[11]
port 157 nsew signal output
rlabel metal2 s 15290 22200 15346 23000 6 chany_top_out[12]
port 158 nsew signal output
rlabel metal2 s 15658 22200 15714 23000 6 chany_top_out[13]
port 159 nsew signal output
rlabel metal2 s 16026 22200 16082 23000 6 chany_top_out[14]
port 160 nsew signal output
rlabel metal2 s 16394 22200 16450 23000 6 chany_top_out[15]
port 161 nsew signal output
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[16]
port 162 nsew signal output
rlabel metal2 s 17130 22200 17186 23000 6 chany_top_out[17]
port 163 nsew signal output
rlabel metal2 s 17498 22200 17554 23000 6 chany_top_out[18]
port 164 nsew signal output
rlabel metal2 s 17866 22200 17922 23000 6 chany_top_out[19]
port 165 nsew signal output
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_out[1]
port 166 nsew signal output
rlabel metal2 s 11610 22200 11666 23000 6 chany_top_out[2]
port 167 nsew signal output
rlabel metal2 s 11978 22200 12034 23000 6 chany_top_out[3]
port 168 nsew signal output
rlabel metal2 s 12346 22200 12402 23000 6 chany_top_out[4]
port 169 nsew signal output
rlabel metal2 s 12714 22200 12770 23000 6 chany_top_out[5]
port 170 nsew signal output
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[6]
port 171 nsew signal output
rlabel metal2 s 13450 22200 13506 23000 6 chany_top_out[7]
port 172 nsew signal output
rlabel metal2 s 13818 22200 13874 23000 6 chany_top_out[8]
port 173 nsew signal output
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[9]
port 174 nsew signal output
rlabel metal3 s 22200 20136 23000 20256 6 clk_1_E_out
port 175 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 clk_1_N_in
port 176 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 clk_1_W_out
port 177 nsew signal output
rlabel metal3 s 22200 20544 23000 20664 6 clk_2_E_out
port 178 nsew signal output
rlabel metal2 s 18970 22200 19026 23000 6 clk_2_N_in
port 179 nsew signal input
rlabel metal2 s 21178 22200 21234 23000 6 clk_2_N_out
port 180 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 clk_2_S_out
port 181 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 clk_2_W_out
port 182 nsew signal output
rlabel metal3 s 22200 20952 23000 21072 6 clk_3_E_out
port 183 nsew signal output
rlabel metal2 s 19338 22200 19394 23000 6 clk_3_N_in
port 184 nsew signal input
rlabel metal2 s 21546 22200 21602 23000 6 clk_3_N_out
port 185 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 clk_3_S_out
port 186 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 clk_3_W_out
port 187 nsew signal output
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_34_
port 188 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_35_
port 189 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 left_bottom_grid_pin_36_
port 190 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 left_bottom_grid_pin_37_
port 191 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_bottom_grid_pin_38_
port 192 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 left_bottom_grid_pin_39_
port 193 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_40_
port 194 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 195 nsew signal input
rlabel metal2 s 19706 22200 19762 23000 6 prog_clk_0_N_in
port 196 nsew signal input
rlabel metal3 s 22200 21360 23000 21480 6 prog_clk_1_E_out
port 197 nsew signal output
rlabel metal2 s 20074 22200 20130 23000 6 prog_clk_1_N_in
port 198 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 prog_clk_1_W_out
port 199 nsew signal output
rlabel metal3 s 22200 21768 23000 21888 6 prog_clk_2_E_out
port 200 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 prog_clk_2_N_in
port 201 nsew signal input
rlabel metal2 s 21914 22200 21970 23000 6 prog_clk_2_N_out
port 202 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 prog_clk_2_S_out
port 203 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 prog_clk_2_W_out
port 204 nsew signal output
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_3_E_out
port 205 nsew signal output
rlabel metal2 s 20810 22200 20866 23000 6 prog_clk_3_N_in
port 206 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_3_N_out
port 207 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 prog_clk_3_S_out
port 208 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 prog_clk_3_W_out
port 209 nsew signal output
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_34_
port 210 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_35_
port 211 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_36_
port 212 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_37_
port 213 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_38_
port 214 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_39_
port 215 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_40_
port 216 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 217 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_42_
port 218 nsew signal input
rlabel metal2 s 938 22200 994 23000 6 top_left_grid_pin_43_
port 219 nsew signal input
rlabel metal2 s 1306 22200 1362 23000 6 top_left_grid_pin_44_
port 220 nsew signal input
rlabel metal2 s 1674 22200 1730 23000 6 top_left_grid_pin_45_
port 221 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 222 nsew signal input
rlabel metal2 s 2410 22200 2466 23000 6 top_left_grid_pin_47_
port 223 nsew signal input
rlabel metal2 s 2778 22200 2834 23000 6 top_left_grid_pin_48_
port 224 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 top_left_grid_pin_49_
port 225 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2663524
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_1__1_/runs/sb_1__1_/results/signoff/sb_1__1_.magic.gds
string GDS_START 79424
<< end >>

