* NGSPICE file created from bottom_left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

.subckt bottom_left_tile VGND VPWR ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23] chanx_right_in[24]
+ chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28] chanx_right_in[29]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21] chanx_right_out[22]
+ chanx_right_out[23] chanx_right_out[24] chanx_right_out[25] chanx_right_out[26]
+ chanx_right_out[27] chanx_right_out[28] chanx_right_out[29] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[20] chany_top_in[21]
+ chany_top_in[22] chany_top_in[23] chany_top_in[24] chany_top_in[25] chany_top_in[26]
+ chany_top_in[27] chany_top_in[28] chany_top_in[29] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[20] chany_top_out[21]
+ chany_top_out[22] chany_top_out[23] chany_top_out[24] chany_top_out[25] chany_top_out[26]
+ chany_top_out[27] chany_top_out[28] chany_top_out[29] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk prog_reset reset right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_0.mux_l1_in_1_ net141 net22 sb_0__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_32.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_131_ sb_0__0_.mux_top_track_0.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input55_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_10.mux_l2_in_0_ net160 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_10.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ sb_0__0_.mux_top_track_34.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mux_right_track_2.mux_l1_in_0_ net64 net53 sb_0__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input18_A chanx_right_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mux_top_track_12.mux_l2_in_0_ net143 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_12.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput75 net75 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput97 net97 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
Xoutput86 net86 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_44.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_44.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l1_in_0_ net70 net67 sb_0__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_130_ sb_0__0_.mux_top_track_2.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chany_top_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ net3 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_44.mux_l2_in_0__153 VGND VGND VPWR VPWR net153 sb_0__0_.mux_top_track_44.mux_l2_in_0__153/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_right_track_10.mux_l1_in_0_ net65 net49 sb_0__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_6 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_12.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput76 net76 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
Xoutput98 net98 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput87 net87 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input30_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_34.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_44.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_12.mux_l1_in_0_ net16 net67 sb_0__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_28.mux_l2_in_0__148 VGND VGND VPWR VPWR net148 sb_0__0_.mux_top_track_28.mux_l2_in_0__148/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_112_ net31 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input60_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput77 net77 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
Xoutput99 net99 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput88 net88 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input23_A chanx_right_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.ccff_head net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_34.mux_l2_in_0_ net133 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_34.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_18.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_18.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_6.mux_l1_in_1__139 VGND VGND VPWR VPWR net139 sb_0__0_.mux_right_track_6.mux_l1_in_1__139/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_6.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_111_ net30 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input53_A chany_top_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput78 net78 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput89 net89 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
XANTENNA_input16_A chanx_right_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_16.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_18.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__075__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_34.mux_l1_in_0_ net66 net36 sb_0__0_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_4.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_30.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_30.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_top_track_12.mux_l2_in_0__143 VGND VGND VPWR VPWR net143 sb_0__0_.mux_top_track_12.mux_l2_in_0__143/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_right_track_46.mux_l2_in_0_ net136 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_110_ net29 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input46_A chany_top_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_right_track_16.mux_l2_in_0__163 VGND VGND VPWR VPWR net163 sb_0__0_.mux_right_track_16.mux_l2_in_0__163/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput79 net79 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mux_top_track_48.mux_l2_in_0_ net155 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_50.mux_l2_in_0_ net156 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_28.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_30.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input39_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mux_right_track_46.mux_l1_in_0_ net64 net59 sb_0__0_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input21_A chanx_right_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_0.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_48.mux_l1_in_0_ net26 net69 sb_0__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input69_A top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_50.mux_l1_in_0_ net25 net70 sb_0__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_34.mux_l2_in_0__133 VGND VGND VPWR VPWR net133 sb_0__0_.mux_right_track_34.mux_l2_in_0__133/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ sb_0__0_.mux_right_track_4.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chany_top_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_44.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_right_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk net1
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input6_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_8.mux_l2_in_0_ net140 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_10.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_6.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_098_ sb_0__0_.mux_right_track_6.out VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_6.mux_l2_in_0_ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input44_A chany_top_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_4.mux_l2_in_0__134 VGND VGND VPWR VPWR net134 sb_0__0_.mux_right_track_4.mux_l2_in_0__134/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_12.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l1_in_1__141 VGND VGND VPWR VPWR net141 sb_0__0_.mux_top_track_0.mux_l1_in_1__141/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_34.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_6.mux_l1_in_1_ net157 net19 sb_0__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_16.mux_l2_in_0_ net163 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_16.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_4.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_8.mux_l1_in_0_ net64 net50 sb_0__0_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ sb_0__0_.mux_right_track_8.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input37_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_10.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_top_track_18.mux_l2_in_0_ net146 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_18.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_30.mux_l2_in_0__149 VGND VGND VPWR VPWR net149 sb_0__0_.mux_top_track_30.mux_l2_in_0__149/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_6.mux_l1_in_0_ net70 net67 sb_0__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_18.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_37_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_2.mux_l2_in_0__147 VGND VGND VPWR VPWR net147 sb_0__0_.mux_top_track_2.mux_l2_in_0__147/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input67_A top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ sb_0__0_.mux_right_track_10.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_0__0_.mux_right_track_16.mux_l1_in_0_ net65 net46 sb_0__0_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_right_track_28.mux_l2_in_0_ net166 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_28.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_079_ sb_0__0_.mux_right_track_44.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_30.mux_l2_in_0_ net167 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_30.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mux_right_track_48.mux_l2_in_0__137 VGND VGND VPWR VPWR net137 sb_0__0_.mux_right_track_48.mux_l2_in_0__137/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mux_top_track_18.mux_l1_in_0_ net12 net70 sb_0__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_16.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_32.mux_l2_in_0_ net150 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_30.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_10.mux_l2_in_0__142 VGND VGND VPWR VPWR net142 sb_0__0_.mux_top_track_10.mux_l2_in_0__142/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_095_ sb_0__0_.mux_right_track_12.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_28.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_28.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_078_ sb_0__0_.mux_right_track_46.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_14.mux_l2_in_0__162 VGND VGND VPWR VPWR net162 sb_0__0_.mux_right_track_14.mux_l2_in_0__162/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_28.mux_l1_in_0_ net63 net39 sb_0__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_30.mux_l1_in_0_ net64 net38 sb_0__0_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_28.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_top_track_32.mux_l1_in_0_ net5 net69 sb_0__0_.mem_top_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_44.mux_l2_in_0_ net153 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_094_ sb_0__0_.mux_right_track_14.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_18.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_28.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_077_ sb_0__0_.mux_right_track_48.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input35_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ sb_0__0_.mux_top_track_4.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_32.mux_l2_in_0__132 VGND VGND VPWR VPWR net132 sb_0__0_.mux_right_track_32.mux_l2_in_0__132/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ sb_0__0_.mux_right_track_16.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input65_A right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_right_track_2.mux_l2_in_0__165 VGND VGND VPWR VPWR net165 sb_0__0_.mux_right_track_2.mux_l2_in_0__165/LO
+ sky130_fd_sc_hd__conb_1
X_076_ sb_0__0_.mux_right_track_50.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_44.mux_l1_in_0_ net28 net67 sb_0__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input28_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_128_ sb_0__0_.mux_top_track_6.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput70 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net70 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk
+ sb_0__0_.mem_right_track_46.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_46.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input10_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input58_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_092_ sb_0__0_.mux_right_track_18.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 chanx_right_in[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_075_ net56 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_127_ sb_0__0_.mux_top_track_8.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_4.mux_l2_in_0_ net134 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_4.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput60 chany_top_in[8] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_14.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_2.mux_l2_in_0_ net147 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_2.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk
+ sb_0__0_.mem_right_track_44.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_46.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_2.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_28.mux_l2_in_0__166 VGND VGND VPWR VPWR net166 sb_0__0_.mux_right_track_28.mux_l2_in_0__166/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_091_ net44 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_right_in[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input70_A top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ net55 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ sb_0__0_.mux_top_track_10.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 chany_top_in[9] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput50 chany_top_in[26] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input33_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_12.mux_l2_in_0_ net161 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_12.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ sb_0__0_.mux_top_track_44.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_12.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_4.mux_l1_in_0_ net65 net52 sb_0__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_14.mux_l2_in_0_ net144 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_14.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ net42 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_right_in[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_2.mux_l1_in_0_ net21 net68 sb_0__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input63_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ net54 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_8.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ sb_0__0_.mux_top_track_12.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput62 prog_reset VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_12
Xsb_0__0_.mux_right_track_46.mux_l2_in_0__136 VGND VGND VPWR VPWR net136 sb_0__0_.mux_right_track_46.mux_l2_in_0__136/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput51 chany_top_in[27] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput40 chany_top_in[17] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input26_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_108_ sb_0__0_.mux_top_track_46.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_12.mux_l1_in_0_ net63 net48 sb_0__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__081__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 chanx_right_in[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_28.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_14.mux_l1_in_0_ net15 net68 sb_0__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_50.mux_l2_in_0__138 VGND VGND VPWR VPWR net138 sb_0__0_.mux_right_track_50.mux_l2_in_0__138/LO
+ sky130_fd_sc_hd__conb_1
X_072_ net43 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_right_track_12.mux_l2_in_0__161 VGND VGND VPWR VPWR net161 sb_0__0_.mux_right_track_12.mux_l2_in_0__161/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_10 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_6.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_32.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_32.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_124_ sb_0__0_.mux_top_track_14.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
Xinput63 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput52 chany_top_in[28] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_right_in[8] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_top_in[18] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_right_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ sb_0__0_.mux_top_track_48.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_right_in[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_18.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input49_A chany_top_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_30.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_32.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ sb_0__0_.mux_top_track_16.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 chanx_right_in[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 chanx_right_in[9] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput64 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chany_top_in[29] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 chany_top_in[19] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_106_ sb_0__0_.mux_top_track_50.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_2.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_right_in[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input61_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__0_.mux_top_track_18.out VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 chany_top_in[2] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput21 chanx_right_in[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 chanx_right_in[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 chany_top_in[0] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 chany_top_in[1] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput65 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ net24 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_48.mux_l2_in_0_ net137 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_50.mux_l2_in_0_ net138 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ net71 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_46.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_50.mem_out\[0\] net62 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfrtp_2
Xsb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_0.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 chanx_right_in[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
X_121_ net11 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input54_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput66 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_8.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xinput33 chany_top_in[10] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput22 chanx_right_in[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_top_in[3] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_right_in[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput44 chany_top_in[20] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ net13 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_14.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input17_A chanx_right_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_44.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input9_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_48.mux_l1_in_0_ net65 net58 sb_0__0_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_50.mux_l1_in_0_ net66 net57 sb_0__0_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_48.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_50.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_right_in[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_0.mux_l2_in_0_ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput121 net121 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
Xoutput110 net110 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
X_120_ net10 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A chany_top_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_0.mux_l1_in_1_ net159 net66 sb_0__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput56 chany_top_in[4] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_6.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xinput67 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput23 chanx_right_in[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_right_in[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_top_in[21] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_top_in[11] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_103_ net2 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_12.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_30.mux_l2_in_0__167 VGND VGND VPWR VPWR net167 sb_0__0_.mux_right_track_30.mux_l2_in_0__167/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 net122 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
Xoutput100 net100 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_0.mux_l1_in_0_ net63 net32 sb_0__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_34.mux_l2_in_0__151 VGND VGND VPWR VPWR net151 sb_0__0_.mux_top_track_34.mux_l2_in_0__151/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 chanx_right_in[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_top_in[5] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput24 chanx_right_in[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_top_in[22] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_top_in[12] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_44.mux_l2_in_0__135 VGND VGND VPWR VPWR net135 sb_0__0_.mux_right_track_44.mux_l2_in_0__135/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ net23 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_10.mux_l2_in_0_ net142 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_10.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_8.mux_l2_in_0_ net158 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_10.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_right_track_0.mux_l1_in_1__159 VGND VGND VPWR VPWR net159 sb_0__0_.mux_right_track_0.mux_l1_in_1__159/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input22_A chanx_right_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_18.mux_l2_in_0__146 VGND VGND VPWR VPWR net146 sb_0__0_.mux_top_track_18.mux_l2_in_0__146/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_10.mux_l2_in_0__160 VGND VGND VPWR VPWR net160 sb_0__0_.mux_right_track_10.mux_l2_in_0__160/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput123 net123 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_32.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 chanx_right_in[3] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 chanx_right_in[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_top_in[13] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput58 chany_top_in[6] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__clkbuf_2
Xinput47 chany_top_in[23] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_18.mux_l2_in_0_ net164 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_18.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_101_ sb_0__0_.mux_right_track_0.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input52_A chany_top_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_top_track_10.mux_l1_in_0_ net17 net69 sb_0__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input15_A chanx_right_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input7_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_8.mux_l1_in_0_ net18 net68 sb_0__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput124 net124 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_30.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xoutput102 net102 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput59 chany_top_in[7] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 chanx_right_in[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_right_in[4] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 chany_top_in[14] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_top_in[24] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_100_ sb_0__0_.mux_right_track_2.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input45_A chany_top_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_8.mux_l2_in_0__158 VGND VGND VPWR VPWR net158 sb_0__0_.mux_top_track_8.mux_l2_in_0__158/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_18.mux_l1_in_0_ net66 net45 sb_0__0_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_32.mux_l2_in_0_ net132 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_32.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_8.mux_l2_in_0__140 VGND VGND VPWR VPWR net140 sb_0__0_.mux_right_track_8.mux_l2_in_0__140/LO
+ sky130_fd_sc_hd__conb_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput103 net103 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mux_top_track_34.mux_l2_in_0_ net151 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput16 chanx_right_in[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 chanx_right_in[5] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 chany_top_in[15] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput49 chany_top_in[25] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input38_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_50.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A chanx_right_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_48.mux_l2_in_0__155 VGND VGND VPWR VPWR net155 sb_0__0_.mux_top_track_48.mux_l2_in_0__155/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_right_track_32.mux_l1_in_0_ net65 net37 sb_0__0_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_input68_A top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_44.mux_l2_in_0_ net135 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput115 net115 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_48.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_48.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput28 chanx_right_in[6] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_right_in[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_top_in[16] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_34.mux_l1_in_0_ net4 net70 sb_0__0_.mem_top_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_089_ net41 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
Xsb_0__0_.mux_top_track_46.mux_l2_in_0_ net154 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A chany_top_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.ccff_head net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_48.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_input13_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_16.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_16.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input5_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput116 net116 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_46.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_48.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_4.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput18 chanx_right_in[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 chanx_right_in[7] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.mux_l1_in_0_ net63 net60 sb_0__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_088_ net40 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_46.mux_l1_in_0_ net27 net68 sb_0__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_14.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_16.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_6.mux_l1_in_1__157 VGND VGND VPWR VPWR net157 sb_0__0_.mux_top_track_6.mux_l1_in_1__157/LO
+ sky130_fd_sc_hd__conb_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput117 net117 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
Xoutput106 net106 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_2.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput19 chanx_right_in[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mux_top_track_32.mux_l2_in_0__150 VGND VGND VPWR VPWR net150 sb_0__0_.mux_top_track_32.mux_l2_in_0__150/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_087_ sb_0__0_.mux_right_track_28.out VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_16.mux_l2_in_0__145 VGND VGND VPWR VPWR net145 sb_0__0_.mux_top_track_16.mux_l2_in_0__145/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_6.mux_l2_in_0_ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_right_track_6.mux_l1_in_1_ net139 net66 sb_0__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input66_A right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_0__0_.mux_top_track_4.mux_l2_in_0_ net152 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_4.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ sb_0__0_.mux_right_track_30.out VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input29_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_34.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_34.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mux_right_track_14.mux_l2_in_0_ net162 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_14.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input11_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xoutput119 net119 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
Xoutput90 net90 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mux_right_track_6.mux_l1_in_0_ net63 net51 sb_0__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input3_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input59_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_16.mux_l2_in_0_ net145 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_16.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_085_ sb_0__0_.mux_right_track_32.out VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
XFILLER_33_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_4.mux_l1_in_0_ net20 net69 sb_0__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk
+ sb_0__0_.mem_right_track_32.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_34.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input41_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
Xoutput80 net80 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
Xoutput91 net91 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mux_right_track_14.mux_l1_in_0_ net64 net47 sb_0__0_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_4.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_084_ sb_0__0_.mux_right_track_34.out VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_10.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_16.mux_l1_in_0_ net14 net69 sb_0__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_28.mux_l2_in_0_ net148 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input34_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ net9 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xsb_0__0_.mux_top_track_30.mux_l2_in_0_ net149 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_46.mux_l2_in_0__154 VGND VGND VPWR VPWR net154 sb_0__0_.mux_top_track_46.mux_l2_in_0__154/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_48.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput81 net81 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_2.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_4.mux_l2_in_0__152 VGND VGND VPWR VPWR net152 sb_0__0_.mux_top_track_4.mux_l2_in_0__152/LO
+ sky130_fd_sc_hd__conb_1
X_083_ net35 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input64_A right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_10.ccff_head
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_50.mux_l2_in_0__156 VGND VGND VPWR VPWR net156 sb_0__0_.mux_top_track_50.mux_l2_in_0__156/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input27_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_118_ net8 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_16.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_28.mux_l1_in_0_ net7 net67 sb_0__0_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__0_.mux_top_track_30.mux_l1_in_0_ net6 net68 sb_0__0_.mem_top_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_46.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xoutput71 net71 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput82 net82 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_082_ net34 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input57_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_1
X_117_ sb_0__0_.mux_top_track_28.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_14.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput94 net94 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
Xoutput72 net72 VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_12
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_081_ net33 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net62 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_14.mux_l2_in_0__144 VGND VGND VPWR VPWR net144 sb_0__0_.mux_top_track_14.mux_l2_in_0__144/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_116_ sb_0__0_.mux_top_track_30.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input32_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_18.mux_l2_in_0__164 VGND VGND VPWR VPWR net164 sb_0__0_.mux_right_track_18.mux_l2_in_0__164/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput84 net84 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
Xoutput73 net73 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
Xoutput95 net95 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_080_ net61 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_2.mux_l2_in_0_ net165 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_2.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_34.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input62_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ sb_0__0_.mux_top_track_32.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l2_in_0_ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net62 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput74 net74 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
Xoutput96 net96 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
Xoutput85 net85 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

