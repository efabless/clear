magic
tech sky130A
magscale 1 2
timestamp 1656943401
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 1104 892 22056 21004
<< metal2 >>
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
<< obsm2 >>
rect 1214 856 22050 21321
rect 1214 734 1986 856
rect 2154 734 2354 856
rect 2522 734 2722 856
rect 2890 734 3090 856
rect 3258 734 3458 856
rect 3626 734 3826 856
rect 3994 734 4194 856
rect 4362 734 4562 856
rect 4730 734 4930 856
rect 5098 734 5298 856
rect 5466 734 5666 856
rect 5834 734 6034 856
rect 6202 734 6402 856
rect 6570 734 6770 856
rect 6938 734 7138 856
rect 7306 734 7506 856
rect 7674 734 7874 856
rect 8042 734 8242 856
rect 8410 734 8610 856
rect 8778 734 8978 856
rect 9146 734 9346 856
rect 9514 734 9714 856
rect 9882 734 10082 856
rect 10250 734 10450 856
rect 10618 734 10818 856
rect 10986 734 11186 856
rect 11354 734 11554 856
rect 11722 734 11922 856
rect 12090 734 12290 856
rect 12458 734 12658 856
rect 12826 734 13026 856
rect 13194 734 13394 856
rect 13562 734 13762 856
rect 13930 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14866 856
rect 15034 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15970 856
rect 16138 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17810 856
rect 17978 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18914 856
rect 19082 734 19282 856
rect 19450 734 19650 856
rect 19818 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20754 856
rect 20922 734 22050 856
<< metal3 >>
rect 0 21224 800 21344
rect 0 20816 800 20936
rect 0 20408 800 20528
rect 0 20000 800 20120
rect 0 19592 800 19712
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18368 800 18488
rect 0 17960 800 18080
rect 0 17552 800 17672
rect 0 17144 800 17264
rect 22200 17144 23000 17264
rect 0 16736 800 16856
rect 0 16328 800 16448
rect 0 15920 800 16040
rect 0 15512 800 15632
rect 0 15104 800 15224
rect 0 14696 800 14816
rect 0 14288 800 14408
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 13064 800 13184
rect 0 12656 800 12776
rect 0 12248 800 12368
rect 0 11840 800 11960
rect 0 11432 800 11552
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 0 10208 800 10328
rect 0 9800 800 9920
rect 0 9392 800 9512
rect 0 8984 800 9104
rect 0 8576 800 8696
rect 0 8168 800 8288
rect 0 7760 800 7880
rect 0 7352 800 7472
rect 0 6944 800 7064
rect 0 6536 800 6656
rect 0 6128 800 6248
rect 0 5720 800 5840
rect 22200 5720 23000 5840
rect 0 5312 800 5432
rect 0 4904 800 5024
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 0 3680 800 3800
rect 0 3272 800 3392
rect 0 2864 800 2984
rect 0 2456 800 2576
rect 0 2048 800 2168
rect 0 1640 800 1760
<< obsm3 >>
rect 880 21144 22200 21317
rect 800 21016 22200 21144
rect 880 20736 22200 21016
rect 800 20608 22200 20736
rect 880 20328 22200 20608
rect 800 20200 22200 20328
rect 880 19920 22200 20200
rect 800 19792 22200 19920
rect 880 19512 22200 19792
rect 800 19384 22200 19512
rect 880 19104 22200 19384
rect 800 18976 22200 19104
rect 880 18696 22200 18976
rect 800 18568 22200 18696
rect 880 18288 22200 18568
rect 800 18160 22200 18288
rect 880 17880 22200 18160
rect 800 17752 22200 17880
rect 880 17472 22200 17752
rect 800 17344 22200 17472
rect 880 17064 22120 17344
rect 800 16936 22200 17064
rect 880 16656 22200 16936
rect 800 16528 22200 16656
rect 880 16248 22200 16528
rect 800 16120 22200 16248
rect 880 15840 22200 16120
rect 800 15712 22200 15840
rect 880 15432 22200 15712
rect 800 15304 22200 15432
rect 880 15024 22200 15304
rect 800 14896 22200 15024
rect 880 14616 22200 14896
rect 800 14488 22200 14616
rect 880 14208 22200 14488
rect 800 14080 22200 14208
rect 880 13800 22200 14080
rect 800 13672 22200 13800
rect 880 13392 22200 13672
rect 800 13264 22200 13392
rect 880 12984 22200 13264
rect 800 12856 22200 12984
rect 880 12576 22200 12856
rect 800 12448 22200 12576
rect 880 12168 22200 12448
rect 800 12040 22200 12168
rect 880 11760 22200 12040
rect 800 11632 22200 11760
rect 880 11352 22200 11632
rect 800 11224 22200 11352
rect 880 10944 22200 11224
rect 800 10816 22200 10944
rect 880 10536 22200 10816
rect 800 10408 22200 10536
rect 880 10128 22200 10408
rect 800 10000 22200 10128
rect 880 9720 22200 10000
rect 800 9592 22200 9720
rect 880 9312 22200 9592
rect 800 9184 22200 9312
rect 880 8904 22200 9184
rect 800 8776 22200 8904
rect 880 8496 22200 8776
rect 800 8368 22200 8496
rect 880 8088 22200 8368
rect 800 7960 22200 8088
rect 880 7680 22200 7960
rect 800 7552 22200 7680
rect 880 7272 22200 7552
rect 800 7144 22200 7272
rect 880 6864 22200 7144
rect 800 6736 22200 6864
rect 880 6456 22200 6736
rect 800 6328 22200 6456
rect 880 6048 22200 6328
rect 800 5920 22200 6048
rect 880 5640 22120 5920
rect 800 5512 22200 5640
rect 880 5232 22200 5512
rect 800 5104 22200 5232
rect 880 4824 22200 5104
rect 800 4696 22200 4824
rect 880 4416 22200 4696
rect 800 4288 22200 4416
rect 880 4008 22200 4288
rect 800 3880 22200 4008
rect 880 3600 22200 3880
rect 800 3472 22200 3600
rect 880 3192 22200 3472
rect 800 3064 22200 3192
rect 880 2784 22200 3064
rect 800 2656 22200 2784
rect 880 2376 22200 2656
rect 800 2248 22200 2376
rect 880 1968 22200 2248
rect 800 1840 22200 1968
rect 880 1667 22200 1840
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 5579 2075 6062 13973
rect 6542 2075 8661 13973
rect 9141 2075 9509 13973
<< labels >>
rlabel metal2 s 20074 0 20130 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 SC_OUT_BOT
port 2 nsew signal output
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_42_
port 5 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_43_
port 6 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_44_
port 7 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 bottom_left_grid_pin_45_
port 8 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 bottom_left_grid_pin_46_
port 9 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 bottom_left_grid_pin_47_
port 10 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 bottom_left_grid_pin_48_
port 11 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 bottom_left_grid_pin_49_
port 12 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 bottom_right_grid_pin_1_
port 13 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 14 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 15 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[0]
port 16 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 17 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 18 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[12]
port 19 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 chanx_left_in[13]
port 20 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 21 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 22 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 chanx_left_in[16]
port 23 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 24 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 25 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[19]
port 26 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[1]
port 27 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[2]
port 28 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[3]
port 29 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 chanx_left_in[4]
port 30 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[5]
port 31 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[6]
port 32 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[7]
port 33 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[8]
port 34 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 35 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_out[0]
port 36 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[10]
port 37 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[11]
port 38 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[12]
port 39 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[13]
port 40 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[14]
port 41 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[15]
port 42 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[16]
port 43 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 chanx_left_out[17]
port 44 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 chanx_left_out[18]
port 45 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 chanx_left_out[19]
port 46 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[1]
port 47 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[2]
port 48 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 chanx_left_out[3]
port 49 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 chanx_left_out[4]
port 50 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[5]
port 51 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[6]
port 52 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[7]
port 53 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[8]
port 54 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[9]
port 55 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[0]
port 56 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[10]
port 57 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[11]
port 58 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[12]
port 59 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[13]
port 60 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 chany_bottom_in[14]
port 61 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[15]
port 62 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[16]
port 63 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[17]
port 64 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[18]
port 65 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_in[19]
port 66 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[1]
port 67 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[2]
port 68 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 chany_bottom_in[3]
port 69 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[4]
port 70 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[5]
port 71 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[6]
port 72 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[7]
port 73 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_in[8]
port 74 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[9]
port 75 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_out[0]
port 76 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[10]
port 77 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[11]
port 78 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 chany_bottom_out[12]
port 79 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[13]
port 80 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[14]
port 81 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[15]
port 82 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[16]
port 83 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[17]
port 84 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[18]
port 85 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[19]
port 86 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[1]
port 87 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[2]
port 88 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_out[3]
port 89 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[4]
port 90 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[5]
port 91 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[6]
port 92 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[7]
port 93 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_out[8]
port 94 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[9]
port 95 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 left_bottom_grid_pin_34_
port 96 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_35_
port 97 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_36_
port 98 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_37_
port 99 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 left_bottom_grid_pin_38_
port 100 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 left_bottom_grid_pin_39_
port 101 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 left_bottom_grid_pin_40_
port 102 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 left_bottom_grid_pin_41_
port 103 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 left_top_grid_pin_1_
port 104 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 prog_clk_0_S_in
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1046956
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_2__2_/runs/sb_2__2_/results/signoff/sb_2__2_.magic.gds
string GDS_START 65026
<< end >>

