magic
tech sky130A
magscale 1 2
timestamp 1656942843
<< viali >>
rect 2145 14569 2179 14603
rect 8769 14569 8803 14603
rect 16405 14569 16439 14603
rect 7389 14365 7423 14399
rect 7656 14365 7690 14399
rect 10333 14365 10367 14399
rect 12653 14365 12687 14399
rect 12909 14365 12943 14399
rect 13093 14365 13127 14399
rect 16313 14365 16347 14399
rect 18061 14365 18095 14399
rect 10066 14297 10100 14331
rect 14749 14297 14783 14331
rect 16046 14297 16080 14331
rect 17816 14297 17850 14331
rect 8953 14229 8987 14263
rect 11529 14229 11563 14263
rect 14933 14229 14967 14263
rect 16681 14229 16715 14263
rect 11529 14025 11563 14059
rect 13001 14025 13035 14059
rect 16681 14025 16715 14059
rect 1593 13957 1627 13991
rect 3065 13957 3099 13991
rect 9496 13957 9530 13991
rect 14718 13957 14752 13991
rect 16221 13957 16255 13991
rect 2145 13889 2179 13923
rect 2697 13889 2731 13923
rect 2789 13889 2823 13923
rect 8870 13889 8904 13923
rect 9137 13889 9171 13923
rect 9229 13889 9263 13923
rect 12642 13889 12676 13923
rect 14114 13889 14148 13923
rect 14381 13889 14415 13923
rect 14473 13889 14507 13923
rect 15945 13889 15979 13923
rect 17794 13889 17828 13923
rect 18153 13889 18187 13923
rect 1869 13821 1903 13855
rect 2421 13821 2455 13855
rect 3433 13821 3467 13855
rect 12909 13821 12943 13855
rect 18061 13821 18095 13855
rect 7757 13685 7791 13719
rect 10609 13685 10643 13719
rect 15853 13685 15887 13719
rect 3893 13481 3927 13515
rect 11713 13413 11747 13447
rect 1593 13345 1627 13379
rect 2973 13345 3007 13379
rect 7389 13345 7423 13379
rect 2145 13277 2179 13311
rect 2697 13277 2731 13311
rect 3065 13277 3099 13311
rect 7656 13277 7690 13311
rect 11621 13277 11655 13311
rect 13093 13277 13127 13311
rect 15485 13277 15519 13311
rect 16957 13277 16991 13311
rect 17049 13277 17083 13311
rect 1869 13209 1903 13243
rect 2421 13209 2455 13243
rect 3157 13209 3191 13243
rect 11354 13209 11388 13243
rect 12826 13209 12860 13243
rect 15218 13209 15252 13243
rect 16690 13209 16724 13243
rect 17294 13209 17328 13243
rect 3525 13141 3559 13175
rect 8769 13141 8803 13175
rect 10241 13141 10275 13175
rect 14105 13141 14139 13175
rect 15577 13141 15611 13175
rect 18429 13141 18463 13175
rect 1593 12937 1627 12971
rect 2421 12937 2455 12971
rect 3249 12937 3283 12971
rect 3709 12937 3743 12971
rect 8125 12937 8159 12971
rect 1961 12869 1995 12903
rect 9238 12869 9272 12903
rect 2053 12801 2087 12835
rect 2513 12801 2547 12835
rect 3341 12801 3375 12835
rect 9505 12801 9539 12835
rect 12642 12801 12676 12835
rect 12909 12801 12943 12835
rect 14114 12801 14148 12835
rect 14381 12801 14415 12835
rect 15586 12801 15620 12835
rect 15853 12801 15887 12835
rect 17794 12801 17828 12835
rect 18061 12801 18095 12835
rect 1869 12733 1903 12767
rect 3525 12733 3559 12767
rect 2697 12665 2731 12699
rect 16681 12665 16715 12699
rect 2881 12597 2915 12631
rect 4077 12597 4111 12631
rect 11529 12597 11563 12631
rect 13001 12597 13035 12631
rect 14473 12597 14507 12631
rect 15945 12597 15979 12631
rect 1777 12393 1811 12427
rect 2605 12393 2639 12427
rect 3801 12393 3835 12427
rect 10241 12393 10275 12427
rect 2421 12257 2455 12291
rect 2973 12257 3007 12291
rect 3157 12257 3191 12291
rect 4353 12257 4387 12291
rect 15577 12257 15611 12291
rect 3249 12189 3283 12223
rect 4169 12189 4203 12223
rect 11621 12189 11655 12223
rect 13369 12189 13403 12223
rect 17049 12189 17083 12223
rect 17141 12189 17175 12223
rect 11376 12121 11410 12155
rect 13102 12121 13136 12155
rect 15332 12121 15366 12155
rect 16793 12121 16827 12155
rect 17386 12121 17420 12155
rect 1685 12053 1719 12087
rect 2145 12053 2179 12087
rect 2237 12053 2271 12087
rect 3617 12053 3651 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 11989 12053 12023 12087
rect 14197 12053 14231 12087
rect 15669 12053 15703 12087
rect 18521 12053 18555 12087
rect 2789 11849 2823 11883
rect 10057 11849 10091 11883
rect 16405 11849 16439 11883
rect 2421 11781 2455 11815
rect 8340 11781 8374 11815
rect 14136 11781 14170 11815
rect 15862 11781 15896 11815
rect 2329 11713 2363 11747
rect 3157 11713 3191 11747
rect 4261 11713 4295 11747
rect 8944 11713 8978 11747
rect 11796 11713 11830 11747
rect 16681 11713 16715 11747
rect 2605 11645 2639 11679
rect 3249 11645 3283 11679
rect 3341 11645 3375 11679
rect 4077 11645 4111 11679
rect 4169 11645 4203 11679
rect 4813 11645 4847 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 11529 11645 11563 11679
rect 14381 11645 14415 11679
rect 16129 11645 16163 11679
rect 17233 11645 17267 11679
rect 7205 11577 7239 11611
rect 14749 11577 14783 11611
rect 1777 11509 1811 11543
rect 1961 11509 1995 11543
rect 3801 11509 3835 11543
rect 4629 11509 4663 11543
rect 4997 11509 5031 11543
rect 11253 11509 11287 11543
rect 12909 11509 12943 11543
rect 13001 11509 13035 11543
rect 2789 11305 2823 11339
rect 2881 11237 2915 11271
rect 4813 11237 4847 11271
rect 8953 11237 8987 11271
rect 13737 11237 13771 11271
rect 14473 11237 14507 11271
rect 2329 11169 2363 11203
rect 2421 11169 2455 11203
rect 3341 11169 3375 11203
rect 3433 11169 3467 11203
rect 4169 11169 4203 11203
rect 4353 11169 4387 11203
rect 5549 11169 5583 11203
rect 2237 11101 2271 11135
rect 4445 11101 4479 11135
rect 5733 11101 5767 11135
rect 10333 11101 10367 11135
rect 10885 11101 10919 11135
rect 12357 11101 12391 11135
rect 15853 11101 15887 11135
rect 17325 11101 17359 11135
rect 3249 11033 3283 11067
rect 3801 11033 3835 11067
rect 5641 11033 5675 11067
rect 6285 11033 6319 11067
rect 10088 11033 10122 11067
rect 11152 11033 11186 11067
rect 12624 11033 12658 11067
rect 15586 11033 15620 11067
rect 17080 11033 17114 11067
rect 1869 10965 1903 10999
rect 6101 10965 6135 10999
rect 12265 10965 12299 10999
rect 15945 10965 15979 10999
rect 2697 10761 2731 10795
rect 3525 10761 3559 10795
rect 4353 10761 4387 10795
rect 6193 10761 6227 10795
rect 6837 10761 6871 10795
rect 9413 10761 9447 10795
rect 3065 10693 3099 10727
rect 3157 10693 3191 10727
rect 4445 10693 4479 10727
rect 8300 10693 8334 10727
rect 2329 10625 2363 10659
rect 3985 10625 4019 10659
rect 5273 10625 5307 10659
rect 5825 10625 5859 10659
rect 6745 10625 6779 10659
rect 11089 10625 11123 10659
rect 11345 10625 11379 10659
rect 13654 10625 13688 10659
rect 15126 10625 15160 10659
rect 15393 10625 15427 10659
rect 2145 10557 2179 10591
rect 2237 10557 2271 10591
rect 2973 10557 3007 10591
rect 3709 10557 3743 10591
rect 3893 10557 3927 10591
rect 5549 10557 5583 10591
rect 5733 10557 5767 10591
rect 6929 10557 6963 10591
rect 8033 10557 8067 10591
rect 13921 10557 13955 10591
rect 1869 10489 1903 10523
rect 6377 10421 6411 10455
rect 9965 10421 9999 10455
rect 12541 10421 12575 10455
rect 14013 10421 14047 10455
rect 17969 10421 18003 10455
rect 18245 10421 18279 10455
rect 18429 10421 18463 10455
rect 2145 10217 2179 10251
rect 3801 10217 3835 10251
rect 4169 10217 4203 10251
rect 13369 10217 13403 10251
rect 17509 10217 17543 10251
rect 14565 10149 14599 10183
rect 18337 10149 18371 10183
rect 2697 10081 2731 10115
rect 2973 10081 3007 10115
rect 4721 10081 4755 10115
rect 5549 10081 5583 10115
rect 6377 10081 6411 10115
rect 17969 10081 18003 10115
rect 18061 10081 18095 10115
rect 3249 10013 3283 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 7656 10013 7690 10047
rect 10149 10013 10183 10047
rect 10416 10013 10450 10047
rect 11989 10013 12023 10047
rect 15945 10013 15979 10047
rect 17417 10013 17451 10047
rect 2053 9945 2087 9979
rect 2605 9945 2639 9979
rect 4077 9945 4111 9979
rect 4537 9945 4571 9979
rect 5641 9945 5675 9979
rect 12234 9945 12268 9979
rect 15678 9945 15712 9979
rect 17150 9945 17184 9979
rect 2513 9877 2547 9911
rect 4629 9877 4663 9911
rect 5733 9877 5767 9911
rect 6101 9877 6135 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 8769 9877 8803 9911
rect 11529 9877 11563 9911
rect 16037 9877 16071 9911
rect 17877 9877 17911 9911
rect 4077 9673 4111 9707
rect 4537 9673 4571 9707
rect 6377 9673 6411 9707
rect 17141 9673 17175 9707
rect 17325 9673 17359 9707
rect 3617 9605 3651 9639
rect 4997 9605 5031 9639
rect 17049 9605 17083 9639
rect 2513 9537 2547 9571
rect 2973 9537 3007 9571
rect 3433 9537 3467 9571
rect 3985 9537 4019 9571
rect 4905 9537 4939 9571
rect 5365 9537 5399 9571
rect 6193 9537 6227 9571
rect 6745 9537 6779 9571
rect 9065 9537 9099 9571
rect 11078 9537 11112 9571
rect 11345 9537 11379 9571
rect 12081 9537 12115 9571
rect 12337 9537 12371 9571
rect 13553 9537 13587 9571
rect 13820 9537 13854 9571
rect 15025 9537 15059 9571
rect 15281 9537 15315 9571
rect 16865 9537 16899 9571
rect 17877 9537 17911 9571
rect 18245 9537 18279 9571
rect 2237 9469 2271 9503
rect 2421 9469 2455 9503
rect 3893 9469 3927 9503
rect 5089 9469 5123 9503
rect 6837 9469 6871 9503
rect 6929 9469 6963 9503
rect 9321 9469 9355 9503
rect 2881 9401 2915 9435
rect 3157 9401 3191 9435
rect 9965 9401 9999 9435
rect 17601 9401 17635 9435
rect 1961 9333 1995 9367
rect 4445 9333 4479 9367
rect 7941 9333 7975 9367
rect 13461 9333 13495 9367
rect 14933 9333 14967 9367
rect 16405 9333 16439 9367
rect 17693 9333 17727 9367
rect 18061 9333 18095 9367
rect 18429 9333 18463 9367
rect 2789 9129 2823 9163
rect 3801 9129 3835 9163
rect 7021 9129 7055 9163
rect 8769 9129 8803 9163
rect 10333 9129 10367 9163
rect 16957 9129 16991 9163
rect 2329 8993 2363 9027
rect 4445 8993 4479 9027
rect 5917 8993 5951 9027
rect 6469 8993 6503 9027
rect 7389 8993 7423 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 13461 8993 13495 9027
rect 14105 8993 14139 9027
rect 2053 8925 2087 8959
rect 4169 8925 4203 8959
rect 6101 8925 6135 8959
rect 6653 8925 6687 8959
rect 7113 8925 7147 8959
rect 8953 8925 8987 8959
rect 11538 8925 11572 8959
rect 14372 8925 14406 8959
rect 15577 8925 15611 8959
rect 17049 8925 17083 8959
rect 4629 8857 4663 8891
rect 5181 8857 5215 8891
rect 5733 8857 5767 8891
rect 7656 8857 7690 8891
rect 9198 8857 9232 8891
rect 12256 8857 12290 8891
rect 15822 8857 15856 8891
rect 17294 8857 17328 8891
rect 1685 8789 1719 8823
rect 2145 8789 2179 8823
rect 2605 8789 2639 8823
rect 3065 8789 3099 8823
rect 4261 8789 4295 8823
rect 5273 8789 5307 8823
rect 5641 8789 5675 8823
rect 6561 8789 6595 8823
rect 10425 8789 10459 8823
rect 13369 8789 13403 8823
rect 15485 8789 15519 8823
rect 18429 8789 18463 8823
rect 1501 8585 1535 8619
rect 2329 8585 2363 8619
rect 2789 8585 2823 8619
rect 3341 8585 3375 8619
rect 4445 8585 4479 8619
rect 5181 8585 5215 8619
rect 6101 8585 6135 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7941 8585 7975 8619
rect 12725 8585 12759 8619
rect 15945 8585 15979 8619
rect 16957 8585 16991 8619
rect 17509 8585 17543 8619
rect 3525 8517 3559 8551
rect 3985 8517 4019 8551
rect 4537 8517 4571 8551
rect 9628 8517 9662 8551
rect 13860 8517 13894 8551
rect 1961 8449 1995 8483
rect 2881 8449 2915 8483
rect 4077 8449 4111 8483
rect 5089 8449 5123 8483
rect 7021 8449 7055 8483
rect 9873 8449 9907 8483
rect 9965 8449 9999 8483
rect 10232 8449 10266 8483
rect 11897 8449 11931 8483
rect 14105 8449 14139 8483
rect 14565 8449 14599 8483
rect 14832 8449 14866 8483
rect 16773 8449 16807 8483
rect 17969 8449 18003 8483
rect 1777 8381 1811 8415
rect 1869 8381 1903 8415
rect 2973 8381 3007 8415
rect 3801 8381 3835 8415
rect 5273 8381 5307 8415
rect 6929 8381 6963 8415
rect 8033 8381 8067 8415
rect 8125 8381 8159 8415
rect 11989 8381 12023 8415
rect 12081 8381 12115 8415
rect 12541 8381 12575 8415
rect 16405 8381 16439 8415
rect 17233 8381 17267 8415
rect 17417 8381 17451 8415
rect 18337 8381 18371 8415
rect 4721 8313 4755 8347
rect 5549 8313 5583 8347
rect 5825 8313 5859 8347
rect 5917 8313 5951 8347
rect 6561 8313 6595 8347
rect 7573 8313 7607 8347
rect 8493 8313 8527 8347
rect 11529 8313 11563 8347
rect 14473 8313 14507 8347
rect 16037 8313 16071 8347
rect 18153 8313 18187 8347
rect 2421 8245 2455 8279
rect 6469 8245 6503 8279
rect 11345 8245 11379 8279
rect 14289 8245 14323 8279
rect 16221 8245 16255 8279
rect 17877 8245 17911 8279
rect 3617 8041 3651 8075
rect 4721 8041 4755 8075
rect 8769 8041 8803 8075
rect 8953 8041 8987 8075
rect 11713 8041 11747 8075
rect 12541 8041 12575 8075
rect 13921 8041 13955 8075
rect 18337 8041 18371 8075
rect 4261 7973 4295 8007
rect 10793 7973 10827 8007
rect 13645 7973 13679 8007
rect 2053 7905 2087 7939
rect 2145 7905 2179 7939
rect 2881 7905 2915 7939
rect 4353 7905 4387 7939
rect 5365 7905 5399 7939
rect 5733 7905 5767 7939
rect 6561 7905 6595 7939
rect 7849 7905 7883 7939
rect 8217 7905 8251 7939
rect 11345 7905 11379 7939
rect 12357 7905 12391 7939
rect 13001 7905 13035 7939
rect 13185 7905 13219 7939
rect 14197 7905 14231 7939
rect 17049 7905 17083 7939
rect 17969 7905 18003 7939
rect 1777 7837 1811 7871
rect 4629 7837 4663 7871
rect 5089 7837 5123 7871
rect 10333 7837 10367 7871
rect 12909 7837 12943 7871
rect 14473 7837 14507 7871
rect 16405 7837 16439 7871
rect 16957 7837 16991 7871
rect 18153 7837 18187 7871
rect 3065 7769 3099 7803
rect 3893 7769 3927 7803
rect 6745 7769 6779 7803
rect 8401 7769 8435 7803
rect 10066 7769 10100 7803
rect 10701 7769 10735 7803
rect 11161 7769 11195 7803
rect 11253 7769 11287 7803
rect 12173 7769 12207 7803
rect 14381 7769 14415 7803
rect 16138 7769 16172 7803
rect 16865 7769 16899 7803
rect 1593 7701 1627 7735
rect 2237 7701 2271 7735
rect 2605 7701 2639 7735
rect 2973 7701 3007 7735
rect 3433 7701 3467 7735
rect 4077 7701 4111 7735
rect 5181 7701 5215 7735
rect 5825 7701 5859 7735
rect 5917 7701 5951 7735
rect 6285 7701 6319 7735
rect 6653 7701 6687 7735
rect 7113 7701 7147 7735
rect 7205 7701 7239 7735
rect 7573 7701 7607 7735
rect 7665 7701 7699 7735
rect 8309 7701 8343 7735
rect 12081 7701 12115 7735
rect 13369 7701 13403 7735
rect 14841 7701 14875 7735
rect 15025 7701 15059 7735
rect 16497 7701 16531 7735
rect 17325 7701 17359 7735
rect 17693 7701 17727 7735
rect 17785 7701 17819 7735
rect 1777 7497 1811 7531
rect 2237 7497 2271 7531
rect 2881 7497 2915 7531
rect 3341 7497 3375 7531
rect 4905 7497 4939 7531
rect 5365 7497 5399 7531
rect 6193 7497 6227 7531
rect 6561 7497 6595 7531
rect 7757 7497 7791 7531
rect 8125 7497 8159 7531
rect 8953 7497 8987 7531
rect 10241 7497 10275 7531
rect 10977 7497 11011 7531
rect 11345 7497 11379 7531
rect 11897 7497 11931 7531
rect 13093 7497 13127 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 14749 7497 14783 7531
rect 15669 7497 15703 7531
rect 17509 7497 17543 7531
rect 17969 7497 18003 7531
rect 1869 7429 1903 7463
rect 7297 7429 7331 7463
rect 12633 7429 12667 7463
rect 14013 7429 14047 7463
rect 18429 7429 18463 7463
rect 2605 7361 2639 7395
rect 3249 7361 3283 7395
rect 4169 7361 4203 7395
rect 4997 7361 5031 7395
rect 5825 7361 5859 7395
rect 7389 7361 7423 7395
rect 8493 7361 8527 7395
rect 8585 7361 8619 7395
rect 9321 7361 9355 7395
rect 10149 7361 10183 7395
rect 11989 7361 12023 7395
rect 13001 7361 13035 7395
rect 15577 7361 15611 7395
rect 16221 7361 16255 7395
rect 17049 7361 17083 7395
rect 17877 7361 17911 7395
rect 1685 7293 1719 7327
rect 3525 7293 3559 7327
rect 3893 7293 3927 7327
rect 4077 7293 4111 7327
rect 4813 7293 4847 7327
rect 5641 7293 5675 7327
rect 5733 7293 5767 7327
rect 7113 7293 7147 7327
rect 8033 7293 8067 7327
rect 8769 7293 8803 7327
rect 9413 7293 9447 7327
rect 9597 7293 9631 7327
rect 10333 7293 10367 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 12081 7293 12115 7327
rect 12909 7293 12943 7327
rect 14105 7293 14139 7327
rect 14841 7293 14875 7327
rect 15025 7293 15059 7327
rect 15853 7293 15887 7327
rect 17141 7293 17175 7327
rect 17233 7293 17267 7327
rect 18153 7293 18187 7327
rect 2421 7225 2455 7259
rect 4537 7225 4571 7259
rect 6929 7225 6963 7259
rect 16405 7225 16439 7259
rect 16681 7225 16715 7259
rect 2789 7157 2823 7191
rect 6653 7157 6687 7191
rect 9781 7157 9815 7191
rect 11529 7157 11563 7191
rect 12449 7157 12483 7191
rect 13553 7157 13587 7191
rect 14381 7157 14415 7191
rect 15209 7157 15243 7191
rect 16037 7157 16071 7191
rect 1501 6953 1535 6987
rect 4905 6953 4939 6987
rect 7941 6953 7975 6987
rect 9321 6953 9355 6987
rect 11437 6953 11471 6987
rect 16681 6953 16715 6987
rect 17509 6953 17543 6987
rect 9505 6885 9539 6919
rect 11161 6885 11195 6919
rect 1777 6817 1811 6851
rect 3065 6817 3099 6851
rect 4537 6817 4571 6851
rect 4721 6817 4755 6851
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 7573 6817 7607 6851
rect 7757 6817 7791 6851
rect 8401 6817 8435 6851
rect 8585 6817 8619 6851
rect 9965 6817 9999 6851
rect 10149 6817 10183 6851
rect 10977 6817 11011 6851
rect 11989 6817 12023 6851
rect 12817 6817 12851 6851
rect 13737 6817 13771 6851
rect 14289 6817 14323 6851
rect 14473 6817 14507 6851
rect 15669 6817 15703 6851
rect 16405 6817 16439 6851
rect 17233 6817 17267 6851
rect 18061 6817 18095 6851
rect 2697 6749 2731 6783
rect 3249 6749 3283 6783
rect 6009 6749 6043 6783
rect 6377 6749 6411 6783
rect 8309 6749 8343 6783
rect 9873 6749 9907 6783
rect 11805 6749 11839 6783
rect 12633 6749 12667 6783
rect 13461 6749 13495 6783
rect 14565 6749 14599 6783
rect 16221 6749 16255 6783
rect 4445 6681 4479 6715
rect 7021 6681 7055 6715
rect 7481 6681 7515 6715
rect 10793 6681 10827 6715
rect 17877 6681 17911 6715
rect 1869 6613 1903 6647
rect 1961 6613 1995 6647
rect 2329 6613 2363 6647
rect 2513 6613 2547 6647
rect 3157 6613 3191 6647
rect 3617 6613 3651 6647
rect 3985 6613 4019 6647
rect 4077 6613 4111 6647
rect 5273 6613 5307 6647
rect 5825 6613 5859 6647
rect 6193 6613 6227 6647
rect 6745 6613 6779 6647
rect 7113 6613 7147 6647
rect 8953 6613 8987 6647
rect 9229 6613 9263 6647
rect 10333 6613 10367 6647
rect 10701 6613 10735 6647
rect 11897 6613 11931 6647
rect 12265 6613 12299 6647
rect 12725 6613 12759 6647
rect 13093 6613 13127 6647
rect 13553 6613 13587 6647
rect 14933 6613 14967 6647
rect 15025 6613 15059 6647
rect 15393 6613 15427 6647
rect 15485 6613 15519 6647
rect 15853 6613 15887 6647
rect 16313 6613 16347 6647
rect 17049 6613 17083 6647
rect 17141 6613 17175 6647
rect 17969 6613 18003 6647
rect 18337 6613 18371 6647
rect 1685 6409 1719 6443
rect 1961 6409 1995 6443
rect 2421 6409 2455 6443
rect 3433 6409 3467 6443
rect 3801 6409 3835 6443
rect 4169 6409 4203 6443
rect 4261 6409 4295 6443
rect 4629 6409 4663 6443
rect 5089 6409 5123 6443
rect 5825 6409 5859 6443
rect 7665 6409 7699 6443
rect 8125 6409 8159 6443
rect 9137 6409 9171 6443
rect 9689 6409 9723 6443
rect 13553 6409 13587 6443
rect 14013 6409 14047 6443
rect 14473 6409 14507 6443
rect 15209 6409 15243 6443
rect 15301 6409 15335 6443
rect 15669 6409 15703 6443
rect 16037 6409 16071 6443
rect 17509 6409 17543 6443
rect 17877 6409 17911 6443
rect 17969 6409 18003 6443
rect 3157 6341 3191 6375
rect 8769 6341 8803 6375
rect 11345 6341 11379 6375
rect 14381 6341 14415 6375
rect 16957 6341 16991 6375
rect 1501 6273 1535 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 3065 6273 3099 6307
rect 3709 6273 3743 6307
rect 4997 6273 5031 6307
rect 6745 6273 6779 6307
rect 8677 6273 8711 6307
rect 10517 6273 10551 6307
rect 11069 6273 11103 6307
rect 11897 6273 11931 6307
rect 12725 6273 12759 6307
rect 17049 6273 17083 6307
rect 2605 6205 2639 6239
rect 4445 6205 4479 6239
rect 5181 6205 5215 6239
rect 5917 6205 5951 6239
rect 6009 6205 6043 6239
rect 6469 6205 6503 6239
rect 6653 6205 6687 6239
rect 7757 6205 7791 6239
rect 7941 6205 7975 6239
rect 8861 6205 8895 6239
rect 9505 6205 9539 6239
rect 9597 6205 9631 6239
rect 10609 6205 10643 6239
rect 10793 6205 10827 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 12817 6205 12851 6239
rect 13001 6205 13035 6239
rect 13369 6205 13403 6239
rect 13461 6205 13495 6239
rect 14657 6205 14691 6239
rect 15393 6205 15427 6239
rect 16129 6205 16163 6239
rect 16221 6205 16255 6239
rect 16773 6205 16807 6239
rect 18153 6205 18187 6239
rect 2881 6137 2915 6171
rect 7297 6137 7331 6171
rect 10057 6137 10091 6171
rect 11529 6137 11563 6171
rect 13921 6137 13955 6171
rect 17417 6137 17451 6171
rect 5457 6069 5491 6103
rect 7113 6069 7147 6103
rect 8309 6069 8343 6103
rect 10149 6069 10183 6103
rect 12357 6069 12391 6103
rect 14841 6069 14875 6103
rect 18337 6069 18371 6103
rect 1593 5865 1627 5899
rect 1869 5865 1903 5899
rect 2697 5865 2731 5899
rect 3065 5865 3099 5899
rect 3341 5865 3375 5899
rect 3893 5865 3927 5899
rect 4537 5865 4571 5899
rect 5917 5865 5951 5899
rect 9965 5865 9999 5899
rect 12081 5865 12115 5899
rect 13829 5865 13863 5899
rect 14105 5865 14139 5899
rect 15209 5865 15243 5899
rect 16037 5865 16071 5899
rect 18061 5865 18095 5899
rect 18429 5865 18463 5899
rect 3433 5797 3467 5831
rect 4353 5797 4387 5831
rect 4905 5797 4939 5831
rect 16865 5797 16899 5831
rect 17693 5797 17727 5831
rect 2513 5729 2547 5763
rect 4997 5729 5031 5763
rect 5365 5729 5399 5763
rect 5457 5729 5491 5763
rect 6561 5729 6595 5763
rect 7113 5729 7147 5763
rect 7297 5729 7331 5763
rect 7941 5729 7975 5763
rect 8585 5729 8619 5763
rect 8953 5729 8987 5763
rect 9413 5729 9447 5763
rect 10333 5729 10367 5763
rect 11529 5729 11563 5763
rect 12541 5729 12575 5763
rect 12725 5729 12759 5763
rect 13553 5729 13587 5763
rect 14749 5729 14783 5763
rect 15761 5729 15795 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 17417 5729 17451 5763
rect 1777 5661 1811 5695
rect 5549 5661 5583 5695
rect 6377 5661 6411 5695
rect 6929 5661 6963 5695
rect 11897 5661 11931 5695
rect 13277 5661 13311 5695
rect 17325 5661 17359 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 2329 5593 2363 5627
rect 6469 5593 6503 5627
rect 8401 5593 8435 5627
rect 11345 5593 11379 5627
rect 14473 5593 14507 5627
rect 15117 5593 15151 5627
rect 15577 5593 15611 5627
rect 2237 5525 2271 5559
rect 2973 5525 3007 5559
rect 4721 5525 4755 5559
rect 6009 5525 6043 5559
rect 7389 5525 7423 5559
rect 7757 5525 7791 5559
rect 8033 5525 8067 5559
rect 8493 5525 8527 5559
rect 9505 5525 9539 5559
rect 9597 5525 9631 5559
rect 10425 5525 10459 5559
rect 10517 5525 10551 5559
rect 10885 5525 10919 5559
rect 10977 5525 11011 5559
rect 11437 5525 11471 5559
rect 12449 5525 12483 5559
rect 12909 5525 12943 5559
rect 13369 5525 13403 5559
rect 14565 5525 14599 5559
rect 15669 5525 15703 5559
rect 16405 5525 16439 5559
rect 17233 5525 17267 5559
rect 1501 5321 1535 5355
rect 1869 5321 1903 5355
rect 4077 5321 4111 5355
rect 4997 5321 5031 5355
rect 5825 5321 5859 5355
rect 6193 5321 6227 5355
rect 6929 5321 6963 5355
rect 7389 5321 7423 5355
rect 7849 5321 7883 5355
rect 8217 5321 8251 5355
rect 9505 5321 9539 5355
rect 10057 5321 10091 5355
rect 10885 5321 10919 5355
rect 11253 5321 11287 5355
rect 13369 5321 13403 5355
rect 15301 5321 15335 5355
rect 16313 5321 16347 5355
rect 17509 5321 17543 5355
rect 18429 5321 18463 5355
rect 1685 5253 1719 5287
rect 2881 5253 2915 5287
rect 3341 5253 3375 5287
rect 5273 5253 5307 5287
rect 6469 5253 6503 5287
rect 6745 5253 6779 5287
rect 9137 5253 9171 5287
rect 10793 5253 10827 5287
rect 11989 5253 12023 5287
rect 13461 5253 13495 5287
rect 17049 5253 17083 5287
rect 2053 5185 2087 5219
rect 2421 5185 2455 5219
rect 2789 5185 2823 5219
rect 4261 5185 4295 5219
rect 7297 5185 7331 5219
rect 8309 5185 8343 5219
rect 9965 5185 9999 5219
rect 11713 5185 11747 5219
rect 12541 5185 12575 5219
rect 14197 5185 14231 5219
rect 14749 5185 14783 5219
rect 15117 5185 15151 5219
rect 15853 5185 15887 5219
rect 17785 5185 17819 5219
rect 3433 5117 3467 5151
rect 5549 5117 5583 5151
rect 5733 5117 5767 5151
rect 7113 5117 7147 5151
rect 8401 5117 8435 5151
rect 8953 5117 8987 5151
rect 9045 5117 9079 5151
rect 10149 5117 10183 5151
rect 10701 5117 10735 5151
rect 12633 5117 12667 5151
rect 12817 5117 12851 5151
rect 13645 5117 13679 5151
rect 14289 5117 14323 5151
rect 14473 5117 14507 5151
rect 15577 5117 15611 5151
rect 15761 5117 15795 5151
rect 17141 5117 17175 5151
rect 17325 5117 17359 5151
rect 18061 5117 18095 5151
rect 2605 5049 2639 5083
rect 4445 5049 4479 5083
rect 7757 5049 7791 5083
rect 12173 5049 12207 5083
rect 13001 5049 13035 5083
rect 13829 5049 13863 5083
rect 14933 5049 14967 5083
rect 2237 4981 2271 5015
rect 3065 4981 3099 5015
rect 9597 4981 9631 5015
rect 11621 4981 11655 5015
rect 16221 4981 16255 5015
rect 16681 4981 16715 5015
rect 2329 4777 2363 4811
rect 2973 4777 3007 4811
rect 5641 4777 5675 4811
rect 8769 4777 8803 4811
rect 9873 4777 9907 4811
rect 11897 4777 11931 4811
rect 12449 4777 12483 4811
rect 12725 4777 12759 4811
rect 13553 4777 13587 4811
rect 17693 4777 17727 4811
rect 18429 4777 18463 4811
rect 6561 4709 6595 4743
rect 15761 4709 15795 4743
rect 16589 4709 16623 4743
rect 18061 4709 18095 4743
rect 3157 4641 3191 4675
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 9597 4641 9631 4675
rect 10333 4641 10367 4675
rect 10517 4641 10551 4675
rect 11161 4641 11195 4675
rect 11253 4641 11287 4675
rect 12633 4641 12667 4675
rect 13185 4641 13219 4675
rect 13369 4641 13403 4675
rect 14657 4641 14691 4675
rect 15025 4641 15059 4675
rect 15209 4641 15243 4675
rect 16313 4641 16347 4675
rect 17233 4641 17267 4675
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 2789 4573 2823 4607
rect 4997 4573 5031 4607
rect 7941 4573 7975 4607
rect 9505 4573 9539 4607
rect 10241 4573 10275 4607
rect 11069 4573 11103 4607
rect 12081 4573 12115 4607
rect 13829 4573 13863 4607
rect 16129 4573 16163 4607
rect 17509 4573 17543 4607
rect 17877 4573 17911 4607
rect 18245 4573 18279 4607
rect 2053 4505 2087 4539
rect 5273 4505 5307 4539
rect 7849 4505 7883 4539
rect 8309 4505 8343 4539
rect 13093 4505 13127 4539
rect 14473 4505 14507 4539
rect 15301 4505 15335 4539
rect 16221 4505 16255 4539
rect 16957 4505 16991 4539
rect 1501 4437 1535 4471
rect 2605 4437 2639 4471
rect 6009 4437 6043 4471
rect 6653 4437 6687 4471
rect 7021 4437 7055 4471
rect 7113 4437 7147 4471
rect 7481 4437 7515 4471
rect 9045 4437 9079 4471
rect 9413 4437 9447 4471
rect 10701 4437 10735 4471
rect 11621 4437 11655 4471
rect 12265 4437 12299 4471
rect 14105 4437 14139 4471
rect 14565 4437 14599 4471
rect 15669 4437 15703 4471
rect 17049 4437 17083 4471
rect 6377 4233 6411 4267
rect 6653 4233 6687 4267
rect 7021 4233 7055 4267
rect 7389 4233 7423 4267
rect 7481 4233 7515 4267
rect 8309 4233 8343 4267
rect 8769 4233 8803 4267
rect 9321 4233 9355 4267
rect 9413 4233 9447 4267
rect 9873 4233 9907 4267
rect 12081 4233 12115 4267
rect 13737 4233 13771 4267
rect 14105 4233 14139 4267
rect 14473 4233 14507 4267
rect 15209 4233 15243 4267
rect 15945 4233 15979 4267
rect 17325 4233 17359 4267
rect 5549 4165 5583 4199
rect 6929 4165 6963 4199
rect 8677 4165 8711 4199
rect 10057 4165 10091 4199
rect 12909 4165 12943 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 2973 4097 3007 4131
rect 3157 4097 3191 4131
rect 6101 4097 6135 4131
rect 11529 4097 11563 4131
rect 13645 4097 13679 4131
rect 15117 4097 15151 4131
rect 16037 4097 16071 4131
rect 16681 4097 16715 4131
rect 17417 4097 17451 4131
rect 17969 4097 18003 4131
rect 7665 4029 7699 4063
rect 7941 4029 7975 4063
rect 9597 4029 9631 4063
rect 11805 4029 11839 4063
rect 12449 4029 12483 4063
rect 12725 4029 12759 4063
rect 12817 4029 12851 4063
rect 13553 4029 13587 4063
rect 14289 4029 14323 4063
rect 15393 4029 15427 4063
rect 16221 4029 16255 4063
rect 16865 4029 16899 4063
rect 17601 4029 17635 4063
rect 1869 3961 1903 3995
rect 2237 3961 2271 3995
rect 2789 3961 2823 3995
rect 8953 3961 8987 3995
rect 10241 3961 10275 3995
rect 13277 3961 13311 3995
rect 14565 3961 14599 3995
rect 15577 3961 15611 3995
rect 18153 3961 18187 3995
rect 8125 3893 8159 3927
rect 10333 3893 10367 3927
rect 10517 3893 10551 3927
rect 14749 3893 14783 3927
rect 16405 3893 16439 3927
rect 18337 3893 18371 3927
rect 2421 3689 2455 3723
rect 4261 3689 4295 3723
rect 8769 3689 8803 3723
rect 9045 3689 9079 3723
rect 9781 3689 9815 3723
rect 10793 3689 10827 3723
rect 13553 3689 13587 3723
rect 14197 3689 14231 3723
rect 14565 3689 14599 3723
rect 14841 3689 14875 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 16589 3689 16623 3723
rect 16957 3689 16991 3723
rect 17325 3689 17359 3723
rect 18245 3689 18279 3723
rect 18521 3689 18555 3723
rect 13645 3621 13679 3655
rect 14933 3621 14967 3655
rect 15485 3621 15519 3655
rect 6929 3553 6963 3587
rect 11253 3553 11287 3587
rect 15945 3553 15979 3587
rect 16129 3553 16163 3587
rect 1501 3485 1535 3519
rect 1869 3485 1903 3519
rect 2237 3485 2271 3519
rect 2605 3485 2639 3519
rect 2973 3485 3007 3519
rect 4077 3485 4111 3519
rect 6653 3485 6687 3519
rect 7573 3485 7607 3519
rect 8125 3485 8159 3519
rect 10977 3485 11011 3519
rect 12909 3485 12943 3519
rect 14289 3485 14323 3519
rect 16773 3485 16807 3519
rect 17141 3485 17175 3519
rect 17509 3485 17543 3519
rect 17785 3485 17819 3519
rect 18061 3485 18095 3519
rect 2697 3417 2731 3451
rect 7849 3417 7883 3451
rect 8401 3417 8435 3451
rect 13185 3417 13219 3451
rect 1685 3349 1719 3383
rect 2053 3349 2087 3383
rect 3893 3349 3927 3383
rect 15209 3349 15243 3383
rect 16405 3349 16439 3383
rect 16221 3145 16255 3179
rect 16773 3145 16807 3179
rect 17325 3145 17359 3179
rect 18245 3145 18279 3179
rect 7849 3077 7883 3111
rect 12265 3077 12299 3111
rect 16405 3077 16439 3111
rect 16957 3077 16991 3111
rect 2053 3009 2087 3043
rect 2145 3009 2179 3043
rect 3801 3009 3835 3043
rect 5825 3009 5859 3043
rect 7021 3009 7055 3043
rect 7573 3009 7607 3043
rect 10885 3009 10919 3043
rect 11989 3009 12023 3043
rect 12541 3009 12575 3043
rect 14749 3009 14783 3043
rect 14841 3009 14875 3043
rect 15393 3009 15427 3043
rect 15945 3009 15979 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 18061 3009 18095 3043
rect 3617 2941 3651 2975
rect 5549 2941 5583 2975
rect 7205 2941 7239 2975
rect 11161 2941 11195 2975
rect 11713 2941 11747 2975
rect 14473 2941 14507 2975
rect 15025 2941 15059 2975
rect 15669 2941 15703 2975
rect 17785 2941 17819 2975
rect 1869 2805 1903 2839
rect 18429 2805 18463 2839
rect 15209 2601 15243 2635
rect 15669 2601 15703 2635
rect 16221 2601 16255 2635
rect 16405 2601 16439 2635
rect 16865 2601 16899 2635
rect 18061 2601 18095 2635
rect 15577 2533 15611 2567
rect 15945 2533 15979 2567
rect 17049 2533 17083 2567
rect 17233 2533 17267 2567
rect 17785 2533 17819 2567
rect 18429 2533 18463 2567
rect 15025 2465 15059 2499
rect 15301 2397 15335 2431
rect 17417 2397 17451 2431
rect 17877 2397 17911 2431
rect 16037 2261 16071 2295
rect 17509 2261 17543 2295
<< metal1 >>
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 10318 15008 10324 15020
rect 9272 14980 10324 15008
rect 9272 14968 9278 14980
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 12618 14940 12624 14952
rect 8628 14912 12624 14940
rect 8628 14900 8634 14912
rect 12618 14900 12624 14912
rect 12676 14940 12682 14952
rect 13078 14940 13084 14952
rect 12676 14912 13084 14940
rect 12676 14900 12682 14912
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 16942 14872 16948 14884
rect 10100 14844 16948 14872
rect 10100 14832 10106 14844
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 11606 14804 11612 14816
rect 6880 14776 11612 14804
rect 6880 14764 6886 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2774 14600 2780 14612
rect 2179 14572 2780 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 8757 14603 8815 14609
rect 8757 14569 8769 14603
rect 8803 14600 8815 14603
rect 10410 14600 10416 14612
rect 8803 14572 10416 14600
rect 8803 14569 8815 14572
rect 8757 14563 8815 14569
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 15930 14600 15936 14612
rect 14332 14572 15936 14600
rect 14332 14560 14338 14572
rect 15930 14560 15936 14572
rect 15988 14600 15994 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 15988 14572 16405 14600
rect 15988 14560 15994 14572
rect 16393 14569 16405 14572
rect 16439 14569 16451 14603
rect 16393 14563 16451 14569
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 15286 14532 15292 14544
rect 12952 14504 15292 14532
rect 12952 14492 12958 14504
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 13814 14464 13820 14476
rect 12820 14436 13820 14464
rect 7374 14396 7380 14408
rect 7335 14368 7380 14396
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 7644 14399 7702 14405
rect 7644 14365 7656 14399
rect 7690 14396 7702 14399
rect 9214 14396 9220 14408
rect 7690 14368 9220 14396
rect 7690 14365 7702 14368
rect 7644 14359 7702 14365
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 9364 14368 10333 14396
rect 9364 14356 9370 14368
rect 10321 14365 10333 14368
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 12641 14399 12699 14405
rect 12641 14365 12653 14399
rect 12687 14396 12699 14399
rect 12820 14396 12848 14436
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 12687 14368 12848 14396
rect 12897 14399 12955 14405
rect 12687 14365 12699 14368
rect 12641 14359 12699 14365
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 12986 14396 12992 14408
rect 12943 14368 12992 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 14826 14396 14832 14408
rect 13136 14368 14832 14396
rect 13136 14356 13142 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 14918 14356 14924 14408
rect 14976 14396 14982 14408
rect 16301 14399 16359 14405
rect 16301 14396 16313 14399
rect 14976 14368 16313 14396
rect 14976 14356 14982 14368
rect 16301 14365 16313 14368
rect 16347 14365 16359 14399
rect 18046 14396 18052 14408
rect 18007 14368 18052 14396
rect 16301 14359 16359 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 8260 14300 9812 14328
rect 8260 14288 8266 14300
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 8846 14260 8852 14272
rect 2372 14232 8852 14260
rect 2372 14220 2378 14232
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 8941 14263 8999 14269
rect 8941 14229 8953 14263
rect 8987 14260 8999 14263
rect 9674 14260 9680 14272
rect 8987 14232 9680 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9784 14260 9812 14300
rect 10042 14288 10048 14340
rect 10100 14337 10106 14340
rect 10100 14328 10112 14337
rect 10502 14328 10508 14340
rect 10100 14300 10508 14328
rect 10100 14291 10112 14300
rect 10100 14288 10106 14291
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 13446 14288 13452 14340
rect 13504 14328 13510 14340
rect 14737 14331 14795 14337
rect 14737 14328 14749 14331
rect 13504 14300 14749 14328
rect 13504 14288 13510 14300
rect 14737 14297 14749 14300
rect 14783 14328 14795 14331
rect 16034 14331 16092 14337
rect 16034 14328 16046 14331
rect 14783 14300 16046 14328
rect 14783 14297 14795 14300
rect 14737 14291 14795 14297
rect 16034 14297 16046 14300
rect 16080 14297 16092 14331
rect 16034 14291 16092 14297
rect 17804 14331 17862 14337
rect 17804 14297 17816 14331
rect 17850 14328 17862 14331
rect 18414 14328 18420 14340
rect 17850 14300 18420 14328
rect 17850 14297 17862 14300
rect 17804 14291 17862 14297
rect 18414 14288 18420 14300
rect 18472 14288 18478 14340
rect 10226 14260 10232 14272
rect 9784 14232 10232 14260
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 11514 14260 11520 14272
rect 11475 14232 11520 14260
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 13964 14232 14933 14260
rect 13964 14220 13970 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 17034 14260 17040 14272
rect 16715 14232 17040 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 9766 14056 9772 14068
rect 3068 14028 9772 14056
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 2958 13988 2964 14000
rect 1627 13960 2964 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 2148 13929 2176 13960
rect 2958 13948 2964 13960
rect 3016 13948 3022 14000
rect 3068 13997 3096 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 10284 14028 11529 14056
rect 10284 14016 10290 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12989 14059 13047 14065
rect 12989 14056 13001 14059
rect 11664 14028 13001 14056
rect 11664 14016 11670 14028
rect 12989 14025 13001 14028
rect 13035 14025 13047 14059
rect 12989 14019 13047 14025
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 14148 14028 14504 14056
rect 14148 14016 14154 14028
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13957 3111 13991
rect 3053 13951 3111 13957
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 9306 13988 9312 14000
rect 7432 13960 9312 13988
rect 7432 13948 7438 13960
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2133 13883 2191 13889
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2406 13852 2412 13864
rect 2367 13824 2412 13852
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2792 13852 2820 13883
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 8478 13920 8484 13932
rect 6236 13892 8484 13920
rect 6236 13880 6242 13892
rect 8478 13880 8484 13892
rect 8536 13880 8542 13932
rect 8846 13880 8852 13932
rect 8904 13929 8910 13932
rect 9140 13929 9168 13960
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 9484 13991 9542 13997
rect 9484 13957 9496 13991
rect 9530 13988 9542 13991
rect 9582 13988 9588 14000
rect 9530 13960 9588 13988
rect 9530 13957 9542 13960
rect 9484 13951 9542 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 12802 13988 12808 14000
rect 10612 13960 12808 13988
rect 8904 13920 8916 13929
rect 9125 13923 9183 13929
rect 8904 13892 8949 13920
rect 8904 13883 8916 13892
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 9171 13892 9229 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 8904 13880 8910 13883
rect 2866 13852 2872 13864
rect 2779 13824 2872 13852
rect 2866 13812 2872 13824
rect 2924 13852 2930 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 2924 13824 3433 13852
rect 2924 13812 2930 13824
rect 3421 13821 3433 13824
rect 3467 13852 3479 13855
rect 3602 13852 3608 13864
rect 3467 13824 3608 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 7745 13719 7803 13725
rect 7745 13685 7757 13719
rect 7791 13716 7803 13719
rect 8386 13716 8392 13728
rect 7791 13688 8392 13716
rect 7791 13685 7803 13688
rect 7745 13679 7803 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 10612 13725 10640 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 12894 13948 12900 14000
rect 12952 13988 12958 14000
rect 14476 13988 14504 14028
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 14884 14028 16681 14056
rect 14884 14016 14890 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 14706 13991 14764 13997
rect 14706 13988 14718 13991
rect 12952 13960 14412 13988
rect 14476 13960 14718 13988
rect 12952 13948 12958 13960
rect 12618 13880 12624 13932
rect 12676 13929 12682 13932
rect 14384 13929 14412 13960
rect 14706 13957 14718 13960
rect 14752 13957 14764 13991
rect 14706 13951 14764 13957
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 16209 13991 16267 13997
rect 15344 13960 16160 13988
rect 15344 13948 15350 13960
rect 12676 13920 12688 13929
rect 14102 13923 14160 13929
rect 14102 13920 14114 13923
rect 12676 13892 12721 13920
rect 13280 13892 14114 13920
rect 12676 13883 12688 13892
rect 12676 13880 12682 13883
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 10597 13719 10655 13725
rect 10597 13716 10609 13719
rect 8536 13688 10609 13716
rect 8536 13676 8542 13688
rect 10597 13685 10609 13688
rect 10643 13685 10655 13719
rect 10597 13679 10655 13685
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 13280 13716 13308 13892
rect 14102 13889 14114 13892
rect 14148 13889 14160 13923
rect 14102 13883 14160 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 14415 13892 14473 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 15930 13920 15936 13932
rect 15891 13892 15936 13920
rect 14461 13883 14519 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16132 13920 16160 13960
rect 16209 13957 16221 13991
rect 16255 13988 16267 13991
rect 17586 13988 17592 14000
rect 16255 13960 17592 13988
rect 16255 13957 16267 13960
rect 16209 13951 16267 13957
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 17782 13923 17840 13929
rect 17782 13920 17794 13923
rect 16132 13892 17794 13920
rect 17782 13889 17794 13892
rect 17828 13920 17840 13923
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17828 13892 18153 13920
rect 17828 13889 17840 13892
rect 17782 13883 17840 13889
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 15838 13716 15844 13728
rect 11940 13688 13308 13716
rect 15799 13688 15844 13716
rect 11940 13676 11946 13688
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 6914 13512 6920 13524
rect 3927 13484 6920 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 1578 13376 1584 13388
rect 1491 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13376 1642 13388
rect 2961 13379 3019 13385
rect 1636 13348 2728 13376
rect 1636 13336 1642 13348
rect 2700 13320 2728 13348
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 3510 13376 3516 13388
rect 3007 13348 3516 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 2130 13308 2136 13320
rect 2091 13280 2136 13308
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3602 13308 3608 13320
rect 3099 13280 3608 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3602 13268 3608 13280
rect 3660 13308 3666 13320
rect 3896 13308 3924 13475
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 9858 13512 9864 13524
rect 8076 13484 9864 13512
rect 8076 13472 8082 13484
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 13170 13512 13176 13524
rect 9968 13484 13176 13512
rect 7374 13376 7380 13388
rect 7335 13348 7380 13376
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 3660 13280 3924 13308
rect 7644 13311 7702 13317
rect 3660 13268 3666 13280
rect 7644 13277 7656 13311
rect 7690 13308 7702 13311
rect 9968 13308 9996 13484
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 15194 13512 15200 13524
rect 13596 13484 15200 13512
rect 13596 13472 13602 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 11698 13444 11704 13456
rect 11659 13416 11704 13444
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 7690 13280 9996 13308
rect 7690 13277 7702 13280
rect 7644 13271 7702 13277
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 11606 13308 11612 13320
rect 10100 13280 11468 13308
rect 11567 13280 11612 13308
rect 10100 13268 10106 13280
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 2406 13240 2412 13252
rect 2367 13212 2412 13240
rect 2406 13200 2412 13212
rect 2464 13200 2470 13252
rect 3145 13243 3203 13249
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 3694 13240 3700 13252
rect 3191 13212 3700 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 3694 13200 3700 13212
rect 3752 13200 3758 13252
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 11342 13243 11400 13249
rect 11342 13240 11354 13243
rect 8168 13212 11354 13240
rect 8168 13200 8174 13212
rect 11342 13209 11354 13212
rect 11388 13209 11400 13243
rect 11440 13240 11468 13280
rect 11606 13268 11612 13280
rect 11664 13308 11670 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 11664 13280 13093 13308
rect 11664 13268 11670 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 14976 13280 15485 13308
rect 14976 13268 14982 13280
rect 15473 13277 15485 13280
rect 15519 13308 15531 13311
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 15519 13280 16957 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 16945 13277 16957 13280
rect 16991 13308 17003 13311
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 16991 13280 17049 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17037 13277 17049 13280
rect 17083 13308 17095 13311
rect 18046 13308 18052 13320
rect 17083 13280 18052 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 12814 13243 12872 13249
rect 12814 13240 12826 13243
rect 11440 13212 12826 13240
rect 11342 13203 11400 13209
rect 12814 13209 12826 13212
rect 12860 13209 12872 13243
rect 12814 13203 12872 13209
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 15206 13243 15264 13249
rect 15206 13240 15218 13243
rect 13412 13212 15218 13240
rect 13412 13200 13418 13212
rect 15206 13209 15218 13212
rect 15252 13209 15264 13243
rect 15206 13203 15264 13209
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 16678 13243 16736 13249
rect 16678 13240 16690 13243
rect 16080 13212 16690 13240
rect 16080 13200 16086 13212
rect 16678 13209 16690 13212
rect 16724 13209 16736 13243
rect 16678 13203 16736 13209
rect 16850 13200 16856 13252
rect 16908 13240 16914 13252
rect 17282 13243 17340 13249
rect 17282 13240 17294 13243
rect 16908 13212 17294 13240
rect 16908 13200 16914 13212
rect 17282 13209 17294 13212
rect 17328 13209 17340 13243
rect 17282 13203 17340 13209
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3292 13144 3525 13172
rect 3292 13132 3298 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 3513 13135 3571 13141
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 9766 13172 9772 13184
rect 8803 13144 9772 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 11238 13172 11244 13184
rect 10275 13144 11244 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 12492 13144 14105 13172
rect 12492 13132 12498 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 15565 13175 15623 13181
rect 15565 13141 15577 13175
rect 15611 13172 15623 13175
rect 15746 13172 15752 13184
rect 15611 13144 15752 13172
rect 15611 13141 15623 13144
rect 15565 13135 15623 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 18196 13144 18429 13172
rect 18196 13132 18202 13144
rect 18417 13141 18429 13144
rect 18463 13141 18475 13175
rect 18417 13135 18475 13141
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2130 12968 2136 12980
rect 1627 12940 2136 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 3050 12968 3056 12980
rect 2455 12940 3056 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3234 12968 3240 12980
rect 3195 12940 3240 12968
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 3694 12968 3700 12980
rect 3655 12940 3700 12968
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 8110 12968 8116 12980
rect 6972 12940 8116 12968
rect 6972 12928 6978 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 17770 12968 17776 12980
rect 8312 12940 17776 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2958 12900 2964 12912
rect 1995 12872 2964 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 8312 12900 8340 12940
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 6420 12872 8340 12900
rect 6420 12860 6426 12872
rect 9214 12860 9220 12912
rect 9272 12909 9278 12912
rect 9272 12900 9284 12909
rect 9272 12872 9317 12900
rect 9272 12863 9284 12872
rect 9272 12860 9278 12863
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 9456 12872 9536 12900
rect 9456 12860 9462 12872
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3786 12832 3792 12844
rect 3375 12804 3792 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 9508 12841 9536 12872
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 14918 12900 14924 12912
rect 11664 12872 14924 12900
rect 11664 12860 11670 12872
rect 9493 12835 9551 12841
rect 6052 12804 9444 12832
rect 6052 12792 6058 12804
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12733 1915 12767
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 1857 12727 1915 12733
rect 2056 12736 3525 12764
rect 1872 12696 1900 12727
rect 2056 12696 2084 12736
rect 3513 12733 3525 12736
rect 3559 12764 3571 12767
rect 8478 12764 8484 12776
rect 3559 12736 8484 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 9416 12764 9444 12804
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11514 12832 11520 12844
rect 11204 12804 11520 12832
rect 11204 12792 11210 12804
rect 11514 12792 11520 12804
rect 11572 12832 11578 12844
rect 12630 12835 12688 12841
rect 12630 12832 12642 12835
rect 11572 12804 12642 12832
rect 11572 12792 11578 12804
rect 12630 12801 12642 12804
rect 12676 12801 12688 12835
rect 12820 12832 12848 12872
rect 12894 12832 12900 12844
rect 12807 12804 12900 12832
rect 12630 12795 12688 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 14384 12841 14412 12872
rect 14918 12860 14924 12872
rect 14976 12900 14982 12912
rect 14976 12872 15884 12900
rect 14976 12860 14982 12872
rect 14102 12835 14160 12841
rect 14102 12832 14114 12835
rect 13372 12804 14114 12832
rect 9416 12736 11652 12764
rect 1872 12668 2084 12696
rect 2685 12699 2743 12705
rect 2685 12665 2697 12699
rect 2731 12696 2743 12699
rect 2774 12696 2780 12708
rect 2731 12668 2780 12696
rect 2731 12665 2743 12668
rect 2685 12659 2743 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 2866 12628 2872 12640
rect 2827 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 4062 12628 4068 12640
rect 4023 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 8352 12600 11529 12628
rect 8352 12588 8358 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11624 12628 11652 12736
rect 13372 12696 13400 12804
rect 14102 12801 14114 12804
rect 14148 12832 14160 12835
rect 14369 12835 14427 12841
rect 14148 12804 14320 12832
rect 14148 12801 14160 12804
rect 14102 12795 14160 12801
rect 14292 12764 14320 12804
rect 14369 12801 14381 12835
rect 14415 12801 14427 12835
rect 15562 12832 15568 12844
rect 15620 12841 15626 12844
rect 15856 12841 15884 12872
rect 15532 12804 15568 12832
rect 14369 12795 14427 12801
rect 15562 12792 15568 12804
rect 15620 12795 15632 12841
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 15620 12792 15626 12795
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 16632 12804 17794 12832
rect 16632 12792 16638 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 17782 12795 17840 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 14292 12736 14596 12764
rect 12912 12668 13400 12696
rect 12912 12628 12940 12668
rect 11624 12600 12940 12628
rect 12989 12631 13047 12637
rect 11517 12591 11575 12597
rect 12989 12597 13001 12631
rect 13035 12628 13047 12631
rect 13078 12628 13084 12640
rect 13035 12600 13084 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13170 12588 13176 12640
rect 13228 12628 13234 12640
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 13228 12600 14473 12628
rect 13228 12588 13234 12600
rect 14461 12597 14473 12600
rect 14507 12597 14519 12631
rect 14568 12628 14596 12736
rect 16669 12699 16727 12705
rect 16669 12665 16681 12699
rect 16715 12696 16727 12699
rect 16942 12696 16948 12708
rect 16715 12668 16948 12696
rect 16715 12665 16727 12668
rect 16669 12659 16727 12665
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 15838 12628 15844 12640
rect 14568 12600 15844 12628
rect 14461 12591 14519 12597
rect 15838 12588 15844 12600
rect 15896 12628 15902 12640
rect 15933 12631 15991 12637
rect 15933 12628 15945 12631
rect 15896 12600 15945 12628
rect 15896 12588 15902 12600
rect 15933 12597 15945 12600
rect 15979 12597 15991 12631
rect 15933 12591 15991 12597
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 2038 12424 2044 12436
rect 1811 12396 2044 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 2593 12427 2651 12433
rect 2593 12424 2605 12427
rect 2556 12396 2605 12424
rect 2556 12384 2562 12396
rect 2593 12393 2605 12396
rect 2639 12393 2651 12427
rect 3418 12424 3424 12436
rect 2593 12387 2651 12393
rect 2746 12396 3424 12424
rect 2746 12356 2774 12396
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 3786 12424 3792 12436
rect 3747 12396 3792 12424
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10318 12424 10324 12436
rect 10275 12396 10324 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 12066 12424 12072 12436
rect 10428 12396 12072 12424
rect 9582 12356 9588 12368
rect 2424 12328 2774 12356
rect 2976 12328 9588 12356
rect 2424 12297 2452 12328
rect 2976 12297 3004 12328
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12257 2467 12291
rect 2409 12251 2467 12257
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 3108 12260 3157 12288
rect 3108 12248 3114 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 3145 12251 3203 12257
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3970 12288 3976 12300
rect 3476 12260 3976 12288
rect 3476 12248 3482 12260
rect 3970 12248 3976 12260
rect 4028 12288 4034 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 4028 12260 4353 12288
rect 4028 12248 4034 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 10428 12288 10456 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 15838 12424 15844 12436
rect 12406 12396 15844 12424
rect 12406 12356 12434 12396
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 18138 12424 18144 12436
rect 16132 12396 18144 12424
rect 11624 12328 12434 12356
rect 11624 12288 11652 12328
rect 15654 12316 15660 12368
rect 15712 12356 15718 12368
rect 16132 12356 16160 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 15712 12328 16160 12356
rect 15712 12316 15718 12328
rect 15565 12291 15623 12297
rect 15565 12288 15577 12291
rect 8168 12260 10456 12288
rect 11532 12260 11652 12288
rect 15488 12260 15577 12288
rect 8168 12248 8174 12260
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2924 12192 3249 12220
rect 2924 12180 2930 12192
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4120 12192 4169 12220
rect 4120 12180 4126 12192
rect 4157 12189 4169 12192
rect 4203 12220 4215 12223
rect 11054 12220 11060 12232
rect 4203 12192 11060 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11532 12220 11560 12260
rect 11164 12192 11560 12220
rect 4798 12152 4804 12164
rect 2148 12124 2912 12152
rect 2148 12093 2176 12124
rect 2884 12096 2912 12124
rect 3620 12124 4804 12152
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 2133 12087 2191 12093
rect 2133 12084 2145 12087
rect 1719 12056 2145 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 2133 12053 2145 12056
rect 2179 12053 2191 12087
rect 2133 12047 2191 12053
rect 2222 12044 2228 12096
rect 2280 12084 2286 12096
rect 2280 12056 2325 12084
rect 2280 12044 2286 12056
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 3620 12093 3648 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 11164 12152 11192 12192
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 11664 12192 13369 12220
rect 11664 12180 11670 12192
rect 13357 12189 13369 12192
rect 13403 12220 13415 12223
rect 15488 12220 15516 12260
rect 15565 12257 15577 12260
rect 15611 12288 15623 12291
rect 15611 12260 15700 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 13403 12192 15516 12220
rect 15672 12220 15700 12260
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 15672 12192 17049 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 17037 12189 17049 12192
rect 17083 12220 17095 12223
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 17083 12192 17141 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 8812 12124 11192 12152
rect 11364 12155 11422 12161
rect 8812 12112 8818 12124
rect 11364 12121 11376 12155
rect 11410 12152 11422 12155
rect 12802 12152 12808 12164
rect 11410 12124 12808 12152
rect 11410 12121 11422 12124
rect 11364 12115 11422 12121
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13090 12155 13148 12161
rect 13090 12152 13102 12155
rect 12952 12124 13102 12152
rect 12952 12112 12958 12124
rect 13090 12121 13102 12124
rect 13136 12121 13148 12155
rect 13090 12115 13148 12121
rect 15320 12155 15378 12161
rect 15320 12121 15332 12155
rect 15366 12152 15378 12155
rect 15746 12152 15752 12164
rect 15366 12124 15752 12152
rect 15366 12121 15378 12124
rect 15320 12115 15378 12121
rect 15746 12112 15752 12124
rect 15804 12112 15810 12164
rect 16781 12155 16839 12161
rect 16781 12121 16793 12155
rect 16827 12152 16839 12155
rect 16827 12124 16896 12152
rect 16827 12121 16839 12124
rect 16781 12115 16839 12121
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 4706 12084 4712 12096
rect 4295 12056 4712 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 11698 12084 11704 12096
rect 5868 12056 11704 12084
rect 5868 12044 5874 12056
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12526 12084 12532 12096
rect 12124 12056 12532 12084
rect 12124 12044 12130 12056
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 14185 12087 14243 12093
rect 14185 12053 14197 12087
rect 14231 12084 14243 12087
rect 14642 12084 14648 12096
rect 14231 12056 14648 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15657 12087 15715 12093
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 16114 12084 16120 12096
rect 15703 12056 16120 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16868 12084 16896 12124
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17374 12155 17432 12161
rect 17374 12152 17386 12155
rect 17000 12124 17386 12152
rect 17000 12112 17006 12124
rect 17374 12121 17386 12124
rect 17420 12121 17432 12155
rect 17374 12115 17432 12121
rect 17034 12084 17040 12096
rect 16868 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 17920 12056 18521 12084
rect 17920 12044 17926 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 2958 11880 2964 11892
rect 2823 11852 2964 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3418 11840 3424 11892
rect 3476 11880 3482 11892
rect 7282 11880 7288 11892
rect 3476 11852 7288 11880
rect 3476 11840 3482 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9640 11852 10057 11880
rect 9640 11840 9646 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 15988 11852 16405 11880
rect 15988 11840 15994 11852
rect 16393 11849 16405 11852
rect 16439 11849 16451 11883
rect 16393 11843 16451 11849
rect 2409 11815 2467 11821
rect 2409 11781 2421 11815
rect 2455 11812 2467 11815
rect 3050 11812 3056 11824
rect 2455 11784 3056 11812
rect 2455 11781 2467 11784
rect 2409 11775 2467 11781
rect 3050 11772 3056 11784
rect 3108 11812 3114 11824
rect 3510 11812 3516 11824
rect 3108 11784 3516 11812
rect 3108 11772 3114 11784
rect 3510 11772 3516 11784
rect 3568 11772 3574 11824
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 8328 11815 8386 11821
rect 8328 11812 8340 11815
rect 3660 11784 8340 11812
rect 3660 11772 3666 11784
rect 8328 11781 8340 11784
rect 8374 11812 8386 11815
rect 11974 11812 11980 11824
rect 8374 11784 11980 11812
rect 8374 11781 8386 11784
rect 8328 11775 8386 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 14124 11815 14182 11821
rect 14124 11781 14136 11815
rect 14170 11812 14182 11815
rect 15654 11812 15660 11824
rect 14170 11784 15660 11812
rect 14170 11781 14182 11784
rect 14124 11775 14182 11781
rect 15654 11772 15660 11784
rect 15712 11772 15718 11824
rect 15850 11815 15908 11821
rect 15850 11781 15862 11815
rect 15896 11812 15908 11815
rect 16114 11812 16120 11824
rect 15896 11784 16120 11812
rect 15896 11781 15908 11784
rect 15850 11775 15908 11781
rect 16114 11772 16120 11784
rect 16172 11772 16178 11824
rect 2317 11747 2375 11753
rect 2317 11744 2329 11747
rect 1780 11716 2329 11744
rect 1780 11552 1808 11716
rect 2317 11713 2329 11716
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2332 11608 2360 11707
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 2740 11716 3157 11744
rect 2740 11704 2746 11716
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3844 11716 4261 11744
rect 3844 11704 3850 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 8018 11744 8024 11756
rect 4249 11707 4307 11713
rect 7208 11716 8024 11744
rect 2590 11676 2596 11688
rect 2551 11648 2596 11676
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 2924 11648 3249 11676
rect 2924 11636 2930 11648
rect 3237 11645 3249 11648
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3878 11676 3884 11688
rect 3375 11648 3884 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4430 11676 4436 11688
rect 4203 11648 4436 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 4430 11636 4436 11648
rect 4488 11676 4494 11688
rect 4801 11679 4859 11685
rect 4801 11676 4813 11679
rect 4488 11648 4813 11676
rect 4488 11636 4494 11648
rect 4801 11645 4813 11648
rect 4847 11676 4859 11679
rect 4890 11676 4896 11688
rect 4847 11648 4896 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6270 11676 6276 11688
rect 6052 11648 6276 11676
rect 6052 11636 6058 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 3418 11608 3424 11620
rect 2332 11580 3424 11608
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 7208 11617 7236 11716
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8938 11753 8944 11756
rect 8932 11744 8944 11753
rect 8536 11716 8944 11744
rect 8536 11704 8542 11716
rect 8932 11707 8944 11716
rect 8938 11704 8944 11707
rect 8996 11704 9002 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11606 11744 11612 11756
rect 11112 11716 11612 11744
rect 11112 11704 11118 11716
rect 11606 11704 11612 11716
rect 11664 11704 11670 11756
rect 11790 11753 11796 11756
rect 11784 11744 11796 11753
rect 11751 11716 11796 11744
rect 11784 11707 11796 11716
rect 11790 11704 11796 11707
rect 11848 11704 11854 11756
rect 13814 11744 13820 11756
rect 12728 11716 13820 11744
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 8662 11676 8668 11688
rect 8619 11648 8668 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 11514 11676 11520 11688
rect 10284 11648 11520 11676
rect 10284 11636 10290 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 3620 11580 7205 11608
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1949 11543 2007 11549
rect 1949 11509 1961 11543
rect 1995 11540 2007 11543
rect 2314 11540 2320 11552
rect 1995 11512 2320 11540
rect 1995 11509 2007 11512
rect 1949 11503 2007 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 3620 11540 3648 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 9646 11580 11560 11608
rect 2556 11512 3648 11540
rect 3789 11543 3847 11549
rect 2556 11500 2562 11512
rect 3789 11509 3801 11543
rect 3835 11540 3847 11543
rect 3878 11540 3884 11552
rect 3835 11512 3884 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4396 11512 4629 11540
rect 4396 11500 4402 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4982 11540 4988 11552
rect 4943 11512 4988 11540
rect 4617 11503 4675 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 9646 11540 9674 11580
rect 11532 11552 11560 11580
rect 5224 11512 9674 11540
rect 5224 11500 5230 11512
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10962 11540 10968 11552
rect 10008 11512 10968 11540
rect 10008 11500 10014 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 11112 11512 11253 11540
rect 11112 11500 11118 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 11514 11500 11520 11552
rect 11572 11500 11578 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12728 11540 12756 11716
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 16408 11744 16436 11843
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15120 11716 16252 11744
rect 16408 11716 16681 11744
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 12894 11540 12900 11552
rect 11756 11512 12756 11540
rect 12855 11512 12900 11540
rect 11756 11500 11762 11512
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 14090 11540 14096 11552
rect 13035 11512 14096 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14384 11540 14412 11639
rect 14737 11611 14795 11617
rect 14737 11577 14749 11611
rect 14783 11608 14795 11611
rect 15120 11608 15148 11716
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16224 11676 16252 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 17126 11676 17132 11688
rect 16224 11648 17132 11676
rect 16117 11639 16175 11645
rect 14783 11580 15148 11608
rect 14783 11577 14795 11580
rect 14737 11571 14795 11577
rect 15838 11540 15844 11552
rect 14384 11512 15844 11540
rect 15838 11500 15844 11512
rect 15896 11540 15902 11552
rect 16132 11540 16160 11639
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 17236 11540 17264 11639
rect 17310 11540 17316 11552
rect 15896 11512 17316 11540
rect 15896 11500 15902 11512
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 3050 11336 3056 11348
rect 2823 11308 3056 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 3786 11296 3792 11348
rect 3844 11336 3850 11348
rect 4982 11336 4988 11348
rect 3844 11308 4988 11336
rect 3844 11296 3850 11308
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 9950 11336 9956 11348
rect 9416 11308 9956 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 2498 11268 2504 11280
rect 1820 11240 2504 11268
rect 1820 11228 1826 11240
rect 2314 11200 2320 11212
rect 2275 11172 2320 11200
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 2424 11209 2452 11240
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 2869 11271 2927 11277
rect 2869 11268 2881 11271
rect 2746 11240 2881 11268
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2746 11132 2774 11240
rect 2869 11237 2881 11240
rect 2915 11237 2927 11271
rect 3878 11268 3884 11280
rect 2869 11231 2927 11237
rect 3344 11240 3884 11268
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3344 11209 3372 11240
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 4522 11268 4528 11280
rect 4172 11240 4528 11268
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 3108 11172 3341 11200
rect 3108 11160 3114 11172
rect 3329 11169 3341 11172
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 3602 11200 3608 11212
rect 3467 11172 3608 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 3436 11132 3464 11163
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 4172 11209 4200 11240
rect 4522 11228 4528 11240
rect 4580 11228 4586 11280
rect 4801 11271 4859 11277
rect 4801 11237 4813 11271
rect 4847 11237 4859 11271
rect 8846 11268 8852 11280
rect 4801 11231 4859 11237
rect 5552 11240 8852 11268
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11169 4215 11203
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4157 11163 4215 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 2271 11104 2774 11132
rect 3160 11104 3464 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2038 11024 2044 11076
rect 2096 11064 2102 11076
rect 2590 11064 2596 11076
rect 2096 11036 2596 11064
rect 2096 11024 2102 11036
rect 2590 11024 2596 11036
rect 2648 11064 2654 11076
rect 3160 11064 3188 11104
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 3568 11104 4445 11132
rect 3568 11092 3574 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4816 11132 4844 11231
rect 5552 11209 5580 11240
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9416 11268 9444 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 11238 11336 11244 11348
rect 10376 11308 11244 11336
rect 10376 11296 10382 11308
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 15930 11336 15936 11348
rect 11572 11308 15936 11336
rect 11572 11296 11578 11308
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 8987 11240 9444 11268
rect 13725 11271 13783 11277
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 13725 11237 13737 11271
rect 13771 11237 13783 11271
rect 13725 11231 13783 11237
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11169 5595 11203
rect 13740 11200 13768 11231
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 14461 11271 14519 11277
rect 14461 11268 14473 11271
rect 13872 11240 14473 11268
rect 13872 11228 13878 11240
rect 14461 11237 14473 11240
rect 14507 11237 14519 11271
rect 14461 11231 14519 11237
rect 13740 11172 14872 11200
rect 5537 11163 5595 11169
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 4816 11104 5733 11132
rect 4433 11095 4491 11101
rect 5721 11101 5733 11104
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 10226 11132 10232 11144
rect 8720 11104 10232 11132
rect 8720 11092 8726 11104
rect 9416 11076 9444 11104
rect 10226 11092 10232 11104
rect 10284 11132 10290 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 10284 11104 10333 11132
rect 10284 11092 10290 11104
rect 10321 11101 10333 11104
rect 10367 11132 10379 11135
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10367 11104 10885 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10873 11101 10885 11104
rect 10919 11132 10931 11135
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 10919 11104 12357 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 12345 11101 12357 11104
rect 12391 11132 12403 11135
rect 12434 11132 12440 11144
rect 12391 11104 12440 11132
rect 12391 11101 12403 11104
rect 12345 11095 12403 11101
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 14844 11132 14872 11172
rect 15838 11132 15844 11144
rect 14844 11104 15700 11132
rect 15799 11104 15844 11132
rect 2648 11036 3188 11064
rect 3237 11067 3295 11073
rect 2648 11024 2654 11036
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 3283 11036 3801 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3789 11027 3847 11033
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 4396 11036 5641 11064
rect 4396 11024 4402 11036
rect 5629 11033 5641 11036
rect 5675 11033 5687 11067
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 5629 11027 5687 11033
rect 5736 11036 6285 11064
rect 5736 11008 5764 11036
rect 6273 11033 6285 11036
rect 6319 11064 6331 11067
rect 6362 11064 6368 11076
rect 6319 11036 6368 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 8478 11024 8484 11076
rect 8536 11064 8542 11076
rect 8754 11064 8760 11076
rect 8536 11036 8760 11064
rect 8536 11024 8542 11036
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 9398 11024 9404 11076
rect 9456 11024 9462 11076
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10076 11067 10134 11073
rect 10076 11064 10088 11067
rect 9824 11036 10088 11064
rect 9824 11024 9830 11036
rect 10076 11033 10088 11036
rect 10122 11064 10134 11067
rect 11140 11067 11198 11073
rect 10122 11036 11100 11064
rect 10122 11033 10134 11036
rect 10076 11027 10134 11033
rect 11072 11008 11100 11036
rect 11140 11033 11152 11067
rect 11186 11064 11198 11067
rect 12612 11067 12670 11073
rect 11186 11036 12572 11064
rect 11186 11033 11198 11036
rect 11140 11027 11198 11033
rect 12544 11008 12572 11036
rect 12612 11033 12624 11067
rect 12658 11064 12670 11067
rect 12710 11064 12716 11076
rect 12658 11036 12716 11064
rect 12658 11033 12670 11036
rect 12612 11027 12670 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15574 11067 15632 11073
rect 15574 11064 15586 11067
rect 15252 11036 15586 11064
rect 15252 11024 15258 11036
rect 15574 11033 15586 11036
rect 15620 11033 15632 11067
rect 15672 11064 15700 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 16850 11064 16856 11076
rect 15672 11036 16856 11064
rect 15574 11027 15632 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 17068 11067 17126 11073
rect 17068 11064 17080 11067
rect 16960 11036 17080 11064
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 5718 10956 5724 11008
rect 5776 10956 5782 11008
rect 6086 10996 6092 11008
rect 6047 10968 6092 10996
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 12250 10996 12256 11008
rect 12211 10968 12256 10996
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 12526 10956 12532 11008
rect 12584 10956 12590 11008
rect 15933 10999 15991 11005
rect 15933 10965 15945 10999
rect 15979 10996 15991 10999
rect 16114 10996 16120 11008
rect 15979 10968 16120 10996
rect 15979 10965 15991 10968
rect 15933 10959 15991 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 16960 10996 16988 11036
rect 17068 11033 17080 11036
rect 17114 11064 17126 11067
rect 17862 11064 17868 11076
rect 17114 11036 17868 11064
rect 17114 11033 17126 11036
rect 17068 11027 17126 11033
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 18782 11024 18788 11076
rect 18840 11064 18846 11076
rect 19150 11064 19156 11076
rect 18840 11036 19156 11064
rect 18840 11024 18846 11036
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 16632 10968 16988 10996
rect 16632 10956 16638 10968
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3510 10792 3516 10804
rect 3471 10764 3516 10792
rect 3510 10752 3516 10764
rect 3568 10752 3574 10804
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 6181 10795 6239 10801
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6227 10764 6837 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9398 10792 9404 10804
rect 8904 10764 9404 10792
rect 8904 10752 8910 10764
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 11882 10792 11888 10804
rect 10152 10764 11888 10792
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 3053 10727 3111 10733
rect 3053 10724 3065 10727
rect 2556 10696 3065 10724
rect 2556 10684 2562 10696
rect 3053 10693 3065 10696
rect 3099 10693 3111 10727
rect 3053 10687 3111 10693
rect 3145 10727 3203 10733
rect 3145 10693 3157 10727
rect 3191 10724 3203 10727
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 3191 10696 4445 10724
rect 3191 10693 3203 10696
rect 3145 10687 3203 10693
rect 4433 10693 4445 10696
rect 4479 10693 4491 10727
rect 4433 10687 4491 10693
rect 4522 10684 4528 10736
rect 4580 10724 4586 10736
rect 8294 10733 8300 10736
rect 8288 10724 8300 10733
rect 4580 10696 8300 10724
rect 4580 10684 4586 10696
rect 8288 10687 8300 10696
rect 8294 10684 8300 10687
rect 8352 10684 8358 10736
rect 2314 10656 2320 10668
rect 2275 10628 2320 10656
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 3602 10656 3608 10668
rect 2746 10628 3608 10656
rect 2130 10588 2136 10600
rect 2091 10560 2136 10588
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2746 10588 2774 10628
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4154 10656 4160 10668
rect 4019 10628 4160 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4304 10628 5273 10656
rect 4304 10616 4310 10628
rect 5261 10625 5273 10628
rect 5307 10656 5319 10659
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5307 10628 5825 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 6638 10656 6644 10668
rect 5859 10628 6644 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7098 10656 7104 10668
rect 6779 10628 7104 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 10152 10656 10180 10764
rect 11882 10752 11888 10764
rect 11940 10792 11946 10804
rect 12250 10792 12256 10804
rect 11940 10764 12256 10792
rect 11940 10752 11946 10764
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 13630 10752 13636 10804
rect 13688 10792 13694 10804
rect 16574 10792 16580 10804
rect 13688 10764 16580 10792
rect 13688 10752 13694 10764
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10870 10724 10876 10736
rect 10284 10696 10876 10724
rect 10284 10684 10290 10696
rect 10870 10684 10876 10696
rect 10928 10724 10934 10736
rect 15838 10724 15844 10736
rect 10928 10696 11376 10724
rect 10928 10684 10934 10696
rect 10502 10656 10508 10668
rect 7300 10628 10180 10656
rect 10336 10628 10508 10656
rect 2271 10560 2774 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2746 10520 2774 10560
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10557 3755 10591
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3697 10551 3755 10557
rect 1903 10492 2774 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2976 10452 3004 10551
rect 3712 10520 3740 10551
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10557 5595 10591
rect 5718 10588 5724 10600
rect 5679 10560 5724 10588
rect 5537 10551 5595 10557
rect 4522 10520 4528 10532
rect 3712 10492 4528 10520
rect 4522 10480 4528 10492
rect 4580 10480 4586 10532
rect 5552 10520 5580 10551
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6288 10560 6929 10588
rect 5902 10520 5908 10532
rect 5552 10492 5908 10520
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 4706 10452 4712 10464
rect 2976 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6288 10452 6316 10560
rect 6917 10557 6929 10560
rect 6963 10588 6975 10591
rect 7300 10588 7328 10628
rect 6963 10560 7328 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7432 10560 8033 10588
rect 7432 10548 7438 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10336 10588 10364 10628
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 11348 10665 11376 10696
rect 13924 10696 15844 10724
rect 11077 10659 11135 10665
rect 11077 10625 11089 10659
rect 11123 10656 11135 10659
rect 11333 10659 11391 10665
rect 11123 10628 11284 10656
rect 11123 10625 11135 10628
rect 11077 10619 11135 10625
rect 10008 10560 10364 10588
rect 11256 10588 11284 10628
rect 11333 10625 11345 10659
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 13642 10659 13700 10665
rect 13642 10656 13654 10659
rect 11572 10628 13654 10656
rect 11572 10616 11578 10628
rect 13642 10625 13654 10628
rect 13688 10625 13700 10659
rect 13642 10619 13700 10625
rect 13924 10600 13952 10696
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 15396 10665 15424 10696
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 15114 10659 15172 10665
rect 15114 10656 15126 10659
rect 14608 10628 15126 10656
rect 14608 10616 14614 10628
rect 15114 10625 15126 10628
rect 15160 10625 15172 10659
rect 15114 10619 15172 10625
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 11422 10588 11428 10600
rect 11256 10560 11428 10588
rect 10008 10548 10014 10560
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 9214 10480 9220 10532
rect 9272 10520 9278 10532
rect 9272 10492 10088 10520
rect 9272 10480 9278 10492
rect 5592 10424 6316 10452
rect 6365 10455 6423 10461
rect 5592 10412 5598 10424
rect 6365 10421 6377 10455
rect 6411 10452 6423 10455
rect 6546 10452 6552 10464
rect 6411 10424 6552 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 9950 10452 9956 10464
rect 9911 10424 9956 10452
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10060 10452 10088 10492
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 10060 10424 12541 10452
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 12529 10415 12587 10421
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14182 10452 14188 10464
rect 14047 10424 14188 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 17957 10455 18015 10461
rect 17957 10452 17969 10455
rect 17552 10424 17969 10452
rect 17552 10412 17558 10424
rect 17957 10421 17969 10424
rect 18003 10421 18015 10455
rect 18230 10452 18236 10464
rect 18191 10424 18236 10452
rect 17957 10415 18015 10421
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 18506 10452 18512 10464
rect 18463 10424 18512 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2222 10248 2228 10260
rect 2179 10220 2228 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 2556 10220 3801 10248
rect 2556 10208 2562 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 3789 10211 3847 10217
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 6196 10220 8340 10248
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 5718 10180 5724 10192
rect 1544 10152 5724 10180
rect 1544 10140 1550 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 2222 10072 2228 10124
rect 2280 10112 2286 10124
rect 2498 10112 2504 10124
rect 2280 10084 2504 10112
rect 2280 10072 2286 10084
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2648 10084 2697 10112
rect 2648 10072 2654 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2685 10075 2743 10081
rect 2958 10072 2964 10084
rect 3016 10112 3022 10124
rect 3970 10112 3976 10124
rect 3016 10084 3976 10112
rect 3016 10072 3022 10084
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 4706 10112 4712 10124
rect 4667 10084 4712 10112
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2608 10044 2636 10072
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2188 10016 2636 10044
rect 2792 10016 3249 10044
rect 2188 10004 2194 10016
rect 1946 9936 1952 9988
rect 2004 9976 2010 9988
rect 2041 9979 2099 9985
rect 2041 9976 2053 9979
rect 2004 9948 2053 9976
rect 2004 9936 2010 9948
rect 2041 9945 2053 9948
rect 2087 9976 2099 9979
rect 2593 9979 2651 9985
rect 2593 9976 2605 9979
rect 2087 9948 2605 9976
rect 2087 9945 2099 9948
rect 2041 9939 2099 9945
rect 2593 9945 2605 9948
rect 2639 9976 2651 9979
rect 2682 9976 2688 9988
rect 2639 9948 2688 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 2498 9908 2504 9920
rect 2411 9880 2504 9908
rect 2498 9868 2504 9880
rect 2556 9908 2562 9920
rect 2792 9908 2820 10016
rect 3237 10013 3249 10016
rect 3283 10044 3295 10047
rect 5166 10044 5172 10056
rect 3283 10016 5172 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 6196 10044 6224 10220
rect 6454 10140 6460 10192
rect 6512 10180 6518 10192
rect 8312 10180 8340 10220
rect 8846 10208 8852 10260
rect 8904 10248 8910 10260
rect 11514 10248 11520 10260
rect 8904 10220 11520 10248
rect 8904 10208 8910 10220
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 13872 10220 17509 10248
rect 13872 10208 13878 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 9122 10180 9128 10192
rect 6512 10152 6960 10180
rect 8312 10152 9128 10180
rect 6512 10140 6518 10152
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 6822 10112 6828 10124
rect 6411 10084 6828 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 6932 10112 6960 10152
rect 9122 10140 9128 10152
rect 9180 10140 9186 10192
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 14550 10180 14556 10192
rect 13780 10152 14556 10180
rect 13780 10140 13786 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 18325 10183 18383 10189
rect 18325 10180 18337 10183
rect 17972 10152 18337 10180
rect 6932 10084 7512 10112
rect 6546 10044 6552 10056
rect 5552 10016 6224 10044
rect 6507 10016 6552 10044
rect 4062 9976 4068 9988
rect 3975 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9976 4126 9988
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 4120 9948 4537 9976
rect 4120 9936 4126 9948
rect 4525 9945 4537 9948
rect 4571 9976 4583 9979
rect 5552 9976 5580 10016
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 7374 10044 7380 10056
rect 7335 10016 7380 10044
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7484 10044 7512 10084
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 17972 10121 18000 10152
rect 18325 10149 18337 10152
rect 18371 10149 18383 10183
rect 18325 10143 18383 10149
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17828 10084 17969 10112
rect 17828 10072 17834 10084
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 7644 10047 7702 10053
rect 7644 10044 7656 10047
rect 7484 10016 7656 10044
rect 7644 10013 7656 10016
rect 7690 10044 7702 10047
rect 8202 10044 8208 10056
rect 7690 10016 8208 10044
rect 7690 10013 7702 10016
rect 7644 10007 7702 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9732 10016 10149 10044
rect 9732 10004 9738 10016
rect 10137 10013 10149 10016
rect 10183 10044 10195 10047
rect 10226 10044 10232 10056
rect 10183 10016 10232 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10410 10053 10416 10056
rect 10404 10007 10416 10053
rect 10468 10044 10474 10056
rect 10468 10016 10504 10044
rect 10410 10004 10416 10007
rect 10468 10004 10474 10016
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 10928 10016 11989 10044
rect 10928 10004 10934 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15896 10016 15945 10044
rect 15896 10004 15902 10016
rect 15933 10013 15945 10016
rect 15979 10044 15991 10047
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 15979 10016 17417 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18064 10044 18092 10075
rect 17920 10016 18092 10044
rect 17920 10004 17926 10016
rect 4571 9948 5580 9976
rect 5629 9979 5687 9985
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 5629 9945 5641 9979
rect 5675 9976 5687 9979
rect 7466 9976 7472 9988
rect 5675 9948 7472 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 10042 9976 10048 9988
rect 8076 9948 10048 9976
rect 8076 9936 8082 9948
rect 10042 9936 10048 9948
rect 10100 9936 10106 9988
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 12222 9979 12280 9985
rect 12222 9976 12234 9979
rect 10744 9948 12234 9976
rect 10744 9936 10750 9948
rect 12222 9945 12234 9948
rect 12268 9945 12280 9979
rect 12222 9939 12280 9945
rect 15654 9936 15660 9988
rect 15712 9985 15718 9988
rect 15712 9976 15724 9985
rect 15712 9948 15757 9976
rect 15712 9939 15724 9948
rect 15712 9936 15718 9939
rect 17126 9936 17132 9988
rect 17184 9985 17190 9988
rect 17184 9976 17196 9985
rect 17184 9948 17229 9976
rect 17184 9939 17196 9948
rect 17184 9936 17190 9939
rect 2556 9880 2820 9908
rect 2556 9868 2562 9880
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 4672 9880 4717 9908
rect 4672 9868 4678 9880
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6089 9911 6147 9917
rect 5776 9880 5821 9908
rect 5776 9868 5782 9880
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6135 9880 6469 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 8202 9908 8208 9920
rect 6963 9880 8208 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 10226 9908 10232 9920
rect 9456 9880 10232 9908
rect 9456 9868 9462 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11882 9908 11888 9920
rect 11563 9880 11888 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 12860 9880 16037 9908
rect 12860 9868 12866 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 17862 9908 17868 9920
rect 17823 9880 17868 9908
rect 16025 9871 16083 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3234 9704 3240 9716
rect 2740 9676 3240 9704
rect 2740 9664 2746 9676
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 4028 9676 4077 9704
rect 4028 9664 4034 9676
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 4065 9667 4123 9673
rect 4525 9707 4583 9713
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 4614 9704 4620 9716
rect 4571 9676 4620 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5776 9676 6377 9704
rect 5776 9664 5782 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 17129 9707 17187 9713
rect 17129 9704 17141 9707
rect 7340 9676 17141 9704
rect 7340 9664 7346 9676
rect 17129 9673 17141 9676
rect 17175 9704 17187 9707
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 17175 9676 17325 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17313 9673 17325 9676
rect 17359 9704 17371 9707
rect 17862 9704 17868 9716
rect 17359 9676 17868 9704
rect 17359 9673 17371 9676
rect 17313 9667 17371 9673
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 3605 9639 3663 9645
rect 3605 9636 3617 9639
rect 3200 9608 3617 9636
rect 3200 9596 3206 9608
rect 3605 9605 3617 9608
rect 3651 9636 3663 9639
rect 4246 9636 4252 9648
rect 3651 9608 4252 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 4246 9596 4252 9608
rect 4304 9636 4310 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4304 9608 4997 9636
rect 4304 9596 4310 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 5258 9596 5264 9648
rect 5316 9636 5322 9648
rect 8386 9636 8392 9648
rect 5316 9608 8392 9636
rect 5316 9596 5322 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 8496 9608 9674 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2682 9568 2688 9580
rect 2547 9540 2688 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2832 9540 2973 9568
rect 2832 9528 2838 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3510 9568 3516 9580
rect 3467 9540 3516 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 3510 9528 3516 9540
rect 3568 9568 3574 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3568 9540 3985 9568
rect 3568 9528 3574 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5166 9568 5172 9580
rect 4939 9540 5172 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5166 9528 5172 9540
rect 5224 9568 5230 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5224 9540 5365 9568
rect 5224 9528 5230 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 6178 9568 6184 9580
rect 6091 9540 6184 9568
rect 5353 9531 5411 9537
rect 6178 9528 6184 9540
rect 6236 9568 6242 9580
rect 6730 9568 6736 9580
rect 6236 9540 6736 9568
rect 6236 9528 6242 9540
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 8018 9568 8024 9580
rect 7432 9540 8024 9568
rect 7432 9528 7438 9540
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8496 9568 8524 9608
rect 8220 9540 8524 9568
rect 9053 9571 9111 9577
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 2225 9503 2283 9509
rect 2225 9500 2237 9503
rect 2188 9472 2237 9500
rect 2188 9460 2194 9472
rect 2225 9469 2237 9472
rect 2271 9469 2283 9503
rect 2225 9463 2283 9469
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5810 9500 5816 9512
rect 5123 9472 5816 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 2424 9432 2452 9463
rect 2866 9432 2872 9444
rect 1964 9404 2452 9432
rect 2827 9404 2872 9432
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 1964 9373 1992 9404
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3694 9432 3700 9444
rect 3191 9404 3700 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 3896 9432 3924 9463
rect 5092 9432 5120 9463
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9500 6975 9503
rect 8110 9500 8116 9512
rect 6963 9472 8116 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 3844 9404 5120 9432
rect 3844 9392 3850 9404
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 6932 9432 6960 9463
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8220 9432 8248 9540
rect 9053 9537 9065 9571
rect 9099 9568 9111 9571
rect 9214 9568 9220 9580
rect 9099 9540 9220 9568
rect 9099 9537 9111 9540
rect 9053 9531 9111 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9646 9568 9674 9608
rect 9766 9596 9772 9648
rect 9824 9636 9830 9648
rect 10226 9636 10232 9648
rect 9824 9608 10232 9636
rect 9824 9596 9830 9608
rect 10226 9596 10232 9608
rect 10284 9636 10290 9648
rect 12434 9636 12440 9648
rect 10284 9608 11284 9636
rect 10284 9596 10290 9608
rect 10686 9568 10692 9580
rect 9646 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9568 10750 9580
rect 11066 9571 11124 9577
rect 11066 9568 11078 9571
rect 10744 9540 11078 9568
rect 10744 9528 10750 9540
rect 11066 9537 11078 9540
rect 11112 9537 11124 9571
rect 11066 9531 11124 9537
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 9674 9500 9680 9512
rect 9355 9472 9680 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 11256 9500 11284 9608
rect 12084 9608 12440 9636
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11790 9568 11796 9580
rect 11379 9540 11796 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11790 9528 11796 9540
rect 11848 9568 11854 9580
rect 12084 9577 12112 9608
rect 12434 9596 12440 9608
rect 12492 9636 12498 9648
rect 13906 9636 13912 9648
rect 12492 9608 13912 9636
rect 12492 9596 12498 9608
rect 13556 9577 13584 9608
rect 13906 9596 13912 9608
rect 13964 9636 13970 9648
rect 15102 9636 15108 9648
rect 13964 9608 15108 9636
rect 13964 9596 13970 9608
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 11848 9540 12081 9568
rect 11848 9528 11854 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 12325 9571 12383 9577
rect 12325 9568 12337 9571
rect 12069 9531 12127 9537
rect 12176 9540 12337 9568
rect 12176 9500 12204 9540
rect 12325 9537 12337 9540
rect 12371 9537 12383 9571
rect 12325 9531 12383 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 13808 9571 13866 9577
rect 13808 9537 13820 9571
rect 13854 9568 13866 9571
rect 14090 9568 14096 9580
rect 13854 9540 14096 9568
rect 13854 9537 13866 9540
rect 13808 9531 13866 9537
rect 14090 9528 14096 9540
rect 14148 9568 14154 9580
rect 14734 9568 14740 9580
rect 14148 9540 14740 9568
rect 14148 9528 14154 9540
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15028 9577 15056 9608
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17402 9636 17408 9648
rect 17083 9608 17408 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15269 9571 15327 9577
rect 15269 9568 15281 9571
rect 15013 9531 15071 9537
rect 15120 9540 15281 9568
rect 15120 9500 15148 9540
rect 15269 9537 15281 9540
rect 15315 9537 15327 9571
rect 15269 9531 15327 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17586 9568 17592 9580
rect 16899 9540 17592 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17736 9540 17877 9568
rect 17736 9528 17742 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 11256 9472 12204 9500
rect 14936 9472 15148 9500
rect 5960 9404 6960 9432
rect 7116 9404 8248 9432
rect 5960 9392 5966 9404
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 1360 9336 1961 9364
rect 1360 9324 1366 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4212 9336 4445 9364
rect 4212 9324 4218 9336
rect 4433 9333 4445 9336
rect 4479 9333 4491 9367
rect 4433 9327 4491 9333
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 7116 9364 7144 9404
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 9953 9435 10011 9441
rect 9953 9432 9965 9435
rect 9824 9404 9965 9432
rect 9824 9392 9830 9404
rect 9953 9401 9965 9404
rect 9999 9432 10011 9435
rect 10134 9432 10140 9444
rect 9999 9404 10140 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 5132 9336 7144 9364
rect 7929 9367 7987 9373
rect 5132 9324 5138 9336
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 8938 9364 8944 9376
rect 7975 9336 8944 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 10042 9364 10048 9376
rect 9088 9336 10048 9364
rect 9088 9324 9094 9336
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14936 9373 14964 9472
rect 17589 9435 17647 9441
rect 17589 9401 17601 9435
rect 17635 9432 17647 9435
rect 18248 9432 18276 9531
rect 18782 9432 18788 9444
rect 17635 9404 18788 9432
rect 17635 9401 17647 9404
rect 17589 9395 17647 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14240 9336 14933 9364
rect 14240 9324 14246 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 15712 9336 16405 9364
rect 15712 9324 15718 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 16393 9327 16451 9333
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 18046 9364 18052 9376
rect 18007 9336 18052 9364
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 18417 9367 18475 9373
rect 18417 9333 18429 9367
rect 18463 9364 18475 9367
rect 18598 9364 18604 9376
rect 18463 9336 18604 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 3789 9163 3847 9169
rect 2832 9132 2877 9160
rect 2832 9120 2838 9132
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 3878 9160 3884 9172
rect 3835 9132 3884 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 5810 9160 5816 9172
rect 3988 9132 5816 9160
rect 2958 9052 2964 9104
rect 3016 9092 3022 9104
rect 3988 9092 4016 9132
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6880 9132 7021 9160
rect 6880 9120 6886 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 8754 9160 8760 9172
rect 7009 9123 7067 9129
rect 7392 9132 8616 9160
rect 8715 9132 8760 9160
rect 3016 9064 4016 9092
rect 3016 9052 3022 9064
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 7392 9092 7420 9132
rect 4120 9064 7420 9092
rect 8588 9092 8616 9132
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 10318 9160 10324 9172
rect 9640 9132 10324 9160
rect 9640 9120 9646 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 13354 9160 13360 9172
rect 10428 9132 13360 9160
rect 8938 9092 8944 9104
rect 8588 9064 8944 9092
rect 4120 9052 4126 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 2406 9024 2412 9036
rect 2363 8996 2412 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4706 9024 4712 9036
rect 4479 8996 4712 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 7006 9024 7012 9036
rect 6503 8996 7012 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1912 8928 2053 8956
rect 1912 8916 1918 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 4154 8956 4160 8968
rect 4115 8928 4160 8956
rect 2041 8919 2099 8925
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 5684 8928 6101 8956
rect 5684 8916 5690 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 6687 8928 7113 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7101 8925 7113 8928
rect 7147 8956 7159 8959
rect 7147 8928 7880 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 2740 8860 3096 8888
rect 2740 8848 2746 8860
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 2133 8823 2191 8829
rect 2133 8789 2145 8823
rect 2179 8820 2191 8823
rect 2314 8820 2320 8832
rect 2179 8792 2320 8820
rect 2179 8789 2191 8792
rect 2133 8783 2191 8789
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8820 2651 8823
rect 2866 8820 2872 8832
rect 2639 8792 2872 8820
rect 2639 8789 2651 8792
rect 2593 8783 2651 8789
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 3068 8829 3096 8860
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4617 8891 4675 8897
rect 4617 8888 4629 8891
rect 4028 8860 4629 8888
rect 4028 8848 4034 8860
rect 4617 8857 4629 8860
rect 4663 8857 4675 8891
rect 5166 8888 5172 8900
rect 5127 8860 5172 8888
rect 4617 8851 4675 8857
rect 5166 8848 5172 8860
rect 5224 8888 5230 8900
rect 5721 8891 5779 8897
rect 5721 8888 5733 8891
rect 5224 8860 5733 8888
rect 5224 8848 5230 8860
rect 5721 8857 5733 8860
rect 5767 8888 5779 8891
rect 6822 8888 6828 8900
rect 5767 8860 6828 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 7644 8891 7702 8897
rect 7644 8888 7656 8891
rect 6972 8860 7656 8888
rect 6972 8848 6978 8860
rect 7644 8857 7656 8860
rect 7690 8857 7702 8891
rect 7852 8888 7880 8928
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8076 8928 8953 8956
rect 8076 8916 8082 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 9674 8956 9680 8968
rect 8987 8928 9680 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 8294 8888 8300 8900
rect 7852 8860 8300 8888
rect 7644 8851 7702 8857
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9186 8891 9244 8897
rect 9186 8888 9198 8891
rect 8536 8860 9198 8888
rect 8536 8848 8542 8860
rect 9186 8857 9198 8860
rect 9232 8857 9244 8891
rect 10428 8888 10456 9132
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 15194 9160 15200 9172
rect 13504 9132 15200 9160
rect 13504 9120 13510 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 9024 11854 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11848 8996 11989 9024
rect 11848 8984 11854 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 13044 8996 13461 9024
rect 13044 8984 13050 8996
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 14090 9024 14096 9036
rect 13964 8996 14096 9024
rect 13964 8984 13970 8996
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11526 8959 11584 8965
rect 11526 8956 11538 8959
rect 11204 8928 11538 8956
rect 11204 8916 11210 8928
rect 11526 8925 11538 8928
rect 11572 8956 11584 8959
rect 11572 8928 11652 8956
rect 11572 8925 11584 8928
rect 11526 8919 11584 8925
rect 11624 8900 11652 8928
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 11940 8928 12434 8956
rect 11940 8916 11946 8928
rect 9186 8851 9244 8857
rect 9646 8860 10456 8888
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3602 8820 3608 8832
rect 3099 8792 3608 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4430 8820 4436 8832
rect 4295 8792 4436 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 4948 8792 5273 8820
rect 4948 8780 4954 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5626 8820 5632 8832
rect 5587 8792 5632 8820
rect 5261 8783 5319 8789
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 5868 8792 6561 8820
rect 5868 8780 5874 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7190 8820 7196 8832
rect 7064 8792 7196 8820
rect 7064 8780 7070 8792
rect 7190 8780 7196 8792
rect 7248 8820 7254 8832
rect 9646 8820 9674 8860
rect 11606 8848 11612 8900
rect 11664 8848 11670 8900
rect 12250 8897 12256 8900
rect 12244 8888 12256 8897
rect 12211 8860 12256 8888
rect 12244 8851 12256 8860
rect 12250 8848 12256 8851
rect 12308 8848 12314 8900
rect 12406 8888 12434 8928
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13998 8956 14004 8968
rect 13412 8928 14004 8956
rect 13412 8916 13418 8928
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14360 8959 14418 8965
rect 14360 8925 14372 8959
rect 14406 8925 14418 8959
rect 14360 8919 14418 8925
rect 12406 8860 13584 8888
rect 7248 8792 9674 8820
rect 7248 8780 7254 8792
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10413 8823 10471 8829
rect 10413 8820 10425 8823
rect 10284 8792 10425 8820
rect 10284 8780 10290 8792
rect 10413 8789 10425 8792
rect 10459 8789 10471 8823
rect 13354 8820 13360 8832
rect 13315 8792 13360 8820
rect 10413 8783 10471 8789
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 13556 8820 13584 8860
rect 14274 8848 14280 8900
rect 14332 8888 14338 8900
rect 14384 8888 14412 8919
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 15160 8928 15577 8956
rect 15160 8916 15166 8928
rect 15565 8925 15577 8928
rect 15611 8956 15623 8959
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 15611 8928 17049 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 15810 8891 15868 8897
rect 15810 8888 15822 8891
rect 14332 8860 14412 8888
rect 14476 8860 15822 8888
rect 14332 8848 14338 8860
rect 14476 8820 14504 8860
rect 15810 8857 15822 8860
rect 15856 8857 15868 8891
rect 17282 8891 17340 8897
rect 17282 8888 17294 8891
rect 15810 8851 15868 8857
rect 15948 8860 17294 8888
rect 13556 8792 14504 8820
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15436 8792 15485 8820
rect 15436 8780 15442 8792
rect 15473 8789 15485 8792
rect 15519 8820 15531 8823
rect 15948 8820 15976 8860
rect 17282 8857 17294 8860
rect 17328 8857 17340 8891
rect 17282 8851 17340 8857
rect 15519 8792 15976 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18414 8820 18420 8832
rect 18012 8792 18420 8820
rect 18012 8780 18018 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2823 8588 3341 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 3329 8585 3341 8588
rect 3375 8616 3387 8619
rect 4154 8616 4160 8628
rect 3375 8588 4160 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 5166 8616 5172 8628
rect 5079 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6089 8619 6147 8625
rect 6089 8616 6101 8619
rect 5868 8588 6101 8616
rect 5868 8576 5874 8588
rect 6089 8585 6101 8588
rect 6135 8585 6147 8619
rect 6089 8579 6147 8585
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 6420 8588 7113 8616
rect 6420 8576 6426 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7515 8588 7941 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 12250 8616 12256 8628
rect 8720 8588 12256 8616
rect 8720 8576 8726 8588
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12710 8616 12716 8628
rect 12623 8588 12716 8616
rect 12710 8576 12716 8588
rect 12768 8616 12774 8628
rect 14550 8616 14556 8628
rect 12768 8588 14556 8616
rect 12768 8576 12774 8588
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16022 8616 16028 8628
rect 15979 8588 16028 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16022 8576 16028 8588
rect 16080 8616 16086 8628
rect 16390 8616 16396 8628
rect 16080 8588 16396 8616
rect 16080 8576 16086 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 3513 8551 3571 8557
rect 3513 8548 3525 8551
rect 1360 8520 3525 8548
rect 1360 8508 1366 8520
rect 3513 8517 3525 8520
rect 3559 8548 3571 8551
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3559 8520 3985 8548
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 3973 8517 3985 8520
rect 4019 8548 4031 8551
rect 4525 8551 4583 8557
rect 4525 8548 4537 8551
rect 4019 8520 4537 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 4525 8517 4537 8520
rect 4571 8548 4583 8551
rect 5184 8548 5212 8576
rect 4571 8520 5212 8548
rect 6656 8520 7420 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2648 8452 2774 8480
rect 2648 8440 2654 8452
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2314 8412 2320 8424
rect 1903 8384 2320 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2746 8344 2774 8452
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 2924 8452 3464 8480
rect 2924 8440 2930 8452
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 2976 8344 3004 8375
rect 2746 8316 3004 8344
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 1820 8248 2421 8276
rect 1820 8236 1826 8248
rect 2409 8245 2421 8248
rect 2455 8245 2467 8279
rect 3436 8276 3464 8452
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3660 8452 4077 8480
rect 3660 8440 3666 8452
rect 4065 8449 4077 8452
rect 4111 8480 4123 8483
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4111 8452 5089 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 3786 8412 3792 8424
rect 3747 8384 3792 8412
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4522 8344 4528 8356
rect 4212 8316 4528 8344
rect 4212 8304 4218 8316
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 4706 8344 4712 8356
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5000 8344 5028 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 6656 8480 6684 8520
rect 5224 8452 6684 8480
rect 5224 8440 5230 8452
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6880 8452 7021 8480
rect 6880 8440 6886 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7392 8480 7420 8520
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 9616 8551 9674 8557
rect 9616 8548 9628 8551
rect 8444 8520 9628 8548
rect 8444 8508 8450 8520
rect 9616 8517 9628 8520
rect 9662 8548 9674 8551
rect 13078 8548 13084 8560
rect 9662 8520 13084 8548
rect 9662 8517 9674 8520
rect 9616 8511 9674 8517
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 13848 8551 13906 8557
rect 13848 8517 13860 8551
rect 13894 8548 13906 8551
rect 14734 8548 14740 8560
rect 13894 8520 14740 8548
rect 13894 8517 13906 8520
rect 13848 8511 13906 8517
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 15010 8508 15016 8560
rect 15068 8508 15074 8560
rect 7392 8452 9812 8480
rect 7009 8443 7067 8449
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 6914 8412 6920 8424
rect 5316 8384 5361 8412
rect 6875 8384 6920 8412
rect 5316 8372 5322 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 9784 8412 9812 8452
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9916 8452 9965 8480
rect 9916 8440 9922 8452
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 10220 8483 10278 8489
rect 10220 8480 10232 8483
rect 9953 8443 10011 8449
rect 10060 8452 10232 8480
rect 10060 8412 10088 8452
rect 10220 8449 10232 8452
rect 10266 8480 10278 8483
rect 10502 8480 10508 8492
rect 10266 8452 10508 8480
rect 10266 8449 10278 8452
rect 10220 8443 10278 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10744 8452 11008 8480
rect 10744 8440 10750 8452
rect 8168 8384 8213 8412
rect 9784 8384 10088 8412
rect 8168 8372 8174 8384
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 5000 8316 5549 8344
rect 5000 8288 5028 8316
rect 5537 8313 5549 8316
rect 5583 8344 5595 8347
rect 5718 8344 5724 8356
rect 5583 8316 5724 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 5902 8344 5908 8356
rect 5859 8316 5908 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 5902 8304 5908 8316
rect 5960 8344 5966 8356
rect 6270 8344 6276 8356
rect 5960 8316 6276 8344
rect 5960 8304 5966 8316
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6420 8316 6561 8344
rect 6420 8304 6426 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 7524 8316 7573 8344
rect 7524 8304 7530 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 8478 8344 8484 8356
rect 8439 8316 8484 8344
rect 7561 8307 7619 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 4430 8276 4436 8288
rect 3436 8248 4436 8276
rect 2409 8239 2467 8245
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 6380 8276 6408 8304
rect 5224 8248 6408 8276
rect 6457 8279 6515 8285
rect 5224 8236 5230 8248
rect 6457 8245 6469 8279
rect 6503 8276 6515 8279
rect 6822 8276 6828 8288
rect 6503 8248 6828 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9858 8276 9864 8288
rect 9732 8248 9864 8276
rect 9732 8236 9738 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10980 8276 11008 8452
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12434 8480 12440 8492
rect 11931 8452 12440 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 14099 8489 14105 8492
rect 14093 8443 14105 8489
rect 14157 8480 14163 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14157 8452 14565 8480
rect 14099 8440 14105 8443
rect 14157 8440 14163 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14820 8483 14878 8489
rect 14820 8449 14832 8483
rect 14866 8480 14878 8483
rect 15028 8480 15056 8508
rect 14866 8452 15056 8480
rect 14866 8449 14878 8452
rect 14820 8443 14878 8449
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 16761 8483 16819 8489
rect 15252 8452 15617 8480
rect 15252 8440 15258 8452
rect 11072 8412 11100 8440
rect 11974 8412 11980 8424
rect 11072 8384 11836 8412
rect 11935 8384 11980 8412
rect 11808 8356 11836 8384
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8381 12127 8415
rect 12526 8412 12532 8424
rect 12487 8384 12532 8412
rect 12069 8375 12127 8381
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11112 8316 11529 8344
rect 11112 8304 11118 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 11790 8304 11796 8356
rect 11848 8344 11854 8356
rect 12084 8344 12112 8375
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 15589 8412 15617 8452
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 16206 8412 16212 8424
rect 15589 8384 16212 8412
rect 16206 8372 16212 8384
rect 16264 8412 16270 8424
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 16264 8384 16405 8412
rect 16264 8372 16270 8384
rect 16393 8381 16405 8384
rect 16439 8412 16451 8415
rect 16776 8412 16804 8443
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 17920 8452 17969 8480
rect 17920 8440 17926 8452
rect 17957 8449 17969 8452
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 16439 8384 16804 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16908 8384 17233 8412
rect 16908 8372 16914 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 14461 8347 14519 8353
rect 14461 8344 14473 8347
rect 11848 8316 12112 8344
rect 14108 8316 14473 8344
rect 11848 8304 11854 8316
rect 11333 8279 11391 8285
rect 11333 8276 11345 8279
rect 10980 8248 11345 8276
rect 11333 8245 11345 8248
rect 11379 8245 11391 8279
rect 11333 8239 11391 8245
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 14108 8276 14136 8316
rect 14461 8313 14473 8316
rect 14507 8344 14519 8347
rect 14507 8316 14596 8344
rect 14507 8313 14519 8316
rect 14461 8307 14519 8313
rect 13044 8248 14136 8276
rect 14277 8279 14335 8285
rect 13044 8236 13050 8248
rect 14277 8245 14289 8279
rect 14323 8276 14335 8279
rect 14366 8276 14372 8288
rect 14323 8248 14372 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14568 8276 14596 8316
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 16025 8347 16083 8353
rect 16025 8344 16037 8347
rect 15620 8316 16037 8344
rect 15620 8304 15626 8316
rect 16025 8313 16037 8316
rect 16071 8344 16083 8347
rect 17420 8344 17448 8375
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 17736 8384 18337 8412
rect 17736 8372 17742 8384
rect 18325 8381 18337 8384
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18138 8344 18144 8356
rect 16071 8316 17448 8344
rect 18099 8316 18144 8344
rect 16071 8313 16083 8316
rect 16025 8307 16083 8313
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 15470 8276 15476 8288
rect 14568 8248 15476 8276
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 15712 8248 16221 8276
rect 15712 8236 15718 8248
rect 16209 8245 16221 8248
rect 16255 8276 16267 8279
rect 17126 8276 17132 8288
rect 16255 8248 17132 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17862 8276 17868 8288
rect 17823 8248 17868 8276
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 2682 8032 2688 8084
rect 2740 8032 2746 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3234 8072 3240 8084
rect 2832 8044 3240 8072
rect 2832 8032 2838 8044
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3605 8075 3663 8081
rect 3605 8072 3617 8075
rect 3476 8044 3617 8072
rect 3476 8032 3482 8044
rect 3605 8041 3617 8044
rect 3651 8072 3663 8075
rect 4062 8072 4068 8084
rect 3651 8044 4068 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 5258 8072 5264 8084
rect 4755 8044 5264 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5902 8072 5908 8084
rect 5644 8044 5908 8072
rect 2700 8004 2728 8032
rect 2700 7976 2912 8004
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2682 7936 2688 7948
rect 2179 7908 2688 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1544 7840 1777 7868
rect 1544 7828 1550 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 2056 7868 2084 7899
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 2884 7945 2912 7976
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 4212 7976 4261 8004
rect 4212 7964 4218 7976
rect 4249 7973 4261 7976
rect 4295 8004 4307 8007
rect 4295 7976 5396 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7905 2927 7939
rect 2869 7899 2927 7905
rect 2774 7868 2780 7880
rect 2056 7840 2780 7868
rect 1765 7831 1823 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 2884 7868 2912 7899
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 5368 7945 5396 7976
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3752 7908 4353 7936
rect 3752 7896 3758 7908
rect 4341 7905 4353 7908
rect 4387 7936 4399 7939
rect 5353 7939 5411 7945
rect 4387 7908 5120 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4430 7868 4436 7880
rect 2884 7840 4436 7868
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4982 7868 4988 7880
rect 4663 7840 4988 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5092 7877 5120 7908
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5644 7936 5672 8044
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 8386 8072 8392 8084
rect 6788 8044 8392 8072
rect 6788 8032 6794 8044
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 8478 8004 8484 8016
rect 5736 7976 8484 8004
rect 5736 7945 5764 7976
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 8772 8004 8800 8035
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 9674 8072 9680 8084
rect 8941 8035 8999 8041
rect 9416 8044 9680 8072
rect 9416 8004 9444 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 11974 8072 11980 8084
rect 11747 8044 11980 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12492 8044 12541 8072
rect 12492 8032 12498 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 13909 8075 13967 8081
rect 13909 8072 13921 8075
rect 12529 8035 12587 8041
rect 13004 8044 13921 8072
rect 8772 7976 9444 8004
rect 10781 8007 10839 8013
rect 10781 7973 10793 8007
rect 10827 8004 10839 8007
rect 11146 8004 11152 8016
rect 10827 7976 11152 8004
rect 10827 7973 10839 7976
rect 10781 7967 10839 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 5399 7908 5672 7936
rect 5721 7939 5779 7945
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 6546 7936 6552 7948
rect 6507 7908 6552 7936
rect 5721 7899 5779 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7834 7936 7840 7948
rect 6880 7908 7328 7936
rect 7795 7908 7840 7936
rect 6880 7896 6886 7908
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 2746 7772 3065 7800
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1452 7704 1593 7732
rect 1452 7692 1458 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 2222 7732 2228 7744
rect 2183 7704 2228 7732
rect 1581 7695 1639 7701
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 2593 7735 2651 7741
rect 2593 7701 2605 7735
rect 2639 7732 2651 7735
rect 2746 7732 2774 7772
rect 3053 7769 3065 7772
rect 3099 7769 3111 7803
rect 3878 7800 3884 7812
rect 3839 7772 3884 7800
rect 3053 7763 3111 7769
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 6733 7803 6791 7809
rect 6733 7769 6745 7803
rect 6779 7800 6791 7803
rect 7300 7800 7328 7908
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8754 7936 8760 7948
rect 8251 7908 8760 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 11296 7908 11345 7936
rect 11296 7896 11302 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12066 7936 12072 7948
rect 11756 7908 12072 7936
rect 11756 7896 11762 7908
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 13004 7945 13032 8044
rect 13909 8041 13921 8044
rect 13955 8072 13967 8075
rect 14918 8072 14924 8084
rect 13955 8044 14924 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 17586 8072 17592 8084
rect 15028 8044 17592 8072
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 13633 8007 13691 8013
rect 13633 8004 13645 8007
rect 13596 7976 13645 8004
rect 13596 7964 13602 7976
rect 13633 7973 13645 7976
rect 13679 7973 13691 8007
rect 13633 7967 13691 7973
rect 14090 7964 14096 8016
rect 14148 8004 14154 8016
rect 15028 8004 15056 8044
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 17862 8032 17868 8084
rect 17920 8032 17926 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 14148 7976 15056 8004
rect 17880 8004 17908 8032
rect 18230 8004 18236 8016
rect 17880 7976 18236 8004
rect 14148 7964 14154 7976
rect 18230 7964 18236 7976
rect 18288 7964 18294 8016
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7905 13047 7939
rect 13170 7936 13176 7948
rect 13131 7908 13176 7936
rect 12989 7899 13047 7905
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 10321 7871 10379 7877
rect 7432 7840 9720 7868
rect 7432 7828 7438 7840
rect 8389 7803 8447 7809
rect 8389 7800 8401 7803
rect 6779 7772 7236 7800
rect 7300 7772 8401 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 2639 7704 2774 7732
rect 2639 7701 2651 7704
rect 2593 7695 2651 7701
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 2961 7735 3019 7741
rect 2961 7732 2973 7735
rect 2924 7704 2973 7732
rect 2924 7692 2930 7704
rect 2961 7701 2973 7704
rect 3007 7701 3019 7735
rect 2961 7695 3019 7701
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3510 7732 3516 7744
rect 3467 7704 3516 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 4062 7732 4068 7744
rect 4023 7704 4068 7732
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4948 7704 5181 7732
rect 4948 7692 4954 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 5810 7732 5816 7744
rect 5771 7704 5816 7732
rect 5169 7695 5227 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 6178 7732 6184 7744
rect 5951 7704 6184 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6638 7732 6644 7744
rect 6328 7704 6373 7732
rect 6599 7704 6644 7732
rect 6328 7692 6334 7704
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7208 7741 7236 7772
rect 8389 7769 8401 7772
rect 8435 7769 8447 7803
rect 9692 7800 9720 7840
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10054 7803 10112 7809
rect 10054 7800 10066 7803
rect 9692 7772 10066 7800
rect 8389 7763 8447 7769
rect 10054 7769 10066 7772
rect 10100 7800 10112 7803
rect 10226 7800 10232 7812
rect 10100 7772 10232 7800
rect 10100 7769 10112 7772
rect 10054 7763 10112 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 6972 7704 7113 7732
rect 6972 7692 6978 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7524 7704 7573 7732
rect 7524 7692 7530 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8110 7732 8116 7744
rect 7699 7704 8116 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9766 7732 9772 7744
rect 8996 7704 9772 7732
rect 8996 7692 9002 7704
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10336 7732 10364 7831
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 10928 7840 11284 7868
rect 10928 7828 10934 7840
rect 11256 7809 11284 7840
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11974 7868 11980 7880
rect 11480 7840 11980 7868
rect 11480 7828 11486 7840
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12360 7868 12388 7899
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 12360 7840 12434 7868
rect 10689 7803 10747 7809
rect 10689 7769 10701 7803
rect 10735 7800 10747 7803
rect 11149 7803 11207 7809
rect 11149 7800 11161 7803
rect 10735 7772 11161 7800
rect 10735 7769 10747 7772
rect 10689 7763 10747 7769
rect 11149 7769 11161 7772
rect 11195 7769 11207 7803
rect 11149 7763 11207 7769
rect 11241 7803 11299 7809
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 12161 7803 12219 7809
rect 12161 7800 12173 7803
rect 11287 7772 12173 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 12161 7769 12173 7772
rect 12207 7769 12219 7803
rect 12406 7800 12434 7840
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12584 7840 12909 7868
rect 12584 7828 12590 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12710 7800 12716 7812
rect 12406 7772 12716 7800
rect 12161 7763 12219 7769
rect 12066 7732 12072 7744
rect 9916 7704 10364 7732
rect 12027 7704 12072 7732
rect 9916 7692 9922 7704
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12176 7732 12204 7763
rect 12710 7760 12716 7772
rect 12768 7800 12774 7812
rect 13188 7800 13216 7896
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 14200 7868 14228 7899
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 15286 7936 15292 7948
rect 14608 7908 15292 7936
rect 14608 7896 14614 7908
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 16632 7908 17049 7936
rect 16632 7896 16638 7908
rect 17037 7905 17049 7908
rect 17083 7905 17095 7939
rect 17037 7899 17095 7905
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 18046 7936 18052 7948
rect 18003 7908 18052 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 18046 7896 18052 7908
rect 18104 7936 18110 7948
rect 18322 7936 18328 7948
rect 18104 7908 18328 7936
rect 18104 7896 18110 7908
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 14458 7868 14464 7880
rect 13688 7840 14228 7868
rect 14419 7840 14464 7868
rect 13688 7828 13694 7840
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 15160 7840 16405 7868
rect 15160 7828 15166 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17126 7868 17132 7880
rect 16991 7840 17132 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17126 7828 17132 7840
rect 17184 7868 17190 7880
rect 17494 7868 17500 7880
rect 17184 7840 17500 7868
rect 17184 7828 17190 7840
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 18138 7868 18144 7880
rect 18099 7840 18144 7868
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 12768 7772 13216 7800
rect 14369 7803 14427 7809
rect 12768 7760 12774 7772
rect 14369 7769 14381 7803
rect 14415 7800 14427 7803
rect 16022 7800 16028 7812
rect 14415 7772 16028 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 16114 7760 16120 7812
rect 16172 7809 16178 7812
rect 16172 7800 16184 7809
rect 16850 7800 16856 7812
rect 16172 7772 16217 7800
rect 16763 7772 16856 7800
rect 16172 7763 16184 7772
rect 16172 7760 16178 7763
rect 16850 7760 16856 7772
rect 16908 7800 16914 7812
rect 17402 7800 17408 7812
rect 16908 7772 17408 7800
rect 16908 7760 16914 7772
rect 17402 7760 17408 7772
rect 17460 7760 17466 7812
rect 12618 7732 12624 7744
rect 12176 7704 12624 7732
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13357 7735 13415 7741
rect 13357 7732 13369 7735
rect 13136 7704 13369 7732
rect 13136 7692 13142 7704
rect 13357 7701 13369 7704
rect 13403 7701 13415 7735
rect 13357 7695 13415 7701
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14792 7704 14841 7732
rect 14792 7692 14798 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 14829 7695 14887 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 16132 7732 16160 7760
rect 15252 7704 16160 7732
rect 15252 7692 15258 7704
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 16448 7704 16497 7732
rect 16448 7692 16454 7704
rect 16485 7701 16497 7704
rect 16531 7701 16543 7735
rect 16485 7695 16543 7701
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17000 7704 17325 7732
rect 17000 7692 17006 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17678 7732 17684 7744
rect 17639 7704 17684 7732
rect 17313 7695 17371 7701
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 18506 7732 18512 7744
rect 17828 7704 18512 7732
rect 17828 7692 17834 7704
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1762 7528 1768 7540
rect 1723 7500 1768 7528
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 1946 7488 1952 7540
rect 2004 7528 2010 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2004 7500 2237 7528
rect 2004 7488 2010 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2866 7528 2872 7540
rect 2827 7500 2872 7528
rect 2225 7491 2283 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3878 7528 3884 7540
rect 3375 7500 3884 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 1857 7463 1915 7469
rect 1857 7460 1869 7463
rect 1636 7432 1869 7460
rect 1636 7420 1642 7432
rect 1857 7429 1869 7432
rect 1903 7429 1915 7463
rect 1857 7423 1915 7429
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 3344 7460 3372 7491
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5810 7528 5816 7540
rect 5399 7500 5816 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6178 7528 6184 7540
rect 6139 7500 6184 7528
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 6546 7528 6552 7540
rect 6507 7500 6552 7528
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 7745 7531 7803 7537
rect 6604 7500 7696 7528
rect 6604 7488 6610 7500
rect 6730 7460 6736 7472
rect 2740 7432 3372 7460
rect 5644 7432 6736 7460
rect 2740 7420 2746 7432
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 2593 7355 2651 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 3602 7392 3608 7404
rect 3528 7364 3608 7392
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2038 7324 2044 7336
rect 1719 7296 2044 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2038 7284 2044 7296
rect 2096 7284 2102 7336
rect 2774 7284 2780 7336
rect 2832 7324 2838 7336
rect 3528 7333 3556 7364
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3988 7364 4169 7392
rect 3513 7327 3571 7333
rect 3513 7324 3525 7327
rect 2832 7296 3525 7324
rect 2832 7284 2838 7296
rect 3513 7293 3525 7296
rect 3559 7293 3571 7327
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3513 7287 3571 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 3050 7256 3056 7268
rect 2455 7228 3056 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 3050 7216 3056 7228
rect 3108 7216 3114 7268
rect 3988 7256 4016 7364
rect 4157 7361 4169 7364
rect 4203 7392 4215 7395
rect 4338 7392 4344 7404
rect 4203 7364 4344 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5258 7392 5264 7404
rect 5031 7364 5264 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 5644 7333 5672 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 6932 7432 7297 7460
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6546 7392 6552 7404
rect 5859 7364 6552 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 4801 7327 4859 7333
rect 4120 7296 4165 7324
rect 4120 7284 4126 7296
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 4847 7296 5641 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 3896 7228 4016 7256
rect 4525 7259 4583 7265
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3896 7188 3924 7228
rect 4525 7225 4537 7259
rect 4571 7256 4583 7259
rect 5736 7256 5764 7287
rect 4571 7228 5764 7256
rect 4571 7225 4583 7228
rect 4525 7219 4583 7225
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 6932 7265 6960 7432
rect 7285 7429 7297 7432
rect 7331 7429 7343 7463
rect 7285 7423 7343 7429
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7558 7392 7564 7404
rect 7423 7364 7564 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 7668 7392 7696 7500
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 7926 7528 7932 7540
rect 7791 7500 7932 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8352 7500 8953 7528
rect 8352 7488 8358 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 9548 7500 10241 7528
rect 9548 7488 9554 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 10229 7491 10287 7497
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 11146 7528 11152 7540
rect 11011 7500 11152 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11885 7531 11943 7537
rect 11885 7528 11897 7531
rect 11379 7500 11897 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11885 7497 11897 7500
rect 11931 7497 11943 7531
rect 13078 7528 13084 7540
rect 13039 7500 13084 7528
rect 11885 7491 11943 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13495 7500 13921 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 14734 7528 14740 7540
rect 14695 7500 14740 7528
rect 13909 7491 13967 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 15703 7500 17509 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 17957 7531 18015 7537
rect 17957 7497 17969 7531
rect 18003 7528 18015 7531
rect 18230 7528 18236 7540
rect 18003 7500 18236 7528
rect 18003 7497 18015 7500
rect 17957 7491 18015 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 12618 7460 12624 7472
rect 8496 7432 12434 7460
rect 12531 7432 12624 7460
rect 8496 7401 8524 7432
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 7668 7364 8493 7392
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8846 7392 8852 7404
rect 8619 7364 8852 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 10134 7392 10140 7404
rect 10095 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 10468 7364 11989 7392
rect 10468 7352 10474 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 6917 7259 6975 7265
rect 6917 7256 6929 7259
rect 5868 7228 6929 7256
rect 5868 7216 5874 7228
rect 6917 7225 6929 7228
rect 6963 7225 6975 7259
rect 7116 7256 7144 7287
rect 7190 7256 7196 7268
rect 7116 7228 7196 7256
rect 6917 7219 6975 7225
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 7576 7256 7604 7352
rect 8018 7324 8024 7336
rect 7979 7296 8024 7324
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 9398 7324 9404 7336
rect 8812 7296 8905 7324
rect 9359 7296 9404 7324
rect 8812 7284 8818 7296
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9582 7324 9588 7336
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 8386 7256 8392 7268
rect 7576 7228 8392 7256
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 8772 7256 8800 7284
rect 10336 7256 10364 7287
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10560 7296 10701 7324
rect 10560 7284 10566 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11422 7324 11428 7336
rect 10919 7296 11428 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11940 7296 12081 7324
rect 11940 7284 11946 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 10594 7256 10600 7268
rect 8772 7228 10600 7256
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 12406 7256 12434 7432
rect 12618 7420 12624 7432
rect 12676 7460 12682 7472
rect 13538 7460 13544 7472
rect 12676 7432 13544 7460
rect 12676 7420 12682 7432
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 13872 7432 14013 7460
rect 13872 7420 13878 7432
rect 14001 7429 14013 7432
rect 14047 7429 14059 7463
rect 14001 7423 14059 7429
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 16666 7460 16672 7472
rect 14608 7432 16672 7460
rect 14608 7420 14614 7432
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 18417 7463 18475 7469
rect 18417 7460 18429 7463
rect 16776 7432 18429 7460
rect 12986 7392 12992 7404
rect 12947 7364 12992 7392
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 15565 7395 15623 7401
rect 14108 7364 15056 7392
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 13354 7324 13360 7336
rect 12943 7296 13360 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 13354 7284 13360 7296
rect 13412 7324 13418 7336
rect 13630 7324 13636 7336
rect 13412 7296 13636 7324
rect 13412 7284 13418 7296
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 14108 7333 14136 7364
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 15028 7333 15056 7364
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16209 7395 16267 7401
rect 15611 7364 16169 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14240 7296 14841 7324
rect 14240 7284 14246 7296
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15194 7324 15200 7336
rect 15059 7296 15200 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7293 15899 7327
rect 16141 7324 16169 7364
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16574 7392 16580 7404
rect 16255 7364 16580 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16574 7352 16580 7364
rect 16632 7392 16638 7404
rect 16776 7392 16804 7432
rect 18417 7429 18429 7432
rect 18463 7429 18475 7463
rect 18417 7423 18475 7429
rect 16632 7364 16804 7392
rect 17037 7395 17095 7401
rect 16632 7352 16638 7364
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17402 7392 17408 7404
rect 17083 7364 17408 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 17586 7352 17592 7404
rect 17644 7392 17650 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17644 7364 17877 7392
rect 17644 7352 17650 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 18322 7392 18328 7404
rect 17865 7355 17923 7361
rect 18156 7364 18328 7392
rect 16758 7324 16764 7336
rect 16141 7296 16764 7324
rect 15841 7287 15899 7293
rect 14734 7256 14740 7268
rect 12406 7228 14740 7256
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 15856 7256 15884 7287
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 18156 7333 18184 7364
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 17221 7327 17279 7333
rect 17221 7293 17233 7327
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 18141 7327 18199 7333
rect 18141 7293 18153 7327
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 16393 7259 16451 7265
rect 14976 7228 16344 7256
rect 14976 7216 14982 7228
rect 2823 7160 3924 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5718 7188 5724 7200
rect 5040 7160 5724 7188
rect 5040 7148 5046 7160
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6604 7160 6653 7188
rect 6604 7148 6610 7160
rect 6641 7157 6653 7160
rect 6687 7188 6699 7191
rect 6822 7188 6828 7200
rect 6687 7160 6828 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 11514 7188 11520 7200
rect 11475 7160 11520 7188
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12434 7188 12440 7200
rect 12124 7160 12440 7188
rect 12124 7148 12130 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 13688 7160 14381 7188
rect 13688 7148 13694 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 14516 7160 15209 7188
rect 14516 7148 14522 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15896 7160 16037 7188
rect 15896 7148 15902 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16316 7188 16344 7228
rect 16393 7225 16405 7259
rect 16439 7256 16451 7259
rect 16482 7256 16488 7268
rect 16439 7228 16488 7256
rect 16439 7225 16451 7228
rect 16393 7219 16451 7225
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 16666 7256 16672 7268
rect 16627 7228 16672 7256
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 16942 7216 16948 7268
rect 17000 7256 17006 7268
rect 17144 7256 17172 7287
rect 17000 7228 17172 7256
rect 17000 7216 17006 7228
rect 17236 7188 17264 7287
rect 16316 7160 17264 7188
rect 16025 7151 16083 7157
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1489 6987 1547 6993
rect 1489 6953 1501 6987
rect 1535 6984 1547 6987
rect 1578 6984 1584 6996
rect 1535 6956 1584 6984
rect 1535 6953 1547 6956
rect 1489 6947 1547 6953
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 2130 6944 2136 6996
rect 2188 6944 2194 6996
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 3602 6984 3608 6996
rect 3476 6956 3608 6984
rect 3476 6944 3482 6956
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 4893 6987 4951 6993
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 5258 6984 5264 6996
rect 4939 6956 5264 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7524 6956 7941 6984
rect 7524 6944 7530 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9306 6984 9312 6996
rect 8444 6956 9312 6984
rect 8444 6944 8450 6956
rect 9306 6944 9312 6956
rect 9364 6984 9370 6996
rect 10226 6984 10232 6996
rect 9364 6956 10232 6984
rect 9364 6944 9370 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12492 6956 15148 6984
rect 12492 6944 12498 6956
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 2038 6848 2044 6860
rect 1811 6820 2044 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2148 6780 2176 6944
rect 8754 6916 8760 6928
rect 4632 6888 5212 6916
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 3142 6848 3148 6860
rect 3099 6820 3148 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 4028 6820 4537 6848
rect 4028 6808 4034 6820
rect 4525 6817 4537 6820
rect 4571 6848 4583 6851
rect 4632 6848 4660 6888
rect 4571 6820 4660 6848
rect 4709 6851 4767 6857
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 5074 6848 5080 6860
rect 4755 6820 5080 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5184 6848 5212 6888
rect 7576 6888 8432 6916
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5184 6820 5365 6848
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 5902 6848 5908 6860
rect 5583 6820 5908 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 7576 6857 7604 6888
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 6380 6820 7573 6848
rect 2056 6752 2176 6780
rect 2685 6783 2743 6789
rect 2056 6724 2084 6752
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2866 6780 2872 6792
rect 2731 6752 2872 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3510 6780 3516 6792
rect 3283 6752 3516 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 6380 6789 6408 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7742 6848 7748 6860
rect 7703 6820 7748 6848
rect 7561 6811 7619 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8404 6857 8432 6888
rect 8588 6888 8760 6916
rect 8588 6857 8616 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 9493 6919 9551 6925
rect 9493 6885 9505 6919
rect 9539 6885 9551 6919
rect 9493 6879 9551 6885
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6817 8631 6851
rect 9306 6848 9312 6860
rect 8573 6811 8631 6817
rect 8864 6820 9312 6848
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 3660 6752 6009 6780
rect 3660 6740 3666 6752
rect 5997 6749 6009 6752
rect 6043 6780 6055 6783
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 6043 6752 6377 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6696 6752 7696 6780
rect 6696 6740 6702 6752
rect 2038 6672 2044 6724
rect 2096 6672 2102 6724
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 3016 6684 4445 6712
rect 3016 6672 3022 6684
rect 4433 6681 4445 6684
rect 4479 6712 4491 6715
rect 6822 6712 6828 6724
rect 4479 6684 6828 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 7009 6715 7067 6721
rect 7009 6681 7021 6715
rect 7055 6712 7067 6715
rect 7469 6715 7527 6721
rect 7469 6712 7481 6715
rect 7055 6684 7481 6712
rect 7055 6681 7067 6684
rect 7009 6675 7067 6681
rect 7469 6681 7481 6684
rect 7515 6681 7527 6715
rect 7668 6712 7696 6752
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8076 6752 8309 6780
rect 8076 6740 8082 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8404 6780 8432 6811
rect 8864 6780 8892 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9508 6848 9536 6879
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 11149 6919 11207 6925
rect 11149 6916 11161 6919
rect 9640 6888 11161 6916
rect 9640 6876 9646 6888
rect 11149 6885 11161 6888
rect 11195 6916 11207 6919
rect 12158 6916 12164 6928
rect 11195 6888 12164 6916
rect 11195 6885 11207 6888
rect 11149 6879 11207 6885
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 15010 6916 15016 6928
rect 13740 6888 15016 6916
rect 9416 6820 9536 6848
rect 9416 6780 9444 6820
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9732 6820 9965 6848
rect 9732 6808 9738 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10965 6851 11023 6857
rect 10965 6817 10977 6851
rect 11011 6848 11023 6851
rect 11238 6848 11244 6860
rect 11011 6820 11244 6848
rect 11011 6817 11023 6820
rect 10965 6811 11023 6817
rect 11238 6808 11244 6820
rect 11296 6848 11302 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11296 6820 11989 6848
rect 11296 6808 11302 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 12802 6848 12808 6860
rect 12763 6820 12808 6848
rect 11977 6811 12035 6817
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13740 6857 13768 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15120 6916 15148 6956
rect 16022 6944 16028 6996
rect 16080 6984 16086 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 16080 6956 16681 6984
rect 16080 6944 16086 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 16669 6947 16727 6953
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17000 6956 17509 6984
rect 17000 6944 17006 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 18138 6916 18144 6928
rect 15120 6888 18144 6916
rect 18138 6876 18144 6888
rect 18196 6876 18202 6928
rect 18322 6876 18328 6928
rect 18380 6876 18386 6928
rect 13725 6851 13783 6857
rect 12952 6820 13676 6848
rect 12952 6808 12958 6820
rect 8404 6752 8892 6780
rect 8956 6752 9444 6780
rect 8297 6743 8355 6749
rect 8956 6712 8984 6752
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9824 6752 9873 6780
rect 9824 6740 9830 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 11146 6780 11152 6792
rect 9861 6743 9919 6749
rect 9968 6752 11152 6780
rect 7668 6684 8984 6712
rect 7469 6675 7527 6681
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 9968 6712 9996 6752
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11480 6752 11805 6780
rect 11480 6740 11486 6752
rect 11793 6749 11805 6752
rect 11839 6780 11851 6783
rect 11882 6780 11888 6792
rect 11839 6752 11888 6780
rect 11839 6749 11851 6752
rect 11793 6743 11851 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 12912 6780 12940 6808
rect 12667 6752 12940 6780
rect 13449 6783 13507 6789
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13538 6780 13544 6792
rect 13495 6752 13544 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13648 6780 13676 6820
rect 13725 6817 13737 6851
rect 13771 6817 13783 6851
rect 14274 6848 14280 6860
rect 14235 6820 14280 6848
rect 13725 6811 13783 6817
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14458 6848 14464 6860
rect 14419 6820 14464 6848
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 14884 6820 15669 6848
rect 14884 6808 14890 6820
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 13998 6780 14004 6792
rect 13648 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14550 6780 14556 6792
rect 14511 6752 14556 6780
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 15672 6780 15700 6811
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 15804 6820 16405 6848
rect 15804 6808 15810 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 17184 6820 17233 6848
rect 17184 6808 17190 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17221 6811 17279 6817
rect 17328 6820 18061 6848
rect 15930 6780 15936 6792
rect 15672 6752 15936 6780
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16206 6780 16212 6792
rect 16167 6752 16212 6780
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17328 6780 17356 6820
rect 18049 6817 18061 6820
rect 18095 6848 18107 6851
rect 18340 6848 18368 6876
rect 18095 6820 18368 6848
rect 18095 6817 18107 6820
rect 18049 6811 18107 6817
rect 18138 6780 18144 6792
rect 16724 6752 17356 6780
rect 17420 6752 18144 6780
rect 16724 6740 16730 6752
rect 10781 6715 10839 6721
rect 9364 6684 9996 6712
rect 10060 6684 10732 6712
rect 9364 6672 9370 6684
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2314 6644 2320 6656
rect 2004 6616 2049 6644
rect 2275 6616 2320 6644
rect 2004 6604 2010 6616
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2774 6644 2780 6656
rect 2547 6616 2780 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3510 6644 3516 6656
rect 3191 6616 3516 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3786 6644 3792 6656
rect 3651 6616 3792 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4154 6644 4160 6656
rect 4111 6616 4160 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 4672 6616 5273 6644
rect 4672 6604 4678 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 5810 6644 5816 6656
rect 5408 6616 5816 6644
rect 5408 6604 5414 6616
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6178 6644 6184 6656
rect 6139 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6730 6644 6736 6656
rect 6691 6616 6736 6644
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 9180 6616 9229 6644
rect 9180 6604 9186 6616
rect 9217 6613 9229 6616
rect 9263 6644 9275 6647
rect 10060 6644 10088 6684
rect 10704 6656 10732 6684
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 10827 6684 12296 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 10318 6644 10324 6656
rect 9263 6616 10088 6644
rect 10279 6616 10324 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10686 6644 10692 6656
rect 10647 6616 10692 6644
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 12268 6653 12296 6684
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13170 6712 13176 6724
rect 12952 6684 13176 6712
rect 12952 6672 12958 6684
rect 13170 6672 13176 6684
rect 13228 6712 13234 6724
rect 17310 6712 17316 6724
rect 13228 6684 16344 6712
rect 13228 6672 13234 6684
rect 12253 6647 12311 6653
rect 11940 6616 11985 6644
rect 11940 6604 11946 6616
rect 12253 6613 12265 6647
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12676 6616 12725 6644
rect 12676 6604 12682 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 13078 6644 13084 6656
rect 13039 6616 13084 6644
rect 12713 6607 12771 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14884 6616 14933 6644
rect 14884 6604 14890 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15194 6644 15200 6656
rect 15059 6616 15200 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 16316 6653 16344 6684
rect 17052 6684 17316 6712
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 15841 6647 15899 6653
rect 15841 6644 15853 6647
rect 15519 6616 15853 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 15841 6613 15853 6616
rect 15887 6613 15899 6647
rect 15841 6607 15899 6613
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 16482 6644 16488 6656
rect 16347 6616 16488 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17052 6653 17080 6684
rect 17310 6672 17316 6684
rect 17368 6672 17374 6724
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 17000 6616 17049 6644
rect 17000 6604 17006 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17420 6644 17448 6752
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18322 6740 18328 6792
rect 18380 6780 18386 6792
rect 19242 6780 19248 6792
rect 18380 6752 19248 6780
rect 18380 6740 18386 6752
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 17862 6712 17868 6724
rect 17823 6684 17868 6712
rect 17862 6672 17868 6684
rect 17920 6712 17926 6724
rect 18782 6712 18788 6724
rect 17920 6684 18788 6712
rect 17920 6672 17926 6684
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 17175 6616 17448 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 17828 6616 17969 6644
rect 17828 6604 17834 6616
rect 17957 6613 17969 6616
rect 18003 6613 18015 6647
rect 18322 6644 18328 6656
rect 18283 6616 18328 6644
rect 17957 6607 18015 6613
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3016 6412 3433 6440
rect 3016 6400 3022 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 3568 6412 3801 6440
rect 3568 6400 3574 6412
rect 3789 6409 3801 6412
rect 3835 6409 3847 6443
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 3789 6403 3847 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4295 6412 4629 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5077 6443 5135 6449
rect 5077 6440 5089 6443
rect 4764 6412 5089 6440
rect 4764 6400 4770 6412
rect 5077 6409 5089 6412
rect 5123 6409 5135 6443
rect 5077 6403 5135 6409
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 6362 6440 6368 6452
rect 5859 6412 6368 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6472 6412 6684 6440
rect 2222 6332 2228 6384
rect 2280 6372 2286 6384
rect 3145 6375 3203 6381
rect 3145 6372 3157 6375
rect 2280 6344 3157 6372
rect 2280 6332 2286 6344
rect 3145 6341 3157 6344
rect 3191 6341 3203 6375
rect 3145 6335 3203 6341
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 6472 6372 6500 6412
rect 5960 6344 6500 6372
rect 5960 6332 5966 6344
rect 6546 6332 6552 6384
rect 6604 6332 6610 6384
rect 6656 6372 6684 6412
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 6788 6412 7665 6440
rect 6788 6400 6794 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 8076 6412 8125 6440
rect 8076 6400 8082 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 8904 6412 9137 6440
rect 8904 6400 8910 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 9125 6403 9183 6409
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9582 6440 9588 6452
rect 9364 6412 9588 6440
rect 9364 6400 9370 6412
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 10318 6440 10324 6452
rect 9723 6412 10324 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10502 6400 10508 6452
rect 10560 6400 10566 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 12802 6440 12808 6452
rect 10652 6412 12808 6440
rect 10652 6400 10658 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13541 6443 13599 6449
rect 13541 6409 13553 6443
rect 13587 6440 13599 6443
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 13587 6412 14013 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 14001 6409 14013 6412
rect 14047 6409 14059 6443
rect 14001 6403 14059 6409
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 14148 6412 14473 6440
rect 14148 6400 14154 6412
rect 14461 6409 14473 6412
rect 14507 6440 14519 6443
rect 15010 6440 15016 6452
rect 14507 6412 15016 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 15194 6440 15200 6452
rect 15155 6412 15200 6440
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 15335 6412 15669 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 15657 6409 15669 6412
rect 15703 6409 15715 6443
rect 15657 6403 15715 6409
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 16071 6412 17509 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 17497 6409 17509 6412
rect 17543 6409 17555 6443
rect 17497 6403 17555 6409
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 17865 6443 17923 6449
rect 17865 6440 17877 6443
rect 17644 6412 17877 6440
rect 17644 6400 17650 6412
rect 17865 6409 17877 6412
rect 17911 6409 17923 6443
rect 17865 6403 17923 6409
rect 17957 6443 18015 6449
rect 17957 6409 17969 6443
rect 18003 6440 18015 6443
rect 19334 6440 19340 6452
rect 18003 6412 19340 6440
rect 18003 6409 18015 6412
rect 17957 6403 18015 6409
rect 8754 6372 8760 6384
rect 6656 6344 7972 6372
rect 8715 6344 8760 6372
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1535 6276 1869 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1857 6273 1869 6276
rect 1903 6304 1915 6307
rect 1946 6304 1952 6316
rect 1903 6276 1952 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3602 6304 3608 6316
rect 3099 6276 3608 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 3752 6276 4997 6304
rect 3752 6264 3758 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 2958 6168 2964 6180
rect 2915 6140 2964 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 5000 6168 5028 6267
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 6564 6304 6592 6332
rect 6730 6304 6736 6316
rect 5684 6276 6592 6304
rect 6691 6276 6736 6304
rect 5684 6264 5690 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7282 6304 7288 6316
rect 7156 6276 7288 6304
rect 7156 6264 7162 6276
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 5132 6208 5181 6236
rect 5132 6196 5138 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5316 6208 5917 6236
rect 5316 6196 5322 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6454 6236 6460 6248
rect 6052 6208 6097 6236
rect 6415 6208 6460 6236
rect 6052 6196 6058 6208
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 6638 6236 6644 6248
rect 6599 6208 6644 6236
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 7742 6236 7748 6248
rect 6748 6208 7420 6236
rect 7703 6208 7748 6236
rect 6748 6168 6776 6208
rect 5000 6140 6776 6168
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 7064 6140 7297 6168
rect 7064 6128 7070 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 5442 6100 5448 6112
rect 5403 6072 5448 6100
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 7101 6103 7159 6109
rect 7101 6069 7113 6103
rect 7147 6100 7159 6103
rect 7190 6100 7196 6112
rect 7147 6072 7196 6100
rect 7147 6069 7159 6072
rect 7101 6063 7159 6069
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7392 6100 7420 6208
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 7944 6245 7972 6344
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 10520 6372 10548 6400
rect 9692 6344 10548 6372
rect 11333 6375 11391 6381
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 8938 6304 8944 6316
rect 8711 6276 8944 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9692 6304 9720 6344
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 11422 6372 11428 6384
rect 11379 6344 11428 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 11790 6332 11796 6384
rect 11848 6372 11854 6384
rect 11848 6344 12112 6372
rect 11848 6332 11854 6344
rect 9508 6276 9720 6304
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8202 6236 8208 6248
rect 7975 6208 8208 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 9508 6245 9536 6276
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 9824 6276 10180 6304
rect 9824 6264 9830 6276
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8628 6208 8861 6236
rect 8628 6196 8634 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 9950 6236 9956 6248
rect 9631 6208 9956 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10152 6236 10180 6276
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10284 6276 10517 6304
rect 10284 6264 10290 6276
rect 10505 6273 10517 6276
rect 10551 6304 10563 6307
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10551 6276 11069 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 11057 6273 11069 6276
rect 11103 6304 11115 6307
rect 11698 6304 11704 6316
rect 11103 6276 11704 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10152 6208 10609 6236
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10778 6236 10784 6248
rect 10739 6208 10784 6236
rect 10597 6199 10655 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 12084 6245 12112 6344
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 14369 6375 14427 6381
rect 14369 6372 14381 6375
rect 12216 6344 14381 6372
rect 12216 6332 12222 6344
rect 14369 6341 14381 6344
rect 14415 6372 14427 6375
rect 15838 6372 15844 6384
rect 14415 6344 15844 6372
rect 14415 6341 14427 6344
rect 14369 6335 14427 6341
rect 15838 6332 15844 6344
rect 15896 6332 15902 6384
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 16945 6375 17003 6381
rect 16945 6372 16957 6375
rect 16816 6344 16957 6372
rect 16816 6332 16822 6344
rect 16945 6341 16957 6344
rect 16991 6341 17003 6375
rect 17972 6372 18000 6403
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 16945 6335 17003 6341
rect 17880 6344 18000 6372
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6304 12771 6307
rect 12894 6304 12900 6316
rect 12759 6276 12900 6304
rect 12759 6273 12771 6276
rect 12713 6267 12771 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13262 6304 13268 6316
rect 13004 6276 13268 6304
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 11480 6208 11989 6236
rect 11480 6196 11486 6208
rect 11977 6205 11989 6208
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12618 6196 12624 6248
rect 12676 6236 12682 6248
rect 13004 6245 13032 6276
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 17037 6307 17095 6313
rect 15988 6276 16252 6304
rect 15988 6264 15994 6276
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12676 6208 12817 6236
rect 12676 6196 12682 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 12989 6199 13047 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 14090 6236 14096 6248
rect 13495 6208 14096 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 7760 6168 7788 6196
rect 8018 6168 8024 6180
rect 7760 6140 8024 6168
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 9858 6168 9864 6180
rect 8128 6140 9864 6168
rect 8128 6100 8156 6140
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 10045 6171 10103 6177
rect 10045 6137 10057 6171
rect 10091 6168 10103 6171
rect 10410 6168 10416 6180
rect 10091 6140 10416 6168
rect 10091 6137 10103 6140
rect 10045 6131 10103 6137
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11204 6140 11529 6168
rect 11204 6128 11210 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 13909 6171 13967 6177
rect 13909 6137 13921 6171
rect 13955 6168 13967 6171
rect 14182 6168 14188 6180
rect 13955 6140 14188 6168
rect 13955 6137 13967 6140
rect 13909 6131 13967 6137
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 14660 6168 14688 6199
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15344 6208 15393 6236
rect 15344 6196 15350 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 16114 6236 16120 6248
rect 16075 6208 16120 6236
rect 15381 6199 15439 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16224 6245 16252 6276
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16724 6208 16773 6236
rect 16724 6196 16730 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 17052 6236 17080 6267
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 17880 6304 17908 6344
rect 18322 6304 18328 6316
rect 17828 6276 17908 6304
rect 18064 6276 18328 6304
rect 17828 6264 17834 6276
rect 18064 6236 18092 6276
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 17052 6208 18092 6236
rect 18141 6239 18199 6245
rect 16761 6199 16819 6205
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 14918 6168 14924 6180
rect 14660 6140 14924 6168
rect 14918 6128 14924 6140
rect 14976 6168 14982 6180
rect 17126 6168 17132 6180
rect 14976 6140 17132 6168
rect 14976 6128 14982 6140
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 17402 6168 17408 6180
rect 17363 6140 17408 6168
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 18156 6168 18184 6199
rect 17972 6140 18184 6168
rect 8294 6100 8300 6112
rect 7392 6072 8156 6100
rect 8255 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10226 6100 10232 6112
rect 10183 6072 10232 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 12345 6103 12403 6109
rect 12345 6069 12357 6103
rect 12391 6100 12403 6103
rect 12526 6100 12532 6112
rect 12391 6072 12532 6100
rect 12391 6069 12403 6072
rect 12345 6063 12403 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14792 6072 14841 6100
rect 14792 6060 14798 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 15654 6100 15660 6112
rect 15160 6072 15660 6100
rect 15160 6060 15166 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 17972 6100 18000 6140
rect 18322 6100 18328 6112
rect 15804 6072 18000 6100
rect 18283 6072 18328 6100
rect 15804 6060 15810 6072
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2556 5868 2697 5896
rect 2556 5856 2562 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 2924 5868 3065 5896
rect 2924 5856 2930 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3053 5859 3111 5865
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 3602 5896 3608 5908
rect 3375 5868 3608 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 3878 5896 3884 5908
rect 3839 5868 3884 5896
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4522 5896 4528 5908
rect 4435 5868 4528 5896
rect 4522 5856 4528 5868
rect 4580 5896 4586 5908
rect 5258 5896 5264 5908
rect 4580 5868 5264 5896
rect 4580 5856 4586 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5905 5899 5963 5905
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6730 5896 6736 5908
rect 5951 5868 6736 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 9950 5896 9956 5908
rect 6880 5868 8800 5896
rect 9911 5868 9956 5896
rect 6880 5856 6886 5868
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 3421 5831 3479 5837
rect 3421 5828 3433 5831
rect 2372 5800 3433 5828
rect 2372 5788 2378 5800
rect 3421 5797 3433 5800
rect 3467 5797 3479 5831
rect 3421 5791 3479 5797
rect 4341 5831 4399 5837
rect 4341 5797 4353 5831
rect 4387 5828 4399 5831
rect 4614 5828 4620 5840
rect 4387 5800 4620 5828
rect 4387 5797 4399 5800
rect 4341 5791 4399 5797
rect 2501 5763 2559 5769
rect 2501 5729 2513 5763
rect 2547 5760 2559 5763
rect 2590 5760 2596 5772
rect 2547 5732 2596 5760
rect 2547 5729 2559 5732
rect 2501 5723 2559 5729
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 3436 5760 3464 5791
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 4893 5831 4951 5837
rect 4893 5797 4905 5831
rect 4939 5828 4951 5831
rect 5810 5828 5816 5840
rect 4939 5800 5816 5828
rect 4939 5797 4951 5800
rect 4893 5791 4951 5797
rect 4985 5763 5043 5769
rect 4985 5760 4997 5763
rect 3436 5732 4997 5760
rect 4985 5729 4997 5732
rect 5031 5760 5043 5763
rect 5166 5760 5172 5772
rect 5031 5732 5172 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1544 5664 1777 5692
rect 1544 5652 1550 5664
rect 1765 5661 1777 5664
rect 1811 5692 1823 5695
rect 2038 5692 2044 5704
rect 1811 5664 2044 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 2130 5624 2136 5636
rect 1360 5596 2136 5624
rect 1360 5584 1366 5596
rect 2130 5584 2136 5596
rect 2188 5624 2194 5636
rect 2317 5627 2375 5633
rect 2317 5624 2329 5627
rect 2188 5596 2329 5624
rect 2188 5584 2194 5596
rect 2317 5593 2329 5596
rect 2363 5593 2375 5627
rect 2317 5587 2375 5593
rect 3970 5584 3976 5636
rect 4028 5624 4034 5636
rect 4028 5596 4752 5624
rect 4028 5584 4034 5596
rect 4724 5568 4752 5596
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2222 5556 2228 5568
rect 2004 5528 2228 5556
rect 2004 5516 2010 5528
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 3510 5556 3516 5568
rect 3007 5528 3516 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 4706 5556 4712 5568
rect 4667 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5000 5556 5028 5723
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5368 5769 5396 5800
rect 5810 5788 5816 5800
rect 5868 5828 5874 5840
rect 8662 5828 8668 5840
rect 5868 5800 6960 5828
rect 5868 5788 5874 5800
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 5500 5732 5545 5760
rect 5500 5720 5506 5732
rect 5994 5720 6000 5772
rect 6052 5760 6058 5772
rect 6454 5760 6460 5772
rect 6052 5732 6460 5760
rect 6052 5720 6058 5732
rect 6454 5720 6460 5732
rect 6512 5760 6518 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6512 5732 6561 5760
rect 6512 5720 6518 5732
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 5534 5692 5540 5704
rect 5495 5664 5540 5692
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 5644 5664 6377 5692
rect 5644 5556 5672 5664
rect 6365 5661 6377 5664
rect 6411 5692 6423 5695
rect 6822 5692 6828 5704
rect 6411 5664 6828 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6932 5701 6960 5800
rect 7116 5800 8668 5828
rect 7116 5769 7144 5800
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5729 7159 5763
rect 7101 5723 7159 5729
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7248 5732 7297 5760
rect 7248 5720 7254 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8570 5760 8576 5772
rect 7975 5732 8576 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7944 5692 7972 5723
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 6963 5664 7972 5692
rect 8772 5692 8800 5868
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11940 5868 12081 5896
rect 11940 5856 11946 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 13814 5896 13820 5908
rect 13775 5868 13820 5896
rect 12069 5859 12127 5865
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 15378 5896 15384 5908
rect 15243 5868 15384 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 16114 5896 16120 5908
rect 16071 5868 16120 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17862 5896 17868 5908
rect 17460 5868 17868 5896
rect 17460 5856 17466 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18414 5896 18420 5908
rect 18375 5868 18420 5896
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 11238 5828 11244 5840
rect 9416 5800 11244 5828
rect 8938 5760 8944 5772
rect 8899 5732 8944 5760
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9416 5769 9444 5800
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 13262 5828 13268 5840
rect 12406 5800 13268 5828
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 10367 5732 11529 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 11517 5729 11529 5732
rect 11563 5760 11575 5763
rect 12406 5760 12434 5800
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 13372 5800 15148 5828
rect 12526 5760 12532 5772
rect 11563 5732 12434 5760
rect 12487 5732 12532 5760
rect 11563 5729 11575 5732
rect 11517 5723 11575 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 11882 5692 11888 5704
rect 8772 5664 11888 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12728 5692 12756 5720
rect 12492 5664 12756 5692
rect 12492 5652 12498 5664
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12860 5664 13277 5692
rect 12860 5652 12866 5664
rect 13265 5661 13277 5664
rect 13311 5692 13323 5695
rect 13372 5692 13400 5800
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5760 13599 5763
rect 13722 5760 13728 5772
rect 13587 5732 13728 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 14918 5760 14924 5772
rect 14783 5732 14924 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 13311 5664 13400 5692
rect 15120 5692 15148 5800
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 16853 5831 16911 5837
rect 16853 5828 16865 5831
rect 15988 5800 16865 5828
rect 15988 5788 15994 5800
rect 16853 5797 16865 5800
rect 16899 5797 16911 5831
rect 16853 5791 16911 5797
rect 17218 5788 17224 5840
rect 17276 5788 17282 5840
rect 17310 5788 17316 5840
rect 17368 5828 17374 5840
rect 17681 5831 17739 5837
rect 17681 5828 17693 5831
rect 17368 5800 17693 5828
rect 17368 5788 17374 5800
rect 17681 5797 17693 5800
rect 17727 5797 17739 5831
rect 17681 5791 17739 5797
rect 15746 5760 15752 5772
rect 15707 5732 15752 5760
rect 15746 5720 15752 5732
rect 15804 5760 15810 5772
rect 15804 5732 16344 5760
rect 15804 5720 15810 5732
rect 16316 5692 16344 5732
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 16485 5763 16543 5769
rect 16485 5760 16497 5763
rect 16448 5732 16497 5760
rect 16448 5720 16454 5732
rect 16485 5729 16497 5732
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5729 16635 5763
rect 17236 5760 17264 5788
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17236 5732 17417 5760
rect 16577 5723 16635 5729
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 16592 5692 16620 5723
rect 15120 5664 16068 5692
rect 16316 5664 16620 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 6457 5627 6515 5633
rect 6457 5624 6469 5627
rect 5736 5596 6469 5624
rect 5736 5568 5764 5596
rect 6457 5593 6469 5596
rect 6503 5624 6515 5627
rect 6730 5624 6736 5636
rect 6503 5596 6736 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7650 5624 7656 5636
rect 7392 5596 7656 5624
rect 5000 5528 5672 5556
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 7392 5565 7420 5596
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 7834 5584 7840 5636
rect 7892 5624 7898 5636
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 7892 5596 8401 5624
rect 7892 5584 7898 5596
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 10318 5584 10324 5636
rect 10376 5624 10382 5636
rect 11333 5627 11391 5633
rect 10376 5596 11192 5624
rect 10376 5584 10382 5596
rect 7377 5559 7435 5565
rect 6052 5528 6097 5556
rect 6052 5516 6058 5528
rect 7377 5525 7389 5559
rect 7423 5525 7435 5559
rect 7377 5519 7435 5525
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7616 5528 7757 5556
rect 7616 5516 7622 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 8018 5556 8024 5568
rect 7979 5528 8024 5556
rect 7745 5519 7803 5525
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 9490 5556 9496 5568
rect 9451 5528 9496 5556
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 9640 5528 9685 5556
rect 9640 5516 9646 5528
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 10410 5556 10416 5568
rect 9916 5528 10416 5556
rect 9916 5516 9922 5528
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 10870 5556 10876 5568
rect 10560 5528 10605 5556
rect 10831 5528 10876 5556
rect 10560 5516 10566 5528
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11164 5556 11192 5596
rect 11333 5593 11345 5627
rect 11379 5624 11391 5627
rect 11379 5596 11652 5624
rect 11379 5593 11391 5596
rect 11333 5587 11391 5593
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 11020 5528 11065 5556
rect 11164 5528 11437 5556
rect 11020 5516 11026 5528
rect 11425 5525 11437 5528
rect 11471 5525 11483 5559
rect 11624 5556 11652 5596
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 11756 5596 14473 5624
rect 11756 5584 11762 5596
rect 14461 5593 14473 5596
rect 14507 5624 14519 5627
rect 15105 5627 15163 5633
rect 14507 5596 15056 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 11790 5556 11796 5568
rect 11624 5528 11796 5556
rect 11425 5519 11483 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12342 5556 12348 5568
rect 12032 5528 12348 5556
rect 12032 5516 12038 5528
rect 12342 5516 12348 5528
rect 12400 5556 12406 5568
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 12400 5528 12449 5556
rect 12400 5516 12406 5528
rect 12437 5525 12449 5528
rect 12483 5556 12495 5559
rect 12526 5556 12532 5568
rect 12483 5528 12532 5556
rect 12483 5525 12495 5528
rect 12437 5519 12495 5525
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 12894 5556 12900 5568
rect 12855 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 13412 5528 13457 5556
rect 13412 5516 13418 5528
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 14553 5559 14611 5565
rect 14553 5556 14565 5559
rect 14148 5528 14565 5556
rect 14148 5516 14154 5528
rect 14553 5525 14565 5528
rect 14599 5556 14611 5559
rect 14918 5556 14924 5568
rect 14599 5528 14924 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15028 5556 15056 5596
rect 15105 5593 15117 5627
rect 15151 5624 15163 5627
rect 15565 5627 15623 5633
rect 15565 5624 15577 5627
rect 15151 5596 15577 5624
rect 15151 5593 15163 5596
rect 15105 5587 15163 5593
rect 15565 5593 15577 5596
rect 15611 5593 15623 5627
rect 15565 5587 15623 5593
rect 16040 5568 16068 5664
rect 17034 5652 17040 5704
rect 17092 5692 17098 5704
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17092 5664 17325 5692
rect 17092 5652 17098 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 15194 5556 15200 5568
rect 15028 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15654 5556 15660 5568
rect 15615 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16022 5516 16028 5568
rect 16080 5556 16086 5568
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 16080 5528 16405 5556
rect 16080 5516 16086 5528
rect 16393 5525 16405 5528
rect 16439 5525 16451 5559
rect 17218 5556 17224 5568
rect 17179 5528 17224 5556
rect 16393 5519 16451 5525
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 17310 5516 17316 5568
rect 17368 5556 17374 5568
rect 17420 5556 17448 5723
rect 17862 5692 17868 5704
rect 17823 5664 17868 5692
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18598 5692 18604 5704
rect 18279 5664 18604 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 17368 5528 17448 5556
rect 17368 5516 17374 5528
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 2406 5352 2412 5364
rect 1964 5324 2412 5352
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 1964 5284 1992 5324
rect 2406 5312 2412 5324
rect 2464 5352 2470 5364
rect 4062 5352 4068 5364
rect 2464 5324 3096 5352
rect 4023 5324 4068 5352
rect 2464 5312 2470 5324
rect 1719 5256 1992 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2222 5244 2228 5296
rect 2280 5284 2286 5296
rect 2869 5287 2927 5293
rect 2869 5284 2881 5287
rect 2280 5256 2881 5284
rect 2280 5244 2286 5256
rect 2869 5253 2881 5256
rect 2915 5253 2927 5287
rect 2869 5247 2927 5253
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2424 5148 2452 5179
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3068 5216 3096 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 5994 5352 6000 5364
rect 5859 5324 6000 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6638 5352 6644 5364
rect 6227 5324 6644 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 7190 5352 7196 5364
rect 6963 5324 7196 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 7190 5312 7196 5324
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 3326 5284 3332 5296
rect 3287 5256 3332 5284
rect 3326 5244 3332 5256
rect 3384 5244 3390 5296
rect 5261 5287 5319 5293
rect 5261 5284 5273 5287
rect 4172 5256 5273 5284
rect 4172 5216 4200 5256
rect 5261 5253 5273 5256
rect 5307 5284 5319 5287
rect 5718 5284 5724 5296
rect 5307 5256 5724 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5718 5244 5724 5256
rect 5776 5244 5782 5296
rect 6454 5284 6460 5296
rect 6415 5256 6460 5284
rect 6454 5244 6460 5256
rect 6512 5284 6518 5296
rect 6733 5287 6791 5293
rect 6733 5284 6745 5287
rect 6512 5256 6745 5284
rect 6512 5244 6518 5256
rect 6733 5253 6745 5256
rect 6779 5253 6791 5287
rect 6733 5247 6791 5253
rect 2832 5188 2877 5216
rect 3068 5188 4200 5216
rect 4249 5219 4307 5225
rect 2832 5176 2838 5188
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 5810 5216 5816 5228
rect 4295 5188 4476 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 3326 5148 3332 5160
rect 2424 5120 3332 5148
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3476 5120 3521 5148
rect 3476 5108 3482 5120
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 2774 5080 2780 5092
rect 2639 5052 2780 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 4448 5089 4476 5188
rect 5552 5188 5816 5216
rect 5552 5157 5580 5188
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7064 5188 7297 5216
rect 7064 5176 7070 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7392 5216 7420 5315
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7800 5324 7849 5352
rect 7800 5312 7806 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8294 5352 8300 5364
rect 8251 5324 8300 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9582 5352 9588 5364
rect 9539 5324 9588 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 10226 5352 10232 5364
rect 10091 5324 10232 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10870 5352 10876 5364
rect 10831 5324 10876 5352
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5352 11299 5355
rect 11422 5352 11428 5364
rect 11287 5324 11428 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 13320 5324 13369 5352
rect 13320 5312 13326 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 15102 5352 15108 5364
rect 13357 5315 13415 5321
rect 13464 5324 15108 5352
rect 9125 5287 9183 5293
rect 9125 5253 9137 5287
rect 9171 5284 9183 5287
rect 10502 5284 10508 5296
rect 9171 5256 10508 5284
rect 9171 5253 9183 5256
rect 9125 5247 9183 5253
rect 7650 5216 7656 5228
rect 7392 5188 7656 5216
rect 7285 5179 7343 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8076 5188 8309 5216
rect 8076 5176 8082 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 9140 5216 9168 5247
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 10962 5284 10968 5296
rect 10827 5256 10968 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11974 5284 11980 5296
rect 11935 5256 11980 5284
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 13464 5293 13492 5324
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15286 5352 15292 5364
rect 15247 5324 15292 5352
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16264 5324 16313 5352
rect 16264 5312 16270 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17497 5355 17555 5361
rect 17497 5352 17509 5355
rect 17276 5324 17509 5352
rect 17276 5312 17282 5324
rect 17497 5321 17509 5324
rect 17543 5321 17555 5355
rect 17497 5315 17555 5321
rect 18417 5355 18475 5361
rect 18417 5321 18429 5355
rect 18463 5352 18475 5355
rect 18782 5352 18788 5364
rect 18463 5324 18788 5352
rect 18463 5321 18475 5324
rect 18417 5315 18475 5321
rect 18782 5312 18788 5324
rect 18840 5352 18846 5364
rect 19150 5352 19156 5364
rect 18840 5324 19156 5352
rect 18840 5312 18846 5324
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 12452 5256 13461 5284
rect 8297 5179 8355 5185
rect 8496 5188 9168 5216
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5684 5120 5733 5148
rect 5684 5108 5690 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 6638 5148 6644 5160
rect 5721 5111 5779 5117
rect 6472 5120 6644 5148
rect 4433 5083 4491 5089
rect 4433 5049 4445 5083
rect 4479 5080 4491 5083
rect 6472 5080 6500 5120
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 8386 5148 8392 5160
rect 7524 5120 7696 5148
rect 8347 5120 8392 5148
rect 7524 5108 7530 5120
rect 4479 5052 6500 5080
rect 7668 5080 7696 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 7668 5052 7757 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 7745 5043 7803 5049
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2924 4984 3065 5012
rect 2924 4972 2930 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 8496 5012 8524 5188
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9732 5188 9965 5216
rect 9732 5176 9738 5188
rect 9953 5185 9965 5188
rect 9999 5216 10011 5219
rect 10226 5216 10232 5228
rect 9999 5188 10232 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 10376 5188 11713 5216
rect 10376 5176 10382 5188
rect 11701 5185 11713 5188
rect 11747 5216 11759 5219
rect 11790 5216 11796 5228
rect 11747 5188 11796 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11790 5176 11796 5188
rect 11848 5216 11854 5228
rect 12452 5216 12480 5256
rect 13449 5253 13461 5256
rect 13495 5253 13507 5287
rect 13449 5247 13507 5253
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14332 5256 15148 5284
rect 14332 5244 14338 5256
rect 11848 5188 12480 5216
rect 12529 5219 12587 5225
rect 11848 5176 11854 5188
rect 12529 5185 12541 5219
rect 12575 5216 12587 5219
rect 12575 5188 13860 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5117 8999 5151
rect 8941 5111 8999 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9858 5148 9864 5160
rect 9079 5120 9864 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 8956 5080 8984 5111
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10134 5148 10140 5160
rect 10095 5120 10140 5148
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5117 10747 5151
rect 12434 5148 12440 5160
rect 10689 5111 10747 5117
rect 10888 5120 12440 5148
rect 10594 5080 10600 5092
rect 8956 5052 10600 5080
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 10704 5080 10732 5111
rect 10888 5080 10916 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12618 5148 12624 5160
rect 12579 5120 12624 5148
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 13446 5148 13452 5160
rect 12851 5120 13452 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13630 5148 13636 5160
rect 13591 5120 13636 5148
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 10704 5052 10916 5080
rect 11882 5040 11888 5092
rect 11940 5080 11946 5092
rect 12161 5083 12219 5089
rect 12161 5080 12173 5083
rect 11940 5052 12173 5080
rect 11940 5040 11946 5052
rect 12161 5049 12173 5052
rect 12207 5049 12219 5083
rect 12161 5043 12219 5049
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 12526 5080 12532 5092
rect 12308 5052 12532 5080
rect 12308 5040 12314 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12989 5083 13047 5089
rect 12989 5049 13001 5083
rect 13035 5080 13047 5083
rect 13354 5080 13360 5092
rect 13035 5052 13360 5080
rect 13035 5049 13047 5052
rect 12989 5043 13047 5049
rect 13354 5040 13360 5052
rect 13412 5040 13418 5092
rect 13832 5089 13860 5188
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13964 5188 14197 5216
rect 13964 5176 13970 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 15120 5225 15148 5256
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 16850 5284 16856 5296
rect 16172 5256 16856 5284
rect 16172 5244 16178 5256
rect 16850 5244 16856 5256
rect 16908 5284 16914 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 16908 5256 17049 5284
rect 16908 5244 16914 5256
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 17037 5247 17095 5253
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14608 5188 14749 5216
rect 14608 5176 14614 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15105 5179 15163 5185
rect 15304 5188 15853 5216
rect 15304 5160 15332 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 17144 5216 17172 5244
rect 17770 5216 17776 5228
rect 17144 5188 17776 5216
rect 15841 5179 15899 5185
rect 17770 5176 17776 5188
rect 17828 5176 17834 5228
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 14148 5120 14289 5148
rect 14148 5108 14154 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14642 5148 14648 5160
rect 14516 5120 14648 5148
rect 14516 5108 14522 5120
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5117 15623 5151
rect 15746 5148 15752 5160
rect 15707 5120 15752 5148
rect 15565 5111 15623 5117
rect 13817 5083 13875 5089
rect 13817 5049 13829 5083
rect 13863 5049 13875 5083
rect 13817 5043 13875 5049
rect 14921 5083 14979 5089
rect 14921 5049 14933 5083
rect 14967 5080 14979 5083
rect 15194 5080 15200 5092
rect 14967 5052 15200 5080
rect 14967 5049 14979 5052
rect 14921 5043 14979 5049
rect 15194 5040 15200 5052
rect 15252 5040 15258 5092
rect 15470 5040 15476 5092
rect 15528 5080 15534 5092
rect 15580 5080 15608 5111
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 17000 5120 17141 5148
rect 17000 5108 17006 5120
rect 17129 5117 17141 5120
rect 17175 5117 17187 5151
rect 17310 5148 17316 5160
rect 17271 5120 17316 5148
rect 17129 5111 17187 5117
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 17328 5080 17356 5108
rect 15528 5052 17356 5080
rect 15528 5040 15534 5052
rect 9582 5012 9588 5024
rect 4764 4984 8524 5012
rect 9543 4984 9588 5012
rect 4764 4972 4770 4984
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10410 5012 10416 5024
rect 9916 4984 10416 5012
rect 9916 4972 9922 4984
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 10560 4984 11621 5012
rect 10560 4972 10566 4984
rect 11609 4981 11621 4984
rect 11655 5012 11667 5015
rect 15102 5012 15108 5024
rect 11655 4984 15108 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 16172 4984 16221 5012
rect 16172 4972 16178 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 16448 4984 16681 5012
rect 16448 4972 16454 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 16669 4975 16727 4981
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 2188 4780 2329 4808
rect 2188 4768 2194 4780
rect 2317 4777 2329 4780
rect 2363 4777 2375 4811
rect 2317 4771 2375 4777
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2832 4780 2973 4808
rect 2832 4768 2838 4780
rect 2961 4777 2973 4780
rect 3007 4808 3019 4811
rect 3878 4808 3884 4820
rect 3007 4780 3884 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 8754 4808 8760 4820
rect 6012 4780 8156 4808
rect 8715 4780 8760 4808
rect 5258 4700 5264 4752
rect 5316 4740 5322 4752
rect 6012 4740 6040 4780
rect 6362 4740 6368 4752
rect 5316 4712 6040 4740
rect 6196 4712 6368 4740
rect 5316 4700 5322 4712
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 1688 4644 3157 4672
rect 1688 4613 1716 4644
rect 3145 4641 3157 4644
rect 3191 4672 3203 4675
rect 3191 4644 5212 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 1820 4576 1865 4604
rect 1820 4564 1826 4576
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 2832 4576 2877 4604
rect 2832 4564 2838 4576
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 5184 4604 5212 4644
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5960 4644 6101 4672
rect 5960 4632 5966 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6196 4604 6224 4712
rect 6362 4700 6368 4712
rect 6420 4740 6426 4752
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 6420 4712 6561 4740
rect 6420 4700 6426 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 8128 4740 8156 4780
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9398 4808 9404 4820
rect 9088 4780 9404 4808
rect 9088 4768 9094 4780
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9548 4780 9873 4808
rect 9548 4768 9554 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 11885 4811 11943 4817
rect 11885 4808 11897 4811
rect 11388 4780 11897 4808
rect 11388 4768 11394 4780
rect 11885 4777 11897 4780
rect 11931 4777 11943 4811
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 11885 4771 11943 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12713 4811 12771 4817
rect 12713 4808 12725 4811
rect 12676 4780 12725 4808
rect 12676 4768 12682 4780
rect 12713 4777 12725 4780
rect 12759 4777 12771 4811
rect 12713 4771 12771 4777
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 13228 4780 13553 4808
rect 13228 4768 13234 4780
rect 13541 4777 13553 4780
rect 13587 4777 13599 4811
rect 13541 4771 13599 4777
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 15470 4808 15476 4820
rect 13872 4780 14688 4808
rect 13872 4768 13878 4780
rect 14550 4740 14556 4752
rect 7156 4712 8064 4740
rect 8128 4712 14556 4740
rect 7156 4700 7162 4712
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6454 4672 6460 4684
rect 6319 4644 6460 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 7374 4672 7380 4684
rect 7331 4644 7380 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 8036 4681 8064 4712
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 8067 4644 9597 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 9585 4641 9597 4644
rect 9631 4672 9643 4675
rect 10134 4672 10140 4684
rect 9631 4644 10140 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10318 4672 10324 4684
rect 10279 4644 10324 4672
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10594 4672 10600 4684
rect 10551 4644 10600 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 12621 4675 12679 4681
rect 11296 4644 11341 4672
rect 11296 4632 11302 4644
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12802 4672 12808 4684
rect 12667 4644 12808 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13173 4675 13231 4681
rect 13173 4672 13185 4675
rect 12952 4644 13185 4672
rect 12952 4632 12958 4644
rect 13173 4641 13185 4644
rect 13219 4641 13231 4675
rect 13173 4635 13231 4641
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 14458 4672 14464 4684
rect 13403 4644 14464 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 14660 4681 14688 4780
rect 15028 4780 15476 4808
rect 15028 4681 15056 4780
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 18506 4808 18512 4820
rect 18463 4780 18512 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 15102 4700 15108 4752
rect 15160 4740 15166 4752
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 15160 4712 15761 4740
rect 15160 4700 15166 4712
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 16577 4743 16635 4749
rect 16577 4740 16589 4743
rect 15749 4703 15807 4709
rect 15856 4712 16589 4740
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 15856 4672 15884 4712
rect 16577 4709 16589 4712
rect 16623 4709 16635 4743
rect 16577 4703 16635 4709
rect 18049 4743 18107 4749
rect 18049 4709 18061 4743
rect 18095 4740 18107 4743
rect 18690 4740 18696 4752
rect 18095 4712 18696 4740
rect 18095 4709 18107 4712
rect 18049 4703 18107 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 16298 4672 16304 4684
rect 15243 4644 15884 4672
rect 16259 4644 16304 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4672 17279 4675
rect 17954 4672 17960 4684
rect 17267 4644 17960 4672
rect 17267 4641 17279 4644
rect 17221 4635 17279 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 5184 4576 6224 4604
rect 4985 4567 5043 4573
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 6696 4576 7941 4604
rect 6696 4564 6702 4576
rect 7929 4573 7941 4576
rect 7975 4604 7987 4607
rect 8754 4604 8760 4616
rect 7975 4576 8760 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9490 4604 9496 4616
rect 9364 4576 9496 4604
rect 9364 4564 9370 4576
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9732 4576 10241 4604
rect 9732 4564 9738 4576
rect 10229 4573 10241 4576
rect 10275 4604 10287 4607
rect 10870 4604 10876 4616
rect 10275 4576 10876 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 12115 4576 13829 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 13817 4573 13829 4576
rect 13863 4604 13875 4607
rect 15838 4604 15844 4616
rect 13863 4576 15844 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16632 4576 17509 4604
rect 16632 4564 16638 4576
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 17586 4604 17592 4616
rect 17543 4576 17592 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 17862 4604 17868 4616
rect 17823 4576 17868 4604
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 2041 4539 2099 4545
rect 2041 4505 2053 4539
rect 2087 4536 2099 4539
rect 2958 4536 2964 4548
rect 2087 4508 2964 4536
rect 2087 4505 2099 4508
rect 2041 4499 2099 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 5258 4536 5264 4548
rect 5219 4508 5264 4536
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 7837 4539 7895 4545
rect 5828 4508 7788 4536
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2590 4468 2596 4480
rect 2551 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 5828 4468 5856 4508
rect 5994 4468 6000 4480
rect 4672 4440 5856 4468
rect 5955 4440 6000 4468
rect 4672 4428 4678 4440
rect 5994 4428 6000 4440
rect 6052 4468 6058 4480
rect 6178 4468 6184 4480
rect 6052 4440 6184 4468
rect 6052 4428 6058 4440
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7006 4468 7012 4480
rect 6967 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7156 4440 7201 4468
rect 7156 4428 7162 4440
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7432 4440 7481 4468
rect 7432 4428 7438 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 7760 4468 7788 4508
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 7883 4508 8309 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 11974 4536 11980 4548
rect 8297 4499 8355 4505
rect 8956 4508 11980 4536
rect 8956 4468 8984 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 13081 4539 13139 4545
rect 13081 4505 13093 4539
rect 13127 4536 13139 4539
rect 13127 4508 14136 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 7760 4440 8984 4468
rect 9033 4471 9091 4477
rect 7469 4431 7527 4437
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9306 4468 9312 4480
rect 9079 4440 9312 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 10689 4471 10747 4477
rect 9456 4440 9501 4468
rect 9456 4428 9462 4440
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 10870 4468 10876 4480
rect 10735 4440 10876 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11609 4471 11667 4477
rect 11609 4468 11621 4471
rect 11020 4440 11621 4468
rect 11020 4428 11026 4440
rect 11609 4437 11621 4440
rect 11655 4468 11667 4471
rect 11698 4468 11704 4480
rect 11655 4440 11704 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 11698 4428 11704 4440
rect 11756 4468 11762 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11756 4440 12265 4468
rect 11756 4428 11762 4440
rect 12253 4437 12265 4440
rect 12299 4468 12311 4471
rect 13262 4468 13268 4480
rect 12299 4440 13268 4468
rect 12299 4437 12311 4440
rect 12253 4431 12311 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 14108 4477 14136 4508
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 14240 4508 14473 4536
rect 14240 4496 14246 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 14461 4499 14519 4505
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 15289 4539 15347 4545
rect 15289 4536 15301 4539
rect 15068 4508 15301 4536
rect 15068 4496 15074 4508
rect 15289 4505 15301 4508
rect 15335 4505 15347 4539
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15289 4499 15347 4505
rect 15672 4508 16221 4536
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 15194 4468 15200 4480
rect 14599 4440 15200 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15672 4477 15700 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 16209 4499 16267 4505
rect 16945 4539 17003 4545
rect 16945 4505 16957 4539
rect 16991 4536 17003 4539
rect 17218 4536 17224 4548
rect 16991 4508 17224 4536
rect 16991 4505 17003 4508
rect 16945 4499 17003 4505
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 18248 4536 18276 4567
rect 18012 4508 18276 4536
rect 18012 4496 18018 4508
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 16816 4440 17049 4468
rect 16816 4428 16822 4440
rect 17037 4437 17049 4440
rect 17083 4437 17095 4471
rect 17037 4431 17095 4437
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 5868 4236 6377 4264
rect 5868 4224 5874 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 6365 4227 6423 4233
rect 6454 4224 6460 4276
rect 6512 4264 6518 4276
rect 6641 4267 6699 4273
rect 6641 4264 6653 4267
rect 6512 4236 6653 4264
rect 6512 4224 6518 4236
rect 6641 4233 6653 4236
rect 6687 4233 6699 4267
rect 7006 4264 7012 4276
rect 6967 4236 7012 4264
rect 6641 4227 6699 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7374 4264 7380 4276
rect 7335 4236 7380 4264
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 8294 4264 8300 4276
rect 7524 4236 7569 4264
rect 8255 4236 8300 4264
rect 7524 4224 7530 4236
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 8478 4264 8484 4276
rect 8404 4236 8484 4264
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 5537 4199 5595 4205
rect 2004 4168 5488 4196
rect 2004 4156 2010 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1719 4100 2053 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2041 4097 2053 4100
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2455 4100 2605 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2593 4097 2605 4100
rect 2639 4128 2651 4131
rect 2682 4128 2688 4140
rect 2639 4100 2688 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4128 3019 4131
rect 3142 4128 3148 4140
rect 3007 4100 3148 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 5460 4128 5488 4168
rect 5537 4165 5549 4199
rect 5583 4196 5595 4199
rect 5902 4196 5908 4208
rect 5583 4168 5908 4196
rect 5583 4165 5595 4168
rect 5537 4159 5595 4165
rect 5902 4156 5908 4168
rect 5960 4156 5966 4208
rect 6917 4199 6975 4205
rect 6917 4165 6929 4199
rect 6963 4196 6975 4199
rect 7190 4196 7196 4208
rect 6963 4168 7196 4196
rect 6963 4165 6975 4168
rect 6917 4159 6975 4165
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 8404 4196 8432 4236
rect 8478 4224 8484 4236
rect 8536 4264 8542 4276
rect 8757 4267 8815 4273
rect 8757 4264 8769 4267
rect 8536 4236 8769 4264
rect 8536 4224 8542 4236
rect 8757 4233 8769 4236
rect 8803 4233 8815 4267
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 8757 4227 8815 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9401 4267 9459 4273
rect 9401 4233 9413 4267
rect 9447 4264 9459 4267
rect 9582 4264 9588 4276
rect 9447 4236 9588 4264
rect 9447 4233 9459 4236
rect 9401 4227 9459 4233
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 9861 4267 9919 4273
rect 9861 4233 9873 4267
rect 9907 4264 9919 4267
rect 10502 4264 10508 4276
rect 9907 4236 10508 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 11790 4224 11796 4276
rect 11848 4264 11854 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 11848 4236 12081 4264
rect 11848 4224 11854 4236
rect 12069 4233 12081 4236
rect 12115 4233 12127 4267
rect 12069 4227 12127 4233
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12584 4236 13676 4264
rect 12584 4224 12590 4236
rect 7300 4168 8432 4196
rect 8665 4199 8723 4205
rect 5994 4128 6000 4140
rect 5460 4100 6000 4128
rect 5994 4088 6000 4100
rect 6052 4128 6058 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 6052 4100 6101 4128
rect 6052 4088 6058 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 7300 4128 7328 4168
rect 8665 4165 8677 4199
rect 8711 4196 8723 4199
rect 10045 4199 10103 4205
rect 10045 4196 10057 4199
rect 8711 4168 10057 4196
rect 8711 4165 8723 4168
rect 8665 4159 8723 4165
rect 10045 4165 10057 4168
rect 10091 4196 10103 4199
rect 10410 4196 10416 4208
rect 10091 4168 10416 4196
rect 10091 4165 10103 4168
rect 10045 4159 10103 4165
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 12897 4199 12955 4205
rect 12897 4196 12909 4199
rect 12636 4168 12909 4196
rect 11514 4128 11520 4140
rect 6089 4091 6147 4097
rect 6380 4100 7328 4128
rect 7668 4100 9628 4128
rect 11475 4100 11520 4128
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 6380 4060 6408 4100
rect 7668 4069 7696 4100
rect 3752 4032 6408 4060
rect 7653 4063 7711 4069
rect 3752 4020 3758 4032
rect 7653 4029 7665 4063
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8202 4060 8208 4072
rect 7975 4032 8208 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 9600 4069 9628 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 11606 4060 11612 4072
rect 9631 4032 11612 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 11974 4060 11980 4072
rect 11839 4032 11980 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12636 4060 12664 4168
rect 12897 4165 12909 4168
rect 12943 4165 12955 4199
rect 13648 4196 13676 4236
rect 13722 4224 13728 4276
rect 13780 4264 13786 4276
rect 14090 4264 14096 4276
rect 13780 4236 13825 4264
rect 14051 4236 14096 4264
rect 13780 4224 13786 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14461 4267 14519 4273
rect 14461 4233 14473 4267
rect 14507 4264 14519 4267
rect 14918 4264 14924 4276
rect 14507 4236 14924 4264
rect 14507 4233 14519 4236
rect 14461 4227 14519 4233
rect 14918 4224 14924 4236
rect 14976 4224 14982 4276
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 15197 4267 15255 4273
rect 15197 4264 15209 4267
rect 15160 4236 15209 4264
rect 15160 4224 15166 4236
rect 15197 4233 15209 4236
rect 15243 4233 15255 4267
rect 15930 4264 15936 4276
rect 15891 4236 15936 4264
rect 15197 4227 15255 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17313 4267 17371 4273
rect 17313 4233 17325 4267
rect 17359 4264 17371 4267
rect 17402 4264 17408 4276
rect 17359 4236 17408 4264
rect 17359 4233 17371 4236
rect 17313 4227 17371 4233
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 13648 4168 15240 4196
rect 12897 4159 12955 4165
rect 13633 4131 13691 4137
rect 12728 4100 13584 4128
rect 12728 4069 12756 4100
rect 13556 4072 13584 4100
rect 13633 4097 13645 4131
rect 13679 4128 13691 4131
rect 13998 4128 14004 4140
rect 13679 4100 14004 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 15105 4131 15163 4137
rect 15105 4097 15117 4131
rect 15151 4097 15163 4131
rect 15212 4128 15240 4168
rect 16850 4156 16856 4208
rect 16908 4196 16914 4208
rect 17034 4196 17040 4208
rect 16908 4168 17040 4196
rect 16908 4156 16914 4168
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 15654 4128 15660 4140
rect 15212 4100 15660 4128
rect 15105 4091 15163 4097
rect 12483 4032 12664 4060
rect 12713 4063 12771 4069
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12713 4029 12725 4063
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13538 4060 13544 4072
rect 12860 4032 12905 4060
rect 13499 4032 13544 4060
rect 12860 4020 12866 4032
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 14277 4063 14335 4069
rect 14277 4029 14289 4063
rect 14323 4060 14335 4063
rect 15010 4060 15016 4072
rect 14323 4032 15016 4060
rect 14323 4029 14335 4032
rect 14277 4023 14335 4029
rect 1854 3992 1860 4004
rect 1815 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3952 1918 4004
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 2271 3964 2636 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 2608 3924 2636 3964
rect 2774 3952 2780 4004
rect 2832 3992 2838 4004
rect 2832 3964 2877 3992
rect 2832 3952 2838 3964
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 7156 3964 8953 3992
rect 7156 3952 7162 3964
rect 8941 3961 8953 3964
rect 8987 3961 8999 3995
rect 10226 3992 10232 4004
rect 10139 3964 10232 3992
rect 8941 3955 8999 3961
rect 10226 3952 10232 3964
rect 10284 3992 10290 4004
rect 13265 3995 13323 4001
rect 10284 3964 12434 3992
rect 10284 3952 10290 3964
rect 2866 3924 2872 3936
rect 2608 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 8076 3896 8125 3924
rect 8076 3884 8082 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 8113 3887 8171 3893
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 9548 3896 10333 3924
rect 9548 3884 9554 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10321 3887 10379 3893
rect 10502 3884 10508 3896
rect 10560 3924 10566 3936
rect 11238 3924 11244 3936
rect 10560 3896 11244 3924
rect 10560 3884 10566 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12406 3924 12434 3964
rect 13265 3961 13277 3995
rect 13311 3992 13323 3995
rect 13906 3992 13912 4004
rect 13311 3964 13912 3992
rect 13311 3961 13323 3964
rect 13265 3955 13323 3961
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 14292 3924 14320 4023
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 14553 3995 14611 4001
rect 14553 3961 14565 3995
rect 14599 3992 14611 3995
rect 15120 3992 15148 4091
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4128 16083 4131
rect 16390 4128 16396 4140
rect 16071 4100 16396 4128
rect 16071 4097 16083 4100
rect 16025 4091 16083 4097
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16715 4100 17172 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 15378 4060 15384 4072
rect 15339 4032 15384 4060
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 16206 4060 16212 4072
rect 16167 4032 16212 4060
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 16298 4020 16304 4072
rect 16356 4060 16362 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 16356 4032 16865 4060
rect 16356 4020 16362 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 14599 3964 14863 3992
rect 15120 3964 15577 3992
rect 14599 3961 14611 3964
rect 14553 3955 14611 3961
rect 12406 3896 14320 3924
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 14737 3927 14795 3933
rect 14737 3924 14749 3927
rect 14700 3896 14749 3924
rect 14700 3884 14706 3896
rect 14737 3893 14749 3896
rect 14783 3893 14795 3927
rect 14835 3924 14863 3964
rect 15565 3961 15577 3964
rect 15611 3961 15623 3995
rect 15565 3955 15623 3961
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 16758 3992 16764 4004
rect 16080 3964 16764 3992
rect 16080 3952 16086 3964
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 17034 3952 17040 4004
rect 17092 3992 17098 4004
rect 17144 3992 17172 4100
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17276 4100 17417 4128
rect 17276 4088 17282 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17736 4100 17969 4128
rect 17736 4088 17742 4100
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4060 17647 4063
rect 17862 4060 17868 4072
rect 17635 4032 17868 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 17862 4020 17868 4032
rect 17920 4020 17926 4072
rect 19058 4060 19064 4072
rect 17972 4032 19064 4060
rect 17972 3992 18000 4032
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 18138 3992 18144 4004
rect 17092 3964 18000 3992
rect 18099 3964 18144 3992
rect 17092 3952 17098 3964
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 15470 3924 15476 3936
rect 14835 3896 15476 3924
rect 14737 3887 14795 3893
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 15988 3896 16405 3924
rect 15988 3884 15994 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 18325 3927 18383 3933
rect 18325 3924 18337 3927
rect 16908 3896 18337 3924
rect 16908 3884 16914 3896
rect 18325 3893 18337 3896
rect 18371 3893 18383 3927
rect 18325 3887 18383 3893
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 2406 3720 2412 3732
rect 2367 3692 2412 3720
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 4080 3692 4261 3720
rect 2240 3556 3004 3584
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1535 3488 1869 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 1857 3485 1869 3488
rect 1903 3516 1915 3519
rect 1946 3516 1952 3528
rect 1903 3488 1952 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2240 3525 2268 3556
rect 2976 3525 3004 3556
rect 4080 3525 4108 3692
rect 4249 3689 4261 3692
rect 4295 3720 4307 3723
rect 8202 3720 8208 3732
rect 4295 3692 8208 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8754 3720 8760 3732
rect 8715 3692 8760 3720
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 10318 3720 10324 3732
rect 9815 3692 10324 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13722 3720 13728 3732
rect 13587 3692 13728 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14182 3720 14188 3732
rect 14143 3692 14188 3720
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14550 3720 14556 3732
rect 14511 3692 14556 3720
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 14829 3723 14887 3729
rect 14829 3689 14841 3723
rect 14875 3720 14887 3723
rect 15010 3720 15016 3732
rect 14875 3692 15016 3720
rect 14875 3689 14887 3692
rect 14829 3683 14887 3689
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15194 3680 15200 3732
rect 15252 3680 15258 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15654 3720 15660 3732
rect 15344 3692 15389 3720
rect 15615 3692 15660 3720
rect 15344 3680 15350 3692
rect 15654 3680 15660 3692
rect 15712 3720 15718 3732
rect 16390 3720 16396 3732
rect 15712 3692 16396 3720
rect 15712 3680 15718 3692
rect 16390 3680 16396 3692
rect 16448 3720 16454 3732
rect 16577 3723 16635 3729
rect 16577 3720 16589 3723
rect 16448 3692 16589 3720
rect 16448 3680 16454 3692
rect 16577 3689 16589 3692
rect 16623 3689 16635 3723
rect 16942 3720 16948 3732
rect 16903 3692 16948 3720
rect 16577 3683 16635 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17310 3720 17316 3732
rect 17271 3692 17316 3720
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 18230 3720 18236 3732
rect 18191 3692 18236 3720
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 19242 3720 19248 3732
rect 18555 3692 19248 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 12802 3612 12808 3664
rect 12860 3652 12866 3664
rect 13633 3655 13691 3661
rect 13633 3652 13645 3655
rect 12860 3624 13645 3652
rect 12860 3612 12866 3624
rect 13633 3621 13645 3624
rect 13679 3621 13691 3655
rect 14200 3652 14228 3680
rect 14921 3655 14979 3661
rect 14921 3652 14933 3655
rect 14200 3624 14933 3652
rect 13633 3615 13691 3621
rect 14921 3621 14933 3624
rect 14967 3621 14979 3655
rect 14921 3615 14979 3621
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 8662 3584 8668 3596
rect 6963 3556 8668 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 15102 3584 15108 3596
rect 11287 3556 15108 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15212 3584 15240 3680
rect 15470 3652 15476 3664
rect 15431 3624 15476 3652
rect 15470 3612 15476 3624
rect 15528 3652 15534 3664
rect 17218 3652 17224 3664
rect 15528 3624 17224 3652
rect 15528 3612 15534 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17494 3652 17500 3664
rect 17328 3624 17500 3652
rect 15562 3584 15568 3596
rect 15212 3556 15568 3584
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 16022 3584 16028 3596
rect 15979 3556 16028 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16172 3556 16217 3584
rect 16172 3544 16178 3556
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 17328 3584 17356 3624
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 18966 3584 18972 3596
rect 16448 3556 17356 3584
rect 16448 3544 16454 3556
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 4065 3519 4123 3525
rect 3007 3488 4016 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 2608 3448 2636 3479
rect 2685 3451 2743 3457
rect 2685 3448 2697 3451
rect 2608 3420 2697 3448
rect 2685 3417 2697 3420
rect 2731 3448 2743 3451
rect 3694 3448 3700 3460
rect 2731 3420 3700 3448
rect 2731 3417 2743 3420
rect 2685 3411 2743 3417
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 3988 3448 4016 3488
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 6144 3488 6653 3516
rect 6144 3476 6150 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 7064 3488 7573 3516
rect 7064 3476 7070 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 7561 3479 7619 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10836 3488 10977 3516
rect 10836 3476 10842 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13078 3516 13084 3528
rect 12943 3488 13084 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14056 3488 14289 3516
rect 14056 3476 14062 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 16206 3516 16212 3528
rect 15068 3488 16212 3516
rect 15068 3476 15074 3488
rect 16206 3476 16212 3488
rect 16264 3516 16270 3528
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16264 3488 16773 3516
rect 16264 3476 16270 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3516 17187 3519
rect 17328 3516 17356 3556
rect 17512 3556 18972 3584
rect 17512 3528 17540 3556
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 17494 3516 17500 3528
rect 17175 3488 17356 3516
rect 17407 3488 17500 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3485 17831 3519
rect 18046 3516 18052 3528
rect 18007 3488 18052 3516
rect 17773 3479 17831 3485
rect 7837 3451 7895 3457
rect 3988 3420 4660 3448
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 2041 3383 2099 3389
rect 2041 3349 2053 3383
rect 2087 3380 2099 3383
rect 2774 3380 2780 3392
rect 2087 3352 2780 3380
rect 2087 3349 2099 3352
rect 2041 3343 2099 3349
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4632 3380 4660 3420
rect 7837 3417 7849 3451
rect 7883 3448 7895 3451
rect 8018 3448 8024 3460
rect 7883 3420 8024 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 8018 3408 8024 3420
rect 8076 3408 8082 3460
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 9490 3448 9496 3460
rect 8435 3420 9496 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 12802 3408 12808 3460
rect 12860 3448 12866 3460
rect 13173 3451 13231 3457
rect 13173 3448 13185 3451
rect 12860 3420 13185 3448
rect 12860 3408 12866 3420
rect 13173 3417 13185 3420
rect 13219 3417 13231 3451
rect 13173 3411 13231 3417
rect 17788 3392 17816 3479
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 4890 3380 4896 3392
rect 4632 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3380 4954 3392
rect 9674 3380 9680 3392
rect 4948 3352 9680 3380
rect 4948 3340 4954 3352
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 15562 3380 15568 3392
rect 15243 3352 15568 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 15804 3352 16405 3380
rect 15804 3340 15810 3352
rect 16393 3349 16405 3352
rect 16439 3380 16451 3383
rect 16482 3380 16488 3392
rect 16439 3352 16488 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 17770 3340 17776 3392
rect 17828 3340 17834 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 16206 3176 16212 3188
rect 16167 3148 16212 3176
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16761 3179 16819 3185
rect 16761 3145 16773 3179
rect 16807 3176 16819 3179
rect 17034 3176 17040 3188
rect 16807 3148 17040 3176
rect 16807 3145 16819 3148
rect 16761 3139 16819 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 17402 3176 17408 3188
rect 17359 3148 17408 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18322 3176 18328 3188
rect 18279 3148 18328 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 6236 3080 7849 3108
rect 6236 3068 6242 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 11204 3080 12265 3108
rect 11204 3068 11210 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 14642 3108 14648 3120
rect 12253 3071 12311 3077
rect 12544 3080 14648 3108
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 2087 3012 2145 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2133 3009 2145 3012
rect 2179 3040 2191 3043
rect 2314 3040 2320 3052
rect 2179 3012 2320 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6638 3040 6644 3052
rect 5859 3012 6644 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6748 3012 7021 3040
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 3694 2972 3700 2984
rect 3651 2944 3700 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 4580 2944 5549 2972
rect 4580 2932 4586 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6748 2972 6776 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7340 3012 7573 3040
rect 7340 3000 7346 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 7561 3003 7619 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11164 3012 11836 3040
rect 11164 2981 11192 3012
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 6328 2944 6776 2972
rect 7024 2944 7205 2972
rect 6328 2932 6334 2944
rect 7024 2916 7052 2944
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 7006 2864 7012 2916
rect 7064 2864 7070 2916
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 11716 2904 11744 2935
rect 10376 2876 11744 2904
rect 10376 2864 10382 2876
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 11808 2836 11836 3012
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12544 3049 12572 3080
rect 14642 3068 14648 3080
rect 14700 3068 14706 3120
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 15654 3108 15660 3120
rect 14976 3080 15660 3108
rect 14976 3068 14982 3080
rect 15654 3068 15660 3080
rect 15712 3108 15718 3120
rect 16393 3111 16451 3117
rect 16393 3108 16405 3111
rect 15712 3080 16405 3108
rect 15712 3068 15718 3080
rect 16393 3077 16405 3080
rect 16439 3077 16451 3111
rect 16393 3071 16451 3077
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11940 3012 11989 3040
rect 11940 3000 11946 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 14734 3040 14740 3052
rect 14695 3012 14740 3040
rect 12529 3003 12587 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 15378 3040 15384 3052
rect 14884 3012 14929 3040
rect 15339 3012 15384 3040
rect 14884 3000 14890 3012
rect 15378 3000 15384 3012
rect 15436 3040 15442 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15436 3012 15945 3040
rect 15436 3000 15442 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 16408 3040 16436 3071
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 16945 3111 17003 3117
rect 16945 3108 16957 3111
rect 16632 3080 16957 3108
rect 16632 3068 16638 3080
rect 16945 3077 16957 3080
rect 16991 3077 17003 3111
rect 16945 3071 17003 3077
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 17954 3108 17960 3120
rect 17736 3080 17960 3108
rect 17736 3068 17742 3080
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 16408 3012 17141 3040
rect 15933 3003 15991 3009
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17129 3003 17187 3009
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 18138 3040 18144 3052
rect 18095 3012 18144 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18138 3000 18144 3012
rect 18196 3040 18202 3052
rect 18414 3040 18420 3052
rect 18196 3012 18420 3040
rect 18196 3000 18202 3012
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 13688 2944 14473 2972
rect 13688 2932 13694 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14700 2944 15025 2972
rect 14700 2932 14706 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 17678 2972 17684 2984
rect 15703 2944 17684 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 17678 2932 17684 2944
rect 17736 2932 17742 2984
rect 17773 2975 17831 2981
rect 17773 2941 17785 2975
rect 17819 2972 17831 2975
rect 18598 2972 18604 2984
rect 17819 2944 18604 2972
rect 17819 2941 17831 2944
rect 17773 2935 17831 2941
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 18138 2904 18144 2916
rect 15620 2876 18144 2904
rect 15620 2864 15626 2876
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 15286 2836 15292 2848
rect 11808 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 16482 2796 16488 2848
rect 16540 2836 16546 2848
rect 18417 2839 18475 2845
rect 18417 2836 18429 2839
rect 16540 2808 18429 2836
rect 16540 2796 16546 2808
rect 18417 2805 18429 2808
rect 18463 2805 18475 2839
rect 18417 2799 18475 2805
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16206 2632 16212 2644
rect 16167 2604 16212 2632
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16390 2632 16396 2644
rect 16351 2604 16396 2632
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 16853 2635 16911 2641
rect 16853 2601 16865 2635
rect 16899 2632 16911 2635
rect 17862 2632 17868 2644
rect 16899 2604 17868 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 18506 2632 18512 2644
rect 18095 2604 18512 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 15565 2567 15623 2573
rect 15565 2533 15577 2567
rect 15611 2564 15623 2567
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15611 2536 15945 2564
rect 15611 2533 15623 2536
rect 15565 2527 15623 2533
rect 15933 2533 15945 2536
rect 15979 2564 15991 2567
rect 16666 2564 16672 2576
rect 15979 2536 16672 2564
rect 15979 2533 15991 2536
rect 15933 2527 15991 2533
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 17034 2564 17040 2576
rect 16995 2536 17040 2564
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 17218 2564 17224 2576
rect 17179 2536 17224 2564
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 17954 2564 17960 2576
rect 17819 2536 17960 2564
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 18138 2524 18144 2576
rect 18196 2564 18202 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 18196 2536 18429 2564
rect 18196 2524 18202 2536
rect 18417 2533 18429 2536
rect 18463 2564 18475 2567
rect 19334 2564 19340 2576
rect 18463 2536 19340 2564
rect 18463 2533 18475 2536
rect 18417 2527 18475 2533
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 15010 2496 15016 2508
rect 14971 2468 15016 2496
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 18046 2496 18052 2508
rect 15304 2468 18052 2496
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 15304 2437 15332 2468
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 15289 2431 15347 2437
rect 15289 2428 15301 2431
rect 4304 2400 15301 2428
rect 4304 2388 4310 2400
rect 15289 2397 15301 2400
rect 15335 2397 15347 2431
rect 16574 2428 16580 2440
rect 15289 2391 15347 2397
rect 15948 2400 16580 2428
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 15948 2360 15976 2400
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 17310 2428 17316 2440
rect 16724 2400 17316 2428
rect 16724 2388 16730 2400
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 17405 2431 17463 2437
rect 17405 2397 17417 2431
rect 17451 2428 17463 2431
rect 17862 2428 17868 2440
rect 17451 2400 17724 2428
rect 17823 2400 17868 2428
rect 17451 2397 17463 2400
rect 17405 2391 17463 2397
rect 17586 2360 17592 2372
rect 8260 2332 15976 2360
rect 16040 2332 17592 2360
rect 8260 2320 8266 2332
rect 16040 2304 16068 2332
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 17696 2360 17724 2400
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18690 2360 18696 2372
rect 17696 2332 18696 2360
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 16850 2292 16856 2304
rect 16632 2264 16856 2292
rect 16632 2252 16638 2264
rect 16850 2252 16856 2264
rect 16908 2292 16914 2304
rect 17497 2295 17555 2301
rect 17497 2292 17509 2295
rect 16908 2264 17509 2292
rect 16908 2252 16914 2264
rect 17497 2261 17509 2264
rect 17543 2261 17555 2295
rect 17497 2255 17555 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 4982 1776 4988 1828
rect 5040 1816 5046 1828
rect 16022 1816 16028 1828
rect 5040 1788 16028 1816
rect 5040 1776 5046 1788
rect 16022 1776 16028 1788
rect 16080 1776 16086 1828
<< via1 >>
rect 9220 14968 9272 15020
rect 10324 14968 10376 15020
rect 8576 14900 8628 14952
rect 12624 14900 12676 14952
rect 13084 14900 13136 14952
rect 10048 14832 10100 14884
rect 16948 14832 17000 14884
rect 6828 14764 6880 14816
rect 11612 14764 11664 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 2780 14560 2832 14612
rect 10416 14560 10468 14612
rect 14280 14560 14332 14612
rect 15936 14560 15988 14612
rect 12900 14492 12952 14544
rect 15292 14492 15344 14544
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 9220 14356 9272 14408
rect 9312 14356 9364 14408
rect 13820 14424 13872 14476
rect 12992 14356 13044 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 14832 14356 14884 14408
rect 14924 14356 14976 14408
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 8208 14288 8260 14340
rect 2320 14220 2372 14272
rect 8852 14220 8904 14272
rect 9680 14220 9732 14272
rect 10048 14331 10100 14340
rect 10048 14297 10066 14331
rect 10066 14297 10100 14331
rect 10048 14288 10100 14297
rect 10508 14288 10560 14340
rect 13452 14288 13504 14340
rect 18420 14288 18472 14340
rect 10232 14220 10284 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 13912 14220 13964 14272
rect 17040 14220 17092 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 2964 13948 3016 14000
rect 9772 14016 9824 14068
rect 10232 14016 10284 14068
rect 11612 14016 11664 14068
rect 14096 14016 14148 14068
rect 7380 13948 7432 14000
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 6184 13880 6236 13932
rect 8484 13880 8536 13932
rect 8852 13923 8904 13932
rect 9312 13948 9364 14000
rect 9588 13948 9640 14000
rect 8852 13889 8870 13923
rect 8870 13889 8904 13923
rect 8852 13880 8904 13889
rect 2872 13812 2924 13864
rect 3608 13812 3660 13864
rect 8392 13676 8444 13728
rect 8484 13676 8536 13728
rect 12808 13948 12860 14000
rect 12900 13948 12952 14000
rect 14832 14016 14884 14068
rect 12624 13923 12676 13932
rect 15292 13948 15344 14000
rect 12624 13889 12642 13923
rect 12642 13889 12676 13923
rect 12624 13880 12676 13889
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 11888 13676 11940 13728
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 17592 13948 17644 14000
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 3516 13336 3568 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 3608 13268 3660 13320
rect 6920 13472 6972 13524
rect 8024 13472 8076 13524
rect 9864 13472 9916 13524
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 13176 13472 13228 13524
rect 13544 13472 13596 13524
rect 15200 13472 15252 13524
rect 11704 13447 11756 13456
rect 11704 13413 11713 13447
rect 11713 13413 11747 13447
rect 11747 13413 11756 13447
rect 11704 13404 11756 13413
rect 10048 13268 10100 13320
rect 11612 13311 11664 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 2412 13243 2464 13252
rect 2412 13209 2421 13243
rect 2421 13209 2455 13243
rect 2455 13209 2464 13243
rect 2412 13200 2464 13209
rect 3700 13200 3752 13252
rect 8116 13200 8168 13252
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 14924 13268 14976 13320
rect 18052 13268 18104 13320
rect 13360 13200 13412 13252
rect 16028 13200 16080 13252
rect 16856 13200 16908 13252
rect 3240 13132 3292 13184
rect 9772 13132 9824 13184
rect 11244 13132 11296 13184
rect 12440 13132 12492 13184
rect 15752 13132 15804 13184
rect 18144 13132 18196 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2136 12928 2188 12980
rect 3056 12928 3108 12980
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 3700 12971 3752 12980
rect 3700 12937 3709 12971
rect 3709 12937 3743 12971
rect 3743 12937 3752 12971
rect 3700 12928 3752 12937
rect 6920 12928 6972 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 2964 12860 3016 12912
rect 6368 12860 6420 12912
rect 17776 12928 17828 12980
rect 9220 12903 9272 12912
rect 9220 12869 9238 12903
rect 9238 12869 9272 12903
rect 9220 12860 9272 12869
rect 9404 12860 9456 12912
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3792 12792 3844 12844
rect 6000 12792 6052 12844
rect 11612 12860 11664 12912
rect 8484 12724 8536 12776
rect 11152 12792 11204 12844
rect 11520 12792 11572 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 14924 12860 14976 12912
rect 2780 12656 2832 12708
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 2872 12588 2924 12597
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 8300 12588 8352 12640
rect 15568 12835 15620 12844
rect 15568 12801 15586 12835
rect 15586 12801 15620 12835
rect 15568 12792 15620 12801
rect 16580 12792 16632 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 13084 12588 13136 12640
rect 13176 12588 13228 12640
rect 16948 12656 17000 12708
rect 15844 12588 15896 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2044 12384 2096 12436
rect 2504 12384 2556 12436
rect 3424 12384 3476 12436
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 10324 12384 10376 12436
rect 9588 12316 9640 12368
rect 3056 12248 3108 12300
rect 3424 12248 3476 12300
rect 3976 12248 4028 12300
rect 8116 12248 8168 12300
rect 12072 12384 12124 12436
rect 15844 12384 15896 12436
rect 15660 12316 15712 12368
rect 18144 12384 18196 12436
rect 2872 12180 2924 12232
rect 4068 12180 4120 12232
rect 11060 12180 11112 12232
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 2872 12044 2924 12096
rect 4804 12112 4856 12164
rect 8760 12112 8812 12164
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 12808 12112 12860 12164
rect 12900 12112 12952 12164
rect 15752 12112 15804 12164
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 5816 12044 5868 12096
rect 11704 12044 11756 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12072 12044 12124 12096
rect 12532 12044 12584 12096
rect 14648 12044 14700 12096
rect 16120 12044 16172 12096
rect 16948 12112 17000 12164
rect 17040 12044 17092 12096
rect 17868 12044 17920 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2964 11840 3016 11892
rect 3424 11840 3476 11892
rect 7288 11840 7340 11892
rect 9588 11840 9640 11892
rect 15936 11840 15988 11892
rect 3056 11772 3108 11824
rect 3516 11772 3568 11824
rect 3608 11772 3660 11824
rect 11980 11772 12032 11824
rect 15660 11772 15712 11824
rect 16120 11772 16172 11824
rect 2688 11704 2740 11756
rect 3792 11704 3844 11756
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 2872 11636 2924 11688
rect 3884 11636 3936 11688
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4436 11636 4488 11688
rect 4896 11636 4948 11688
rect 6000 11636 6052 11688
rect 6276 11636 6328 11688
rect 3424 11568 3476 11620
rect 8024 11704 8076 11756
rect 8484 11704 8536 11756
rect 8944 11747 8996 11756
rect 8944 11713 8978 11747
rect 8978 11713 8996 11747
rect 8944 11704 8996 11713
rect 11060 11704 11112 11756
rect 11612 11704 11664 11756
rect 11796 11747 11848 11756
rect 11796 11713 11830 11747
rect 11830 11713 11848 11747
rect 11796 11704 11848 11713
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 10232 11636 10284 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 2320 11500 2372 11552
rect 2504 11500 2556 11552
rect 3884 11500 3936 11552
rect 4344 11500 4396 11552
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 4988 11500 5040 11509
rect 5172 11500 5224 11552
rect 9956 11500 10008 11552
rect 10968 11500 11020 11552
rect 11060 11500 11112 11552
rect 11520 11500 11572 11552
rect 11704 11500 11756 11552
rect 13820 11704 13872 11756
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 14096 11500 14148 11552
rect 15844 11500 15896 11552
rect 17132 11636 17184 11688
rect 17316 11500 17368 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 3056 11296 3108 11348
rect 3792 11296 3844 11348
rect 4988 11296 5040 11348
rect 1768 11228 1820 11280
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 2504 11228 2556 11280
rect 3056 11160 3108 11212
rect 3884 11228 3936 11280
rect 3608 11160 3660 11212
rect 4528 11228 4580 11280
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 2044 11024 2096 11076
rect 2596 11024 2648 11076
rect 3516 11092 3568 11144
rect 8852 11228 8904 11280
rect 9956 11296 10008 11348
rect 10324 11296 10376 11348
rect 11244 11296 11296 11348
rect 11520 11296 11572 11348
rect 15936 11296 15988 11348
rect 13820 11228 13872 11280
rect 8668 11092 8720 11144
rect 10232 11092 10284 11144
rect 12440 11092 12492 11144
rect 15844 11135 15896 11144
rect 4344 11024 4396 11076
rect 6368 11024 6420 11076
rect 8484 11024 8536 11076
rect 8760 11024 8812 11076
rect 9404 11024 9456 11076
rect 9772 11024 9824 11076
rect 12716 11024 12768 11076
rect 15200 11024 15252 11076
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 16856 11024 16908 11076
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 5724 10956 5776 11008
rect 6092 10999 6144 11008
rect 6092 10965 6101 10999
rect 6101 10965 6135 10999
rect 6135 10965 6144 10999
rect 6092 10956 6144 10965
rect 11060 10956 11112 11008
rect 12256 10999 12308 11008
rect 12256 10965 12265 10999
rect 12265 10965 12299 10999
rect 12299 10965 12308 10999
rect 12256 10956 12308 10965
rect 12532 10956 12584 11008
rect 16120 10956 16172 11008
rect 16580 10956 16632 11008
rect 17868 11024 17920 11076
rect 18788 11024 18840 11076
rect 19156 11024 19208 11076
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 3516 10795 3568 10804
rect 3516 10761 3525 10795
rect 3525 10761 3559 10795
rect 3559 10761 3568 10795
rect 3516 10752 3568 10761
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 8852 10752 8904 10804
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 2504 10684 2556 10736
rect 4528 10684 4580 10736
rect 8300 10727 8352 10736
rect 8300 10693 8334 10727
rect 8334 10693 8352 10727
rect 8300 10684 8352 10693
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2136 10591 2188 10600
rect 2136 10557 2145 10591
rect 2145 10557 2179 10591
rect 2179 10557 2188 10591
rect 2136 10548 2188 10557
rect 3608 10616 3660 10668
rect 4160 10616 4212 10668
rect 4252 10616 4304 10668
rect 6644 10616 6696 10668
rect 7104 10616 7156 10668
rect 11888 10752 11940 10804
rect 12256 10752 12308 10804
rect 13636 10752 13688 10804
rect 16580 10752 16632 10804
rect 10232 10684 10284 10736
rect 10876 10684 10928 10736
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 5724 10591 5776 10600
rect 4528 10480 4580 10532
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 5908 10480 5960 10532
rect 4712 10412 4764 10464
rect 5540 10412 5592 10464
rect 7380 10548 7432 10600
rect 9956 10548 10008 10600
rect 10508 10616 10560 10668
rect 11520 10616 11572 10668
rect 14556 10616 14608 10668
rect 15844 10684 15896 10736
rect 11428 10548 11480 10600
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 9220 10480 9272 10532
rect 6552 10412 6604 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 14188 10412 14240 10464
rect 17500 10412 17552 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 18512 10412 18564 10464
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 2228 10208 2280 10260
rect 2504 10208 2556 10260
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 1492 10140 1544 10192
rect 5724 10140 5776 10192
rect 2228 10072 2280 10124
rect 2504 10072 2556 10124
rect 2596 10072 2648 10124
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3976 10072 4028 10124
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 2136 10004 2188 10056
rect 1952 9936 2004 9988
rect 2688 9936 2740 9988
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 5172 10004 5224 10056
rect 6460 10140 6512 10192
rect 8852 10208 8904 10260
rect 11520 10208 11572 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13820 10208 13872 10260
rect 6828 10072 6880 10124
rect 9128 10140 9180 10192
rect 13728 10140 13780 10192
rect 14556 10183 14608 10192
rect 14556 10149 14565 10183
rect 14565 10149 14599 10183
rect 14599 10149 14608 10183
rect 14556 10140 14608 10149
rect 6552 10047 6604 10056
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 17776 10072 17828 10124
rect 8208 10004 8260 10056
rect 9680 10004 9732 10056
rect 10232 10004 10284 10056
rect 10416 10047 10468 10056
rect 10416 10013 10450 10047
rect 10450 10013 10468 10047
rect 10416 10004 10468 10013
rect 10876 10004 10928 10056
rect 15844 10004 15896 10056
rect 17868 10004 17920 10056
rect 7472 9936 7524 9988
rect 8024 9936 8076 9988
rect 10048 9936 10100 9988
rect 10692 9936 10744 9988
rect 15660 9979 15712 9988
rect 15660 9945 15678 9979
rect 15678 9945 15712 9979
rect 15660 9936 15712 9945
rect 17132 9979 17184 9988
rect 17132 9945 17150 9979
rect 17150 9945 17184 9979
rect 17132 9936 17184 9945
rect 2504 9868 2556 9877
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 8208 9868 8260 9920
rect 8668 9868 8720 9920
rect 9404 9868 9456 9920
rect 10232 9868 10284 9920
rect 11888 9868 11940 9920
rect 12808 9868 12860 9920
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 2688 9664 2740 9716
rect 3240 9664 3292 9716
rect 3976 9664 4028 9716
rect 4620 9664 4672 9716
rect 5724 9664 5776 9716
rect 7288 9664 7340 9716
rect 17868 9664 17920 9716
rect 3148 9596 3200 9648
rect 4252 9596 4304 9648
rect 5264 9596 5316 9648
rect 8392 9596 8444 9648
rect 2688 9528 2740 9580
rect 2780 9528 2832 9580
rect 3516 9528 3568 9580
rect 5172 9528 5224 9580
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6736 9571 6788 9580
rect 6184 9528 6236 9537
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7380 9528 7432 9580
rect 8024 9528 8076 9580
rect 2136 9460 2188 9512
rect 2872 9435 2924 9444
rect 1308 9324 1360 9376
rect 2872 9401 2881 9435
rect 2881 9401 2915 9435
rect 2915 9401 2924 9435
rect 2872 9392 2924 9401
rect 3700 9392 3752 9444
rect 3792 9392 3844 9444
rect 5816 9460 5868 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 5908 9392 5960 9444
rect 8116 9460 8168 9512
rect 9220 9528 9272 9580
rect 9772 9596 9824 9648
rect 10232 9596 10284 9648
rect 10692 9528 10744 9580
rect 9680 9460 9732 9512
rect 11796 9528 11848 9580
rect 12440 9596 12492 9648
rect 13912 9596 13964 9648
rect 14096 9528 14148 9580
rect 14740 9528 14792 9580
rect 15108 9596 15160 9648
rect 17408 9596 17460 9648
rect 17592 9528 17644 9580
rect 17684 9528 17736 9580
rect 4160 9324 4212 9376
rect 5080 9324 5132 9376
rect 9772 9392 9824 9444
rect 10140 9392 10192 9444
rect 8944 9324 8996 9376
rect 9036 9324 9088 9376
rect 10048 9324 10100 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 14188 9324 14240 9376
rect 18788 9392 18840 9444
rect 15660 9324 15712 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 18604 9324 18656 9376
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 3884 9120 3936 9172
rect 2964 9052 3016 9104
rect 5816 9120 5868 9172
rect 6828 9120 6880 9172
rect 8760 9163 8812 9172
rect 4068 9052 4120 9104
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 9588 9120 9640 9172
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 8944 9052 8996 9104
rect 2412 8984 2464 9036
rect 4712 8984 4764 9036
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 7012 8984 7064 9036
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 1860 8916 1912 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5632 8916 5684 8968
rect 2688 8848 2740 8900
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 2320 8780 2372 8832
rect 2872 8780 2924 8832
rect 3976 8848 4028 8900
rect 5172 8891 5224 8900
rect 5172 8857 5181 8891
rect 5181 8857 5215 8891
rect 5215 8857 5224 8891
rect 5172 8848 5224 8857
rect 6828 8848 6880 8900
rect 6920 8848 6972 8900
rect 8024 8916 8076 8968
rect 9680 8916 9732 8968
rect 8300 8848 8352 8900
rect 8484 8848 8536 8900
rect 13360 9120 13412 9172
rect 13452 9120 13504 9172
rect 15200 9120 15252 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 12992 8984 13044 9036
rect 13912 8984 13964 9036
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 11152 8916 11204 8968
rect 11888 8916 11940 8968
rect 3608 8780 3660 8832
rect 4436 8780 4488 8832
rect 4896 8780 4948 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 5816 8780 5868 8832
rect 7012 8780 7064 8832
rect 7196 8780 7248 8832
rect 11612 8848 11664 8900
rect 12256 8891 12308 8900
rect 12256 8857 12290 8891
rect 12290 8857 12308 8891
rect 12256 8848 12308 8857
rect 13360 8916 13412 8968
rect 14004 8916 14056 8968
rect 10232 8780 10284 8832
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 14280 8848 14332 8900
rect 15108 8916 15160 8968
rect 15384 8780 15436 8832
rect 17960 8780 18012 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 1492 8576 1544 8585
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 4160 8576 4212 8628
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5816 8576 5868 8628
rect 6368 8576 6420 8628
rect 8668 8576 8720 8628
rect 12256 8576 12308 8628
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 14556 8576 14608 8628
rect 16028 8576 16080 8628
rect 16396 8576 16448 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 1308 8508 1360 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2596 8440 2648 8492
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 2320 8372 2372 8424
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 1768 8236 1820 8288
rect 3608 8440 3660 8492
rect 3792 8415 3844 8424
rect 3792 8381 3801 8415
rect 3801 8381 3835 8415
rect 3835 8381 3844 8415
rect 3792 8372 3844 8381
rect 4160 8304 4212 8356
rect 4528 8304 4580 8356
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 5172 8440 5224 8492
rect 6828 8440 6880 8492
rect 8392 8508 8444 8560
rect 13084 8508 13136 8560
rect 14740 8508 14792 8560
rect 15016 8508 15068 8560
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 6920 8415 6972 8424
rect 5264 8372 5316 8381
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10508 8440 10560 8492
rect 10692 8440 10744 8492
rect 8116 8372 8168 8381
rect 5724 8304 5776 8356
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 6276 8304 6328 8356
rect 6368 8304 6420 8356
rect 7472 8304 7524 8356
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 4436 8236 4488 8288
rect 4988 8236 5040 8288
rect 5172 8236 5224 8288
rect 6828 8236 6880 8288
rect 9680 8236 9732 8288
rect 9864 8236 9916 8288
rect 11060 8440 11112 8492
rect 12440 8440 12492 8492
rect 14105 8483 14157 8492
rect 14105 8449 14139 8483
rect 14139 8449 14157 8483
rect 14105 8440 14157 8449
rect 15200 8440 15252 8492
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 12532 8415 12584 8424
rect 11060 8304 11112 8356
rect 11796 8304 11848 8356
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 16212 8372 16264 8424
rect 17868 8440 17920 8492
rect 16856 8372 16908 8424
rect 12992 8236 13044 8288
rect 14372 8236 14424 8288
rect 15568 8304 15620 8356
rect 17684 8372 17736 8424
rect 18144 8347 18196 8356
rect 18144 8313 18153 8347
rect 18153 8313 18187 8347
rect 18187 8313 18196 8347
rect 18144 8304 18196 8313
rect 15476 8236 15528 8288
rect 15660 8236 15712 8288
rect 17132 8236 17184 8288
rect 17868 8279 17920 8288
rect 17868 8245 17877 8279
rect 17877 8245 17911 8279
rect 17911 8245 17920 8279
rect 17868 8236 17920 8245
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 2688 8032 2740 8084
rect 2780 8032 2832 8084
rect 3240 8032 3292 8084
rect 3424 8032 3476 8084
rect 4068 8032 4120 8084
rect 5264 8032 5316 8084
rect 1492 7828 1544 7880
rect 2688 7896 2740 7948
rect 4160 7964 4212 8016
rect 2780 7828 2832 7880
rect 3700 7896 3752 7948
rect 4436 7828 4488 7880
rect 4988 7828 5040 7880
rect 5908 8032 5960 8084
rect 6736 8032 6788 8084
rect 8392 8032 8444 8084
rect 8484 7964 8536 8016
rect 8852 8032 8904 8084
rect 9680 8032 9732 8084
rect 11980 8032 12032 8084
rect 12440 8032 12492 8084
rect 11152 7964 11204 8016
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 6828 7896 6880 7948
rect 7840 7939 7892 7948
rect 1400 7692 1452 7744
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 3884 7803 3936 7812
rect 3884 7769 3893 7803
rect 3893 7769 3927 7803
rect 3927 7769 3936 7803
rect 3884 7760 3936 7769
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 8760 7896 8812 7948
rect 11244 7896 11296 7948
rect 11704 7896 11756 7948
rect 12072 7896 12124 7948
rect 14924 8032 14976 8084
rect 13544 7964 13596 8016
rect 14096 7964 14148 8016
rect 17592 8032 17644 8084
rect 17868 8032 17920 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 18236 7964 18288 8016
rect 13176 7939 13228 7948
rect 7380 7828 7432 7880
rect 2872 7692 2924 7744
rect 3516 7692 3568 7744
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 4896 7692 4948 7744
rect 5816 7735 5868 7744
rect 5816 7701 5825 7735
rect 5825 7701 5859 7735
rect 5859 7701 5868 7735
rect 5816 7692 5868 7701
rect 6184 7692 6236 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6644 7735 6696 7744
rect 6276 7692 6328 7701
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 6920 7692 6972 7744
rect 10232 7760 10284 7812
rect 7472 7692 7524 7744
rect 8116 7692 8168 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8944 7692 8996 7744
rect 9772 7692 9824 7744
rect 9864 7692 9916 7744
rect 10876 7828 10928 7880
rect 11428 7828 11480 7880
rect 11980 7828 12032 7880
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 12532 7828 12584 7880
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 12716 7760 12768 7812
rect 13636 7828 13688 7880
rect 14556 7896 14608 7948
rect 15292 7896 15344 7948
rect 16580 7896 16632 7948
rect 18052 7896 18104 7948
rect 18328 7896 18380 7948
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 15108 7828 15160 7880
rect 17132 7828 17184 7880
rect 17500 7828 17552 7880
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 16028 7760 16080 7812
rect 16120 7803 16172 7812
rect 16120 7769 16138 7803
rect 16138 7769 16172 7803
rect 16856 7803 16908 7812
rect 16120 7760 16172 7769
rect 16856 7769 16865 7803
rect 16865 7769 16899 7803
rect 16899 7769 16908 7803
rect 16856 7760 16908 7769
rect 17408 7760 17460 7812
rect 12624 7692 12676 7744
rect 13084 7692 13136 7744
rect 14740 7692 14792 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 15200 7692 15252 7744
rect 16396 7692 16448 7744
rect 16948 7692 17000 7744
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 17776 7735 17828 7744
rect 17776 7701 17785 7735
rect 17785 7701 17819 7735
rect 17819 7701 17828 7735
rect 17776 7692 17828 7701
rect 18512 7692 18564 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 1952 7488 2004 7540
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 1584 7420 1636 7472
rect 2688 7420 2740 7472
rect 3884 7488 3936 7540
rect 5264 7488 5316 7540
rect 5816 7488 5868 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 2504 7352 2556 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 2044 7284 2096 7336
rect 2780 7284 2832 7336
rect 3608 7352 3660 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 3056 7216 3108 7268
rect 4344 7352 4396 7404
rect 5264 7352 5316 7404
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 6736 7420 6788 7472
rect 6552 7352 6604 7404
rect 4068 7284 4120 7293
rect 5816 7216 5868 7268
rect 7564 7352 7616 7404
rect 7932 7488 7984 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8300 7488 8352 7540
rect 9496 7488 9548 7540
rect 11152 7488 11204 7540
rect 13084 7531 13136 7540
rect 13084 7497 13093 7531
rect 13093 7497 13127 7531
rect 13127 7497 13136 7531
rect 13084 7488 13136 7497
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 18236 7488 18288 7540
rect 12624 7463 12676 7472
rect 8852 7352 8904 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10416 7352 10468 7404
rect 7196 7216 7248 7268
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 9404 7327 9456 7336
rect 8760 7284 8812 7293
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 8392 7216 8444 7268
rect 10508 7284 10560 7336
rect 11428 7284 11480 7336
rect 11888 7284 11940 7336
rect 10600 7216 10652 7268
rect 12624 7429 12633 7463
rect 12633 7429 12667 7463
rect 12667 7429 12676 7463
rect 12624 7420 12676 7429
rect 13544 7420 13596 7472
rect 13820 7420 13872 7472
rect 14556 7420 14608 7472
rect 16672 7420 16724 7472
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13360 7284 13412 7336
rect 13636 7284 13688 7336
rect 14188 7284 14240 7336
rect 15200 7284 15252 7336
rect 16580 7352 16632 7404
rect 17408 7352 17460 7404
rect 17592 7352 17644 7404
rect 14740 7216 14792 7268
rect 14924 7216 14976 7268
rect 16764 7284 16816 7336
rect 18328 7352 18380 7404
rect 4988 7148 5040 7200
rect 5724 7148 5776 7200
rect 6552 7148 6604 7200
rect 6828 7148 6880 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 12072 7148 12124 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 13636 7148 13688 7200
rect 14464 7148 14516 7200
rect 15844 7148 15896 7200
rect 16488 7216 16540 7268
rect 16672 7259 16724 7268
rect 16672 7225 16681 7259
rect 16681 7225 16715 7259
rect 16715 7225 16724 7259
rect 16672 7216 16724 7225
rect 16948 7216 17000 7268
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1584 6944 1636 6996
rect 2136 6944 2188 6996
rect 3424 6944 3476 6996
rect 3608 6944 3660 6996
rect 5264 6944 5316 6996
rect 7472 6944 7524 6996
rect 8392 6944 8444 6996
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 10232 6944 10284 6996
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 12440 6944 12492 6996
rect 2044 6808 2096 6860
rect 3148 6808 3200 6860
rect 3976 6808 4028 6860
rect 5080 6808 5132 6860
rect 5908 6808 5960 6860
rect 2872 6740 2924 6792
rect 3516 6740 3568 6792
rect 3608 6740 3660 6792
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 8760 6876 8812 6928
rect 6644 6740 6696 6792
rect 2044 6672 2096 6724
rect 2964 6672 3016 6724
rect 6828 6672 6880 6724
rect 8024 6740 8076 6792
rect 9312 6808 9364 6860
rect 9588 6876 9640 6928
rect 12164 6876 12216 6928
rect 9680 6808 9732 6860
rect 10324 6808 10376 6860
rect 11244 6808 11296 6860
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 12900 6808 12952 6860
rect 15016 6876 15068 6928
rect 16028 6944 16080 6996
rect 16948 6944 17000 6996
rect 18144 6876 18196 6928
rect 18328 6876 18380 6928
rect 9772 6740 9824 6792
rect 9312 6672 9364 6724
rect 11152 6740 11204 6792
rect 11428 6740 11480 6792
rect 11888 6740 11940 6792
rect 13544 6740 13596 6792
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 14464 6851 14516 6860
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 14832 6808 14884 6860
rect 14004 6740 14056 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 15752 6808 15804 6860
rect 17132 6808 17184 6860
rect 15936 6740 15988 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 16672 6740 16724 6792
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 2320 6647 2372 6656
rect 1952 6604 2004 6613
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2780 6604 2832 6656
rect 3516 6604 3568 6656
rect 3792 6604 3844 6656
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4160 6604 4212 6656
rect 4620 6604 4672 6656
rect 5356 6604 5408 6656
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 6184 6647 6236 6656
rect 6184 6613 6193 6647
rect 6193 6613 6227 6647
rect 6227 6613 6236 6647
rect 6184 6604 6236 6613
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9128 6604 9180 6656
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 12900 6672 12952 6724
rect 13176 6672 13228 6724
rect 11888 6604 11940 6613
rect 12624 6604 12676 6656
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13084 6604 13136 6613
rect 13636 6604 13688 6656
rect 14832 6604 14884 6656
rect 15200 6604 15252 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 16488 6604 16540 6656
rect 16948 6604 17000 6656
rect 17316 6672 17368 6724
rect 18144 6740 18196 6792
rect 18328 6740 18380 6792
rect 19248 6740 19300 6792
rect 17868 6715 17920 6724
rect 17868 6681 17877 6715
rect 17877 6681 17911 6715
rect 17911 6681 17920 6715
rect 17868 6672 17920 6681
rect 18788 6672 18840 6724
rect 17776 6604 17828 6656
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 2964 6400 3016 6452
rect 3516 6400 3568 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 4712 6400 4764 6452
rect 6368 6400 6420 6452
rect 2228 6332 2280 6384
rect 5908 6332 5960 6384
rect 6552 6332 6604 6384
rect 6736 6400 6788 6452
rect 8024 6400 8076 6452
rect 8852 6400 8904 6452
rect 9312 6400 9364 6452
rect 9588 6400 9640 6452
rect 10324 6400 10376 6452
rect 10508 6400 10560 6452
rect 10600 6400 10652 6452
rect 12808 6400 12860 6452
rect 14096 6400 14148 6452
rect 15016 6400 15068 6452
rect 15200 6443 15252 6452
rect 15200 6409 15209 6443
rect 15209 6409 15243 6443
rect 15243 6409 15252 6443
rect 15200 6400 15252 6409
rect 17592 6400 17644 6452
rect 8760 6375 8812 6384
rect 1952 6264 2004 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3608 6264 3660 6316
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 2964 6128 3016 6180
rect 5632 6264 5684 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7104 6264 7156 6316
rect 7288 6264 7340 6316
rect 5080 6196 5132 6248
rect 5264 6196 5316 6248
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6460 6239 6512 6248
rect 6000 6196 6052 6205
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 7748 6239 7800 6248
rect 7012 6128 7064 6180
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 7196 6060 7248 6112
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 8760 6341 8769 6375
rect 8769 6341 8803 6375
rect 8803 6341 8812 6375
rect 8760 6332 8812 6341
rect 8944 6264 8996 6316
rect 11428 6332 11480 6384
rect 11796 6332 11848 6384
rect 8208 6196 8260 6248
rect 8576 6196 8628 6248
rect 9772 6264 9824 6316
rect 9956 6196 10008 6248
rect 10232 6264 10284 6316
rect 11704 6264 11756 6316
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11428 6196 11480 6248
rect 12164 6332 12216 6384
rect 15844 6332 15896 6384
rect 16764 6332 16816 6384
rect 19340 6400 19392 6452
rect 12900 6264 12952 6316
rect 12624 6196 12676 6248
rect 13268 6264 13320 6316
rect 15936 6264 15988 6316
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 14096 6196 14148 6248
rect 8024 6128 8076 6180
rect 9864 6128 9916 6180
rect 10416 6128 10468 6180
rect 11152 6128 11204 6180
rect 14188 6128 14240 6180
rect 15292 6196 15344 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16672 6196 16724 6248
rect 17776 6264 17828 6316
rect 18328 6264 18380 6316
rect 14924 6128 14976 6180
rect 17132 6128 17184 6180
rect 17408 6171 17460 6180
rect 17408 6137 17417 6171
rect 17417 6137 17451 6171
rect 17451 6137 17460 6171
rect 17408 6128 17460 6137
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 10232 6060 10284 6112
rect 12532 6060 12584 6112
rect 14740 6060 14792 6112
rect 15108 6060 15160 6112
rect 15660 6060 15712 6112
rect 15752 6060 15804 6112
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 2504 5856 2556 5908
rect 2872 5856 2924 5908
rect 3608 5856 3660 5908
rect 3884 5899 3936 5908
rect 3884 5865 3893 5899
rect 3893 5865 3927 5899
rect 3927 5865 3936 5899
rect 3884 5856 3936 5865
rect 4528 5899 4580 5908
rect 4528 5865 4537 5899
rect 4537 5865 4571 5899
rect 4571 5865 4580 5899
rect 4528 5856 4580 5865
rect 5264 5856 5316 5908
rect 6736 5856 6788 5908
rect 6828 5856 6880 5908
rect 9956 5899 10008 5908
rect 2320 5788 2372 5840
rect 2596 5720 2648 5772
rect 4620 5788 4672 5840
rect 1492 5652 1544 5704
rect 2044 5652 2096 5704
rect 1308 5584 1360 5636
rect 2136 5584 2188 5636
rect 3976 5584 4028 5636
rect 1952 5516 2004 5568
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3516 5516 3568 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 5172 5720 5224 5772
rect 5816 5788 5868 5840
rect 5448 5763 5500 5772
rect 5448 5729 5457 5763
rect 5457 5729 5491 5763
rect 5491 5729 5500 5763
rect 5448 5720 5500 5729
rect 6000 5720 6052 5772
rect 6460 5720 6512 5772
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6828 5652 6880 5704
rect 8668 5788 8720 5840
rect 7196 5720 7248 5772
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 11888 5856 11940 5908
rect 13820 5899 13872 5908
rect 13820 5865 13829 5899
rect 13829 5865 13863 5899
rect 13863 5865 13872 5899
rect 13820 5856 13872 5865
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 15384 5856 15436 5908
rect 16120 5856 16172 5908
rect 17408 5856 17460 5908
rect 17868 5856 17920 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 8944 5763 8996 5772
rect 8944 5729 8953 5763
rect 8953 5729 8987 5763
rect 8987 5729 8996 5763
rect 8944 5720 8996 5729
rect 11244 5788 11296 5840
rect 13268 5788 13320 5840
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 12440 5652 12492 5704
rect 12808 5652 12860 5704
rect 13728 5720 13780 5772
rect 14924 5720 14976 5772
rect 15936 5788 15988 5840
rect 17224 5788 17276 5840
rect 17316 5788 17368 5840
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 16396 5720 16448 5772
rect 6736 5584 6788 5636
rect 5724 5516 5776 5568
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 7656 5584 7708 5636
rect 7840 5584 7892 5636
rect 10324 5584 10376 5636
rect 6000 5516 6052 5525
rect 7564 5516 7616 5568
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 9864 5516 9916 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 10508 5559 10560 5568
rect 10508 5525 10517 5559
rect 10517 5525 10551 5559
rect 10551 5525 10560 5559
rect 10876 5559 10928 5568
rect 10508 5516 10560 5525
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 11704 5584 11756 5636
rect 11796 5516 11848 5568
rect 11980 5516 12032 5568
rect 12348 5516 12400 5568
rect 12532 5516 12584 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 14096 5516 14148 5568
rect 14924 5516 14976 5568
rect 17040 5652 17092 5704
rect 15200 5516 15252 5568
rect 15660 5559 15712 5568
rect 15660 5525 15669 5559
rect 15669 5525 15703 5559
rect 15703 5525 15712 5559
rect 15660 5516 15712 5525
rect 16028 5516 16080 5568
rect 17224 5559 17276 5568
rect 17224 5525 17233 5559
rect 17233 5525 17267 5559
rect 17267 5525 17276 5559
rect 17224 5516 17276 5525
rect 17316 5516 17368 5568
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18604 5652 18656 5704
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 2412 5312 2464 5364
rect 4068 5355 4120 5364
rect 2228 5244 2280 5296
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 6000 5312 6052 5364
rect 6644 5312 6696 5364
rect 7196 5312 7248 5364
rect 3332 5287 3384 5296
rect 3332 5253 3341 5287
rect 3341 5253 3375 5287
rect 3375 5253 3384 5287
rect 3332 5244 3384 5253
rect 5724 5244 5776 5296
rect 6460 5287 6512 5296
rect 6460 5253 6469 5287
rect 6469 5253 6503 5287
rect 6503 5253 6512 5287
rect 6460 5244 6512 5253
rect 2780 5176 2832 5185
rect 3332 5108 3384 5160
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 2780 5040 2832 5092
rect 5816 5176 5868 5228
rect 7012 5176 7064 5228
rect 7748 5312 7800 5364
rect 8300 5312 8352 5364
rect 9588 5312 9640 5364
rect 10232 5312 10284 5364
rect 10876 5355 10928 5364
rect 10876 5321 10885 5355
rect 10885 5321 10919 5355
rect 10919 5321 10928 5355
rect 10876 5312 10928 5321
rect 11428 5312 11480 5364
rect 13268 5312 13320 5364
rect 7656 5176 7708 5228
rect 8024 5176 8076 5228
rect 10508 5244 10560 5296
rect 10968 5244 11020 5296
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 15108 5312 15160 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 16212 5312 16264 5364
rect 17224 5312 17276 5364
rect 18788 5312 18840 5364
rect 19156 5312 19208 5364
rect 5632 5108 5684 5160
rect 6644 5108 6696 5160
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7472 5108 7524 5160
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2872 4972 2924 5024
rect 4712 4972 4764 5024
rect 9680 5176 9732 5228
rect 10232 5176 10284 5228
rect 10324 5176 10376 5228
rect 11796 5176 11848 5228
rect 14280 5244 14332 5296
rect 9864 5108 9916 5160
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 10600 5040 10652 5092
rect 12440 5108 12492 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 13452 5108 13504 5160
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 11888 5040 11940 5092
rect 12256 5040 12308 5092
rect 12532 5040 12584 5092
rect 13360 5040 13412 5092
rect 13912 5176 13964 5228
rect 14556 5176 14608 5228
rect 16120 5244 16172 5296
rect 16856 5244 16908 5296
rect 17132 5244 17184 5296
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 14096 5108 14148 5160
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 14648 5108 14700 5160
rect 15292 5108 15344 5160
rect 15752 5151 15804 5160
rect 15200 5040 15252 5092
rect 15476 5040 15528 5092
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 16948 5108 17000 5160
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 9864 4972 9916 5024
rect 10416 4972 10468 5024
rect 10508 4972 10560 5024
rect 15108 4972 15160 5024
rect 16120 4972 16172 5024
rect 16396 4972 16448 5024
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 2136 4768 2188 4820
rect 2780 4768 2832 4820
rect 3884 4768 3936 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 8760 4811 8812 4820
rect 5264 4700 5316 4752
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 2780 4564 2832 4573
rect 4804 4564 4856 4616
rect 5908 4632 5960 4684
rect 6368 4700 6420 4752
rect 7104 4700 7156 4752
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 9036 4768 9088 4820
rect 9404 4768 9456 4820
rect 9496 4768 9548 4820
rect 11336 4768 11388 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 12624 4768 12676 4820
rect 13176 4768 13228 4820
rect 13820 4768 13872 4820
rect 6460 4632 6512 4684
rect 7380 4632 7432 4684
rect 14556 4700 14608 4752
rect 10140 4632 10192 4684
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10600 4632 10652 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 12808 4632 12860 4684
rect 12900 4632 12952 4684
rect 14464 4632 14516 4684
rect 15476 4768 15528 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 18512 4768 18564 4820
rect 15108 4700 15160 4752
rect 18696 4700 18748 4752
rect 16304 4675 16356 4684
rect 16304 4641 16313 4675
rect 16313 4641 16347 4675
rect 16347 4641 16356 4675
rect 16304 4632 16356 4641
rect 17960 4632 18012 4684
rect 6644 4564 6696 4616
rect 8760 4564 8812 4616
rect 9312 4564 9364 4616
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9680 4564 9732 4616
rect 10876 4564 10928 4616
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 15844 4564 15896 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16580 4564 16632 4616
rect 17592 4564 17644 4616
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 2964 4496 3016 4548
rect 5264 4539 5316 4548
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 4620 4428 4672 4480
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 6184 4428 6236 4480
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7380 4428 7432 4480
rect 11980 4496 12032 4548
rect 9312 4428 9364 4480
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 10876 4428 10928 4480
rect 10968 4428 11020 4480
rect 11704 4428 11756 4480
rect 13268 4428 13320 4480
rect 14188 4496 14240 4548
rect 15016 4496 15068 4548
rect 15200 4428 15252 4480
rect 17224 4496 17276 4548
rect 17960 4496 18012 4548
rect 16764 4428 16816 4480
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 5816 4224 5868 4276
rect 6460 4224 6512 4276
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 7380 4267 7432 4276
rect 7380 4233 7389 4267
rect 7389 4233 7423 4267
rect 7423 4233 7432 4267
rect 7380 4224 7432 4233
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 8300 4267 8352 4276
rect 7472 4224 7524 4233
rect 8300 4233 8309 4267
rect 8309 4233 8343 4267
rect 8343 4233 8352 4267
rect 8300 4224 8352 4233
rect 1952 4156 2004 4208
rect 2136 4088 2188 4140
rect 2688 4088 2740 4140
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 5908 4156 5960 4208
rect 7196 4156 7248 4208
rect 8484 4224 8536 4276
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 9588 4224 9640 4276
rect 10508 4224 10560 4276
rect 11796 4224 11848 4276
rect 12532 4224 12584 4276
rect 6000 4088 6052 4140
rect 10416 4156 10468 4208
rect 11520 4131 11572 4140
rect 3700 4020 3752 4072
rect 8208 4020 8260 4072
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 11612 4020 11664 4072
rect 11980 4020 12032 4072
rect 13728 4267 13780 4276
rect 13728 4233 13737 4267
rect 13737 4233 13771 4267
rect 13771 4233 13780 4267
rect 14096 4267 14148 4276
rect 13728 4224 13780 4233
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 14924 4224 14976 4276
rect 15108 4224 15160 4276
rect 15936 4267 15988 4276
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 17408 4224 17460 4276
rect 14004 4088 14056 4140
rect 16856 4156 16908 4208
rect 17040 4156 17092 4208
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 13544 4063 13596 4072
rect 12808 4020 12860 4029
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 2780 3995 2832 4004
rect 2780 3961 2789 3995
rect 2789 3961 2823 3995
rect 2823 3961 2832 3995
rect 2780 3952 2832 3961
rect 7104 3952 7156 4004
rect 10232 3995 10284 4004
rect 10232 3961 10241 3995
rect 10241 3961 10275 3995
rect 10275 3961 10284 3995
rect 10232 3952 10284 3961
rect 2872 3884 2924 3936
rect 8024 3884 8076 3936
rect 9496 3884 9548 3936
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 11244 3884 11296 3936
rect 13912 3952 13964 4004
rect 15016 4020 15068 4072
rect 15660 4088 15712 4140
rect 16396 4088 16448 4140
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 16304 4020 16356 4072
rect 14648 3884 14700 3936
rect 16028 3952 16080 4004
rect 16764 3952 16816 4004
rect 17040 3952 17092 4004
rect 17224 4088 17276 4140
rect 17684 4088 17736 4140
rect 17868 4020 17920 4072
rect 19064 4020 19116 4072
rect 18144 3995 18196 4004
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 15476 3884 15528 3936
rect 15936 3884 15988 3936
rect 16856 3884 16908 3936
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 1952 3476 2004 3528
rect 8208 3680 8260 3732
rect 8760 3723 8812 3732
rect 8760 3689 8769 3723
rect 8769 3689 8803 3723
rect 8803 3689 8812 3723
rect 8760 3680 8812 3689
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 10324 3680 10376 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 13728 3680 13780 3732
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 14556 3723 14608 3732
rect 14556 3689 14565 3723
rect 14565 3689 14599 3723
rect 14599 3689 14608 3723
rect 14556 3680 14608 3689
rect 15016 3680 15068 3732
rect 15200 3680 15252 3732
rect 15292 3723 15344 3732
rect 15292 3689 15301 3723
rect 15301 3689 15335 3723
rect 15335 3689 15344 3723
rect 15660 3723 15712 3732
rect 15292 3680 15344 3689
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16396 3680 16448 3732
rect 16948 3723 17000 3732
rect 16948 3689 16957 3723
rect 16957 3689 16991 3723
rect 16991 3689 17000 3723
rect 16948 3680 17000 3689
rect 17316 3723 17368 3732
rect 17316 3689 17325 3723
rect 17325 3689 17359 3723
rect 17359 3689 17368 3723
rect 17316 3680 17368 3689
rect 18236 3723 18288 3732
rect 18236 3689 18245 3723
rect 18245 3689 18279 3723
rect 18279 3689 18288 3723
rect 18236 3680 18288 3689
rect 19248 3680 19300 3732
rect 12808 3612 12860 3664
rect 8668 3544 8720 3596
rect 15108 3544 15160 3596
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 17224 3612 17276 3664
rect 15568 3544 15620 3596
rect 16028 3544 16080 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 16396 3544 16448 3596
rect 17500 3612 17552 3664
rect 3700 3408 3752 3460
rect 6092 3476 6144 3528
rect 7012 3476 7064 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 10784 3476 10836 3528
rect 13084 3476 13136 3528
rect 14004 3476 14056 3528
rect 15016 3476 15068 3528
rect 16212 3476 16264 3528
rect 18972 3544 19024 3596
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 18052 3519 18104 3528
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 2780 3340 2832 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 8024 3408 8076 3460
rect 9496 3408 9548 3460
rect 12808 3408 12860 3460
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 4896 3340 4948 3392
rect 9680 3340 9732 3392
rect 15568 3340 15620 3392
rect 15752 3340 15804 3392
rect 16488 3340 16540 3392
rect 17776 3340 17828 3392
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16212 3136 16264 3145
rect 17040 3136 17092 3188
rect 17408 3136 17460 3188
rect 18328 3136 18380 3188
rect 6184 3068 6236 3120
rect 11152 3068 11204 3120
rect 2320 3000 2372 3052
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 6644 3000 6696 3052
rect 3700 2932 3752 2984
rect 4528 2932 4580 2984
rect 6276 2932 6328 2984
rect 7288 3000 7340 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 7012 2864 7064 2916
rect 10324 2864 10376 2916
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 11888 3000 11940 3052
rect 14648 3068 14700 3120
rect 14924 3068 14976 3120
rect 15660 3068 15712 3120
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 15384 3043 15436 3052
rect 14832 3000 14884 3009
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 16580 3068 16632 3120
rect 17684 3068 17736 3120
rect 17960 3068 18012 3120
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 18144 3000 18196 3052
rect 18420 3000 18472 3052
rect 13636 2932 13688 2984
rect 14648 2932 14700 2984
rect 17684 2932 17736 2984
rect 18604 2932 18656 2984
rect 15568 2864 15620 2916
rect 18144 2864 18196 2916
rect 15292 2796 15344 2848
rect 16488 2796 16540 2848
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 17868 2592 17920 2644
rect 18512 2592 18564 2644
rect 16672 2524 16724 2576
rect 17040 2567 17092 2576
rect 17040 2533 17049 2567
rect 17049 2533 17083 2567
rect 17083 2533 17092 2567
rect 17040 2524 17092 2533
rect 17224 2567 17276 2576
rect 17224 2533 17233 2567
rect 17233 2533 17267 2567
rect 17267 2533 17276 2567
rect 17224 2524 17276 2533
rect 17960 2524 18012 2576
rect 18144 2524 18196 2576
rect 19340 2524 19392 2576
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 4252 2388 4304 2440
rect 18052 2456 18104 2508
rect 8208 2320 8260 2372
rect 16580 2388 16632 2440
rect 16672 2388 16724 2440
rect 17316 2388 17368 2440
rect 17868 2431 17920 2440
rect 17592 2320 17644 2372
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18696 2320 18748 2372
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 16580 2252 16632 2304
rect 16856 2252 16908 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 4988 1776 5040 1828
rect 16028 1776 16080 1828
<< metal2 >>
rect 2042 16538 2098 17200
rect 2042 16510 2636 16538
rect 2042 16400 2098 16510
rect 2134 14376 2190 14385
rect 2134 14311 2190 14320
rect 1582 14104 1638 14113
rect 1582 14039 1638 14048
rect 1596 13394 1624 14039
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13569 1900 13806
rect 1858 13560 1914 13569
rect 1858 13495 1914 13504
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2148 13326 2176 14311
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2136 13320 2188 13326
rect 1858 13288 1914 13297
rect 2136 13262 2188 13268
rect 1858 13223 1860 13232
rect 1912 13223 1914 13232
rect 1860 13194 1912 13200
rect 2148 12986 2176 13262
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12442 2084 12786
rect 2044 12436 2096 12442
rect 2332 12434 2360 14214
rect 2412 13864 2464 13870
rect 2410 13832 2412 13841
rect 2464 13832 2466 13841
rect 2410 13767 2466 13776
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2424 13025 2452 13194
rect 2410 13016 2466 13025
rect 2410 12951 2466 12960
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 12753 2544 12786
rect 2502 12744 2558 12753
rect 2502 12679 2558 12688
rect 2516 12442 2544 12679
rect 2608 12458 2636 16510
rect 5998 16400 6054 17200
rect 9954 16538 10010 17200
rect 9784 16510 10010 16538
rect 2870 15464 2926 15473
rect 2870 15399 2926 15408
rect 2778 15192 2834 15201
rect 2778 15127 2834 15136
rect 2792 14618 2820 15127
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2792 13954 2820 14554
rect 2700 13938 2820 13954
rect 2688 13932 2820 13938
rect 2740 13926 2820 13932
rect 2688 13874 2740 13880
rect 2884 13870 2912 15399
rect 3054 14920 3110 14929
rect 3054 14855 3110 14864
rect 2962 14648 3018 14657
rect 2962 14583 3018 14592
rect 2976 14385 3004 14583
rect 2962 14376 3018 14385
rect 2962 14311 3018 14320
rect 2964 14000 3016 14006
rect 3068 13988 3096 14855
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 3016 13960 3096 13988
rect 2964 13942 3016 13948
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3620 13705 3648 13806
rect 3606 13696 3662 13705
rect 3174 13628 3482 13637
rect 3606 13631 3662 13640
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 6012 13433 6040 16400
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 5998 13424 6054 13433
rect 3516 13388 3568 13394
rect 5998 13359 6054 13368
rect 3516 13330 3568 13336
rect 2688 13320 2740 13326
rect 2686 13288 2688 13297
rect 2740 13288 2742 13297
rect 2686 13223 2742 13232
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 12986 3280 13126
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12481 2820 12650
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2778 12472 2834 12481
rect 2504 12436 2556 12442
rect 2332 12406 2452 12434
rect 2044 12378 2096 12384
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 11393 1808 11494
rect 1766 11384 1822 11393
rect 1766 11319 1822 11328
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1320 8566 1348 9318
rect 1504 8634 1532 10134
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1320 7313 1348 8502
rect 1504 7886 1532 8570
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 1306 7032 1362 7041
rect 1306 6967 1362 6976
rect 1320 6633 1348 6967
rect 1306 6624 1362 6633
rect 1306 6559 1362 6568
rect 1320 5642 1348 6559
rect 1308 5636 1360 5642
rect 1308 5578 1360 5584
rect 1412 4865 1440 7686
rect 1596 7478 1624 9687
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1596 7002 1624 7414
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1688 6848 1716 8774
rect 1780 8430 1808 11222
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 8974 1900 10950
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1860 8968 1912 8974
rect 1964 8945 1992 9930
rect 1860 8910 1912 8916
rect 1950 8936 2006 8945
rect 1950 8871 2006 8880
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 7546 1808 8230
rect 1964 7546 1992 8434
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2056 7342 2084 11018
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2148 10062 2176 10542
rect 2240 10266 2268 12038
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11218 2360 11494
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 10441 2360 10610
rect 2318 10432 2374 10441
rect 2318 10367 2374 10376
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9518 2176 9998
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2240 9330 2268 10066
rect 2148 9302 2268 9330
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2056 6866 2084 7278
rect 2148 7002 2176 9302
rect 2424 9042 2452 12406
rect 2608 12430 2728 12458
rect 2504 12378 2556 12384
rect 2700 12322 2728 12430
rect 2778 12407 2834 12416
rect 2700 12294 2820 12322
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11286 2544 11494
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2608 11082 2636 11630
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2700 10810 2728 11698
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2516 10266 2544 10678
rect 2594 10568 2650 10577
rect 2594 10503 2650 10512
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2516 10130 2544 10202
rect 2608 10130 2636 10503
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2594 9888 2650 9897
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2044 6860 2096 6866
rect 1688 6820 1808 6848
rect 1674 6760 1730 6769
rect 1674 6695 1730 6704
rect 1688 6458 1716 6695
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 1596 5914 1624 6151
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1504 5370 1532 5646
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1780 4622 1808 6820
rect 2044 6802 2096 6808
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1872 5914 1900 6598
rect 1964 6458 1992 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1950 6352 2006 6361
rect 1950 6287 1952 6296
rect 2004 6287 2006 6296
rect 1952 6258 2004 6264
rect 2056 6225 2084 6666
rect 2240 6390 2268 7686
rect 2332 6662 2360 8366
rect 2410 7576 2466 7585
rect 2410 7511 2466 7520
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2424 6458 2452 7511
rect 2516 7410 2544 9862
rect 2594 9823 2650 9832
rect 2608 8498 2636 9823
rect 2700 9722 2728 9930
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2792 9586 2820 12294
rect 2884 12238 2912 12582
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11778 2912 12038
rect 2976 11898 3004 12854
rect 3068 12306 3096 12922
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 3424 12436 3476 12442
rect 3528 12434 3556 13330
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3476 12406 3556 12434
rect 3620 12434 3648 13262
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3712 12986 3740 13194
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 3804 12442 3832 12786
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3792 12436 3844 12442
rect 3620 12406 3740 12434
rect 3424 12378 3476 12384
rect 3436 12306 3464 12378
rect 3514 12336 3570 12345
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3424 12300 3476 12306
rect 3514 12271 3570 12280
rect 3424 12242 3476 12248
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3056 11824 3108 11830
rect 2884 11750 3004 11778
rect 3056 11766 3108 11772
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2700 8906 2728 9522
rect 2792 9178 2820 9522
rect 2884 9450 2912 11630
rect 2976 10713 3004 11750
rect 3068 11354 3096 11766
rect 3436 11626 3464 11834
rect 3528 11830 3556 12271
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3620 11218 3648 11766
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 2962 10704 3018 10713
rect 2962 10639 3018 10648
rect 2962 10432 3018 10441
rect 2962 10367 3018 10376
rect 2976 10130 3004 10367
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2962 9752 3018 9761
rect 2962 9687 3018 9696
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2976 9330 3004 9687
rect 2884 9302 3004 9330
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 9058 2912 9302
rect 2962 9208 3018 9217
rect 2962 9143 3018 9152
rect 2976 9110 3004 9143
rect 2792 9030 2912 9058
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2686 8800 2742 8809
rect 2686 8735 2742 8744
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2042 6216 2098 6225
rect 2042 6151 2098 6160
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2056 5710 2084 6151
rect 2332 5846 2360 6258
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2044 5704 2096 5710
rect 1858 5672 1914 5681
rect 2044 5646 2096 5652
rect 1858 5607 1914 5616
rect 2136 5636 2188 5642
rect 1872 5370 1900 5607
rect 2136 5578 2188 5584
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1858 4584 1914 4593
rect 1858 4519 1914 4528
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1214 3088 1270 3097
rect 1214 3023 1270 3032
rect 1228 800 1256 3023
rect 1504 2689 1532 4422
rect 1872 4010 1900 4519
rect 1964 4214 1992 5510
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2056 5001 2084 5170
rect 2042 4992 2098 5001
rect 2042 4927 2098 4936
rect 2148 4826 2176 5578
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 5302 2268 5510
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2240 4321 2268 4966
rect 2226 4312 2282 4321
rect 2226 4247 2282 4256
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1964 3534 1992 4150
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2042 3904 2098 3913
rect 2042 3839 2098 3848
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1490 2680 1546 2689
rect 1490 2615 1546 2624
rect 1688 1601 1716 3334
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 2145 1900 2790
rect 1858 2136 1914 2145
rect 1858 2071 1914 2080
rect 1674 1592 1730 1601
rect 1674 1527 1730 1536
rect 2056 800 2084 3839
rect 2148 3641 2176 4082
rect 2134 3632 2190 3641
rect 2134 3567 2190 3576
rect 2332 3058 2360 5782
rect 2424 5370 2452 6394
rect 2516 5914 2544 7346
rect 2608 6254 2636 8434
rect 2700 8090 2728 8735
rect 2792 8090 2820 9030
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8498 2912 8774
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2884 8129 2912 8434
rect 2962 8392 3018 8401
rect 2962 8327 3018 8336
rect 2870 8120 2926 8129
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2780 8084 2832 8090
rect 2870 8055 2926 8064
rect 2780 8026 2832 8032
rect 2686 7984 2742 7993
rect 2686 7919 2688 7928
rect 2740 7919 2742 7928
rect 2688 7890 2740 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 5778 2636 6190
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2410 3768 2466 3777
rect 2410 3703 2412 3712
rect 2464 3703 2466 3712
rect 2412 3674 2464 3680
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2608 2417 2636 4422
rect 2700 4146 2728 7414
rect 2792 7342 2820 7822
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7546 2912 7686
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2870 7440 2926 7449
rect 2870 7375 2926 7384
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2884 6798 2912 7375
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 5953 2820 6598
rect 2778 5944 2834 5953
rect 2884 5914 2912 6734
rect 2976 6730 3004 8327
rect 3068 7449 3096 11154
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 10810 3556 11086
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3514 10704 3570 10713
rect 3514 10639 3570 10648
rect 3608 10668 3660 10674
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3528 9761 3556 10639
rect 3608 10610 3660 10616
rect 3514 9752 3570 9761
rect 3240 9716 3292 9722
rect 3160 9664 3240 9674
rect 3514 9687 3570 9696
rect 3160 9658 3292 9664
rect 3160 9654 3280 9658
rect 3148 9648 3280 9654
rect 3200 9646 3280 9648
rect 3148 9590 3200 9596
rect 3516 9580 3568 9586
rect 3620 9568 3648 10610
rect 3712 9625 3740 12406
rect 3792 12378 3844 12384
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 11665 3832 11698
rect 3884 11688 3936 11694
rect 3790 11656 3846 11665
rect 3988 11676 4016 12242
rect 4080 12238 4108 12582
rect 4068 12232 4120 12238
rect 4066 12200 4068 12209
rect 4120 12200 4122 12209
rect 4066 12135 4122 12144
rect 4710 12200 4766 12209
rect 4710 12135 4766 12144
rect 4804 12164 4856 12170
rect 4080 12109 4108 12135
rect 4724 12102 4752 12135
rect 4804 12106 4856 12112
rect 4712 12096 4764 12102
rect 4632 12056 4712 12084
rect 4158 11792 4214 11801
rect 4158 11727 4214 11736
rect 3936 11648 4016 11676
rect 3884 11630 3936 11636
rect 3790 11591 3846 11600
rect 3804 11354 3832 11591
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11286 3924 11494
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3988 10713 4016 11648
rect 4068 11688 4120 11694
rect 4172 11676 4200 11727
rect 4120 11648 4200 11676
rect 4436 11688 4488 11694
rect 4068 11630 4120 11636
rect 4436 11630 4488 11636
rect 4344 11552 4396 11558
rect 4066 11520 4122 11529
rect 4344 11494 4396 11500
rect 4066 11455 4122 11464
rect 4080 11064 4108 11455
rect 4356 11218 4384 11494
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4344 11076 4396 11082
rect 4080 11036 4292 11064
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3568 9540 3648 9568
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3516 9522 3568 9528
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3054 7440 3110 7449
rect 3252 7410 3280 8026
rect 3436 7993 3464 8026
rect 3422 7984 3478 7993
rect 3422 7919 3478 7928
rect 3528 7936 3556 9522
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8498 3648 8774
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3712 8401 3740 9386
rect 3804 8430 3832 9386
rect 3896 9178 3924 10542
rect 3976 10124 4028 10130
rect 4080 10112 4108 10775
rect 4264 10674 4292 11036
rect 4344 11018 4396 11024
rect 4356 10810 4384 11018
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4172 10266 4200 10610
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4080 10084 4200 10112
rect 3976 10066 4028 10072
rect 3988 9722 4016 10066
rect 4066 10024 4122 10033
rect 4066 9959 4068 9968
rect 4120 9959 4122 9968
rect 4068 9930 4120 9936
rect 4172 9874 4200 10084
rect 4080 9846 4200 9874
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3882 9072 3938 9081
rect 3882 9007 3938 9016
rect 3792 8424 3844 8430
rect 3698 8392 3754 8401
rect 3792 8366 3844 8372
rect 3698 8327 3754 8336
rect 3700 7948 3752 7954
rect 3528 7908 3700 7936
rect 3528 7857 3556 7908
rect 3896 7936 3924 9007
rect 3988 8906 4016 9658
rect 4080 9217 4108 9846
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4066 9208 4122 9217
rect 4066 9143 4122 9152
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3700 7890 3752 7896
rect 3804 7908 3924 7936
rect 3514 7848 3570 7857
rect 3514 7783 3570 7792
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3054 7375 3110 7384
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 7313 3280 7346
rect 3238 7304 3294 7313
rect 3056 7268 3108 7274
rect 3238 7239 3294 7248
rect 3056 7210 3108 7216
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6458 3004 6666
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2962 6352 3018 6361
rect 2962 6287 3018 6296
rect 2976 6186 3004 6287
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2778 5879 2834 5888
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2778 5264 2834 5273
rect 2834 5222 2912 5250
rect 2778 5199 2780 5208
rect 2832 5199 2834 5208
rect 2780 5170 2832 5176
rect 2778 5128 2834 5137
rect 2778 5063 2780 5072
rect 2832 5063 2834 5072
rect 2780 5034 2832 5040
rect 2884 5030 2912 5222
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2792 4622 2820 4762
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2778 4040 2834 4049
rect 2778 3975 2780 3984
rect 2832 3975 2834 3984
rect 2780 3946 2832 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2594 2408 2650 2417
rect 2594 2343 2650 2352
rect 2792 1873 2820 3334
rect 2884 2961 2912 3878
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2976 2258 3004 4490
rect 3068 3505 3096 7210
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3146 6896 3202 6905
rect 3146 6831 3148 6840
rect 3200 6831 3202 6840
rect 3148 6802 3200 6808
rect 3436 6338 3464 6938
rect 3528 6798 3556 7686
rect 3606 7576 3662 7585
rect 3606 7511 3662 7520
rect 3620 7410 3648 7511
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3606 7168 3662 7177
rect 3606 7103 3662 7112
rect 3620 7002 3648 7103
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6458 3556 6598
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3436 6310 3556 6338
rect 3620 6322 3648 6734
rect 3712 6322 3740 7890
rect 3804 7041 3832 7908
rect 3882 7848 3938 7857
rect 3882 7783 3884 7792
rect 3936 7783 3938 7792
rect 3884 7754 3936 7760
rect 3896 7546 3924 7754
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3884 7336 3936 7342
rect 3882 7304 3884 7313
rect 3936 7304 3938 7313
rect 3882 7239 3938 7248
rect 3790 7032 3846 7041
rect 3790 6967 3846 6976
rect 3882 6896 3938 6905
rect 3988 6866 4016 8842
rect 4080 8673 4108 9046
rect 4172 8974 4200 9318
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4066 8664 4122 8673
rect 4066 8599 4122 8608
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4172 8537 4200 8570
rect 4158 8528 4214 8537
rect 4158 8463 4214 8472
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 8106 4200 8298
rect 4080 8090 4200 8106
rect 4068 8084 4200 8090
rect 4120 8078 4200 8084
rect 4068 8026 4120 8032
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7342 4108 7686
rect 4068 7336 4120 7342
rect 4172 7313 4200 7958
rect 4068 7278 4120 7284
rect 4158 7304 4214 7313
rect 3882 6831 3938 6840
rect 3976 6860 4028 6866
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3528 5574 3556 6310
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3620 5914 3648 6258
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3332 5296 3384 5302
rect 3330 5264 3332 5273
rect 3384 5264 3386 5273
rect 3330 5199 3386 5208
rect 3344 5166 3372 5199
rect 3332 5160 3384 5166
rect 3424 5160 3476 5166
rect 3332 5102 3384 5108
rect 3422 5128 3424 5137
rect 3476 5128 3478 5137
rect 3422 5063 3478 5072
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 3146 4584 3202 4593
rect 3146 4519 3202 4528
rect 3160 4146 3188 4519
rect 3528 4185 3556 5510
rect 3514 4176 3570 4185
rect 3148 4140 3200 4146
rect 3514 4111 3570 4120
rect 3148 4082 3200 4088
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3054 3496 3110 3505
rect 3712 3466 3740 4014
rect 3054 3431 3110 3440
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3804 3058 3832 6598
rect 3896 5914 3924 6831
rect 3976 6802 4028 6808
rect 3988 6662 4016 6802
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3988 5658 4016 6598
rect 3896 5642 4016 5658
rect 3896 5636 4028 5642
rect 3896 5630 3976 5636
rect 3896 4826 3924 5630
rect 3976 5578 4028 5584
rect 4080 5522 4108 7278
rect 4158 7239 4214 7248
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6458 4200 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3988 5494 4108 5522
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3988 4593 4016 5494
rect 4066 5400 4122 5409
rect 4066 5335 4068 5344
rect 4120 5335 4122 5344
rect 4068 5306 4120 5312
rect 3974 4584 4030 4593
rect 3974 4519 4030 4528
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3233 3924 3334
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 2884 2230 3004 2258
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 2884 800 2912 2230
rect 3712 800 3740 2926
rect 4264 2446 4292 9590
rect 4448 8945 4476 11630
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4540 10742 4568 11222
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4540 10538 4568 10678
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4632 10010 4660 12056
rect 4712 12038 4764 12044
rect 4710 11792 4766 11801
rect 4710 11727 4766 11736
rect 4724 10470 4752 11727
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 10130 4752 10406
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4540 9982 4660 10010
rect 4434 8936 4490 8945
rect 4434 8871 4490 8880
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8634 4476 8774
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4342 8392 4398 8401
rect 4540 8362 4568 9982
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9722 4660 9862
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4618 9480 4674 9489
rect 4618 9415 4674 9424
rect 4342 8327 4398 8336
rect 4528 8356 4580 8362
rect 4356 7410 4384 8327
rect 4528 8298 4580 8304
rect 4436 8288 4488 8294
rect 4488 8236 4568 8242
rect 4436 8230 4568 8236
rect 4448 8214 4568 8230
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4448 6254 4476 7822
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4540 5914 4568 8214
rect 4632 6662 4660 9415
rect 4724 9042 4752 10066
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4632 5846 4660 6598
rect 4724 6458 4752 8298
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4632 4486 4660 5782
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5030 4752 5510
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4816 4622 4844 12106
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 4896 11688 4948 11694
rect 4894 11656 4896 11665
rect 4948 11656 4950 11665
rect 4894 11591 4950 11600
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5000 11354 5028 11494
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 7750 4936 8774
rect 5000 8401 5028 11290
rect 5184 10062 5212 11494
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 5736 10606 5764 10950
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10130 5580 10406
rect 5736 10198 5764 10542
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9586 5212 9998
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 5736 9722 5764 9862
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5092 8809 5120 9318
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5078 8800 5134 8809
rect 5078 8735 5134 8744
rect 5184 8634 5212 8842
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5172 8492 5224 8498
rect 5092 8452 5172 8480
rect 4986 8392 5042 8401
rect 4986 8327 5042 8336
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 7886 5028 8230
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 5000 7562 5028 7822
rect 5092 7585 5120 8452
rect 5172 8434 5224 8440
rect 5276 8430 5304 9590
rect 5828 9518 5856 12038
rect 6012 11694 6040 12786
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6196 11098 6224 13874
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6012 11070 6224 11098
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5920 9450 5948 10474
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8838 5672 8910
rect 5828 8838 5856 9114
rect 5906 9072 5962 9081
rect 5906 9007 5908 9016
rect 5960 9007 5962 9016
rect 5908 8978 5960 8984
rect 5632 8832 5684 8838
rect 5816 8832 5868 8838
rect 5684 8792 5764 8820
rect 5632 8774 5684 8780
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5736 8362 5764 8792
rect 5816 8774 5868 8780
rect 5828 8634 5856 8774
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 4908 7534 5028 7562
rect 5078 7576 5134 7585
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4908 3398 4936 7534
rect 5078 7511 5134 7520
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 5681 5028 7142
rect 5092 6866 5120 7511
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 6254 5120 6802
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5184 5778 5212 8230
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5276 7546 5304 8026
rect 5828 7834 5856 8570
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5920 8090 5948 8298
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5736 7806 5856 7834
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 7002 5304 7346
rect 5736 7206 5764 7806
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7546 5856 7686
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5828 6662 5856 7210
rect 5920 6866 5948 8026
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5356 6656 5408 6662
rect 5276 6633 5356 6644
rect 5262 6624 5356 6633
rect 5318 6616 5356 6624
rect 5356 6598 5408 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5262 6559 5318 6568
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5828 6497 5856 6598
rect 5814 6488 5870 6497
rect 5814 6423 5870 6432
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5914 5304 6190
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4986 5672 5042 5681
rect 4986 5607 5042 5616
rect 5000 5370 5028 5607
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4540 800 4568 2926
rect 5000 1834 5028 5306
rect 5276 4758 5304 5850
rect 5460 5778 5488 6054
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5540 5704 5592 5710
rect 5538 5672 5540 5681
rect 5592 5672 5594 5681
rect 5538 5607 5594 5616
rect 5644 5556 5672 6258
rect 5828 5930 5856 6423
rect 5920 6390 5948 6802
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6012 6254 6040 11070
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6288 10962 6316 11630
rect 6380 11082 6408 12854
rect 6734 11248 6790 11257
rect 6734 11183 6790 11192
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5828 5902 5948 5930
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5724 5568 5776 5574
rect 5644 5528 5724 5556
rect 5724 5510 5776 5516
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5736 5302 5764 5510
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5828 5234 5856 5782
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4826 5672 5102
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5276 1986 5304 4490
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5828 4282 5856 5170
rect 5920 4690 5948 5902
rect 6012 5778 6040 6190
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5370 6040 5510
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5920 4214 5948 4626
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 6012 4146 6040 4422
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6104 3534 6132 10950
rect 6288 10934 6408 10962
rect 6182 10160 6238 10169
rect 6182 10095 6238 10104
rect 6196 9586 6224 10095
rect 6380 10010 6408 10934
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6288 9982 6408 10010
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6196 8537 6224 9415
rect 6182 8528 6238 8537
rect 6182 8463 6238 8472
rect 6196 7834 6224 8463
rect 6288 8362 6316 9982
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6380 8362 6408 8570
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6196 7806 6408 7834
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6182 7168 6238 7177
rect 6182 7103 6238 7112
rect 6196 6662 6224 7103
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 4486 6224 6598
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5276 1958 5396 1986
rect 4988 1828 5040 1834
rect 4988 1770 5040 1776
rect 5368 800 5396 1958
rect 6196 800 6224 3062
rect 6288 2990 6316 7686
rect 6380 6458 6408 7806
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6380 4758 6408 6394
rect 6472 6361 6500 10134
rect 6564 10062 6592 10406
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6550 8936 6606 8945
rect 6550 8871 6606 8880
rect 6564 7954 6592 8871
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6656 7834 6684 10610
rect 6748 10033 6776 11183
rect 6840 10130 6868 14758
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 14006 7420 14350
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 7380 14000 7432 14006
rect 6918 13968 6974 13977
rect 7380 13942 7432 13948
rect 6918 13903 6974 13912
rect 6932 13530 6960 13903
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7392 13394 7420 13942
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6932 12434 6960 12922
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 6932 12406 7236 12434
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6828 10124 6880 10130
rect 6880 10084 6960 10112
rect 6828 10066 6880 10072
rect 6734 10024 6790 10033
rect 6734 9959 6790 9968
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 8537 6776 9522
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9178 6868 9454
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 8906 6960 10084
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6840 8809 6868 8842
rect 7024 8838 7052 8978
rect 7012 8832 7064 8838
rect 6826 8800 6882 8809
rect 7012 8774 7064 8780
rect 6826 8735 6882 8744
rect 6734 8528 6790 8537
rect 6734 8463 6790 8472
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6840 8294 6868 8434
rect 6920 8424 6972 8430
rect 7024 8412 7052 8774
rect 6972 8384 7052 8412
rect 6920 8366 6972 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6564 7806 6684 7834
rect 6564 7546 6592 7806
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6564 7313 6592 7346
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6390 6592 7142
rect 6656 6798 6684 7686
rect 6748 7478 6776 8026
rect 6840 7954 6868 8230
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6840 7206 6868 7890
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6458 6776 6598
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6552 6384 6604 6390
rect 6458 6352 6514 6361
rect 6552 6326 6604 6332
rect 6458 6287 6514 6296
rect 6736 6316 6788 6322
rect 6472 6254 6500 6287
rect 6736 6258 6788 6264
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6472 5302 6500 5714
rect 6656 5370 6684 6190
rect 6748 5914 6776 6258
rect 6840 5914 6868 6666
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6828 5704 6880 5710
rect 6734 5672 6790 5681
rect 6828 5646 6880 5652
rect 6734 5607 6736 5616
rect 6788 5607 6790 5616
rect 6736 5578 6788 5584
rect 6840 5545 6868 5646
rect 6826 5536 6882 5545
rect 6826 5471 6882 5480
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6472 4690 6500 5238
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 4282 6500 4626
rect 6656 4622 6684 5102
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6656 3058 6684 4422
rect 6932 3516 6960 7686
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 7024 6186 7052 7239
rect 7116 6662 7144 10610
rect 7208 9194 7236 12406
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7300 9722 7328 11834
rect 8036 11762 8064 13466
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8128 12986 8156 13194
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 8022 11112 8078 11121
rect 8022 11047 8078 11056
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 10062 7420 10542
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7392 9586 7420 9998
rect 8036 9994 8064 11047
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7208 9166 7328 9194
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7208 7274 7236 8774
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7194 7032 7250 7041
rect 7194 6967 7250 6976
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7024 4729 7052 5170
rect 7116 5166 7144 6258
rect 7208 6202 7236 6967
rect 7300 6322 7328 9166
rect 7392 9042 7420 9522
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7484 8362 7512 9930
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 8036 8974 8064 9522
rect 8128 9518 8156 12242
rect 8220 10062 8248 14282
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8496 13734 8524 13874
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8312 10742 8340 12582
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8404 10577 8432 13670
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 11762 8524 12718
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8390 10568 8446 10577
rect 8390 10503 8446 10512
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8128 8430 8156 9454
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 7838 7984 7894 7993
rect 7838 7919 7840 7928
rect 7892 7919 7894 7928
rect 7840 7890 7892 7896
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 6882 7420 7822
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7002 7512 7686
rect 7562 7576 7618 7585
rect 8036 7562 8064 8366
rect 8128 8129 8156 8366
rect 8114 8120 8170 8129
rect 8114 8055 8170 8064
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7944 7546 8064 7562
rect 8128 7546 8156 7686
rect 7562 7511 7618 7520
rect 7932 7540 8064 7546
rect 7576 7410 7604 7511
rect 7984 7534 8064 7540
rect 8116 7540 8168 7546
rect 7932 7482 7984 7488
rect 8116 7482 8168 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7392 6854 7512 6882
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7208 6174 7328 6202
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 5778 7236 6054
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7300 5522 7328 6174
rect 7208 5494 7328 5522
rect 7208 5370 7236 5494
rect 7286 5400 7342 5409
rect 7196 5364 7248 5370
rect 7286 5335 7342 5344
rect 7196 5306 7248 5312
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4758 7144 5102
rect 7104 4752 7156 4758
rect 7010 4720 7066 4729
rect 7104 4694 7156 4700
rect 7010 4655 7066 4664
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7024 4282 7052 4422
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7116 4010 7144 4422
rect 7208 4214 7236 5306
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7012 3528 7064 3534
rect 6932 3488 7012 3516
rect 7012 3470 7064 3476
rect 7300 3058 7328 5335
rect 7484 5250 7512 6854
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 6633 7788 6802
rect 8036 6798 8064 7278
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8220 6712 8248 9862
rect 8404 9654 8432 10503
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8496 9500 8524 11018
rect 8312 9472 8524 9500
rect 8312 8906 8340 9472
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8312 7868 8340 8842
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8404 8090 8432 8502
rect 8496 8362 8524 8842
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8496 8022 8524 8298
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8312 7840 8524 7868
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 7002 8432 7210
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8128 6684 8248 6712
rect 7746 6624 7802 6633
rect 7746 6559 7802 6568
rect 8022 6488 8078 6497
rect 8022 6423 8024 6432
rect 8076 6423 8078 6432
rect 8024 6394 8076 6400
rect 7748 6248 7800 6254
rect 7746 6216 7748 6225
rect 7800 6216 7802 6225
rect 7746 6151 7802 6160
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 8036 5658 8064 6122
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7944 5630 8064 5658
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7576 5409 7604 5510
rect 7562 5400 7618 5409
rect 7562 5335 7618 5344
rect 7668 5352 7696 5578
rect 7748 5364 7800 5370
rect 7668 5324 7748 5352
rect 7748 5306 7800 5312
rect 7852 5250 7880 5578
rect 7392 5222 7512 5250
rect 7668 5234 7880 5250
rect 7656 5228 7880 5234
rect 7392 4690 7420 5222
rect 7708 5222 7880 5228
rect 7656 5170 7708 5176
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4282 7420 4422
rect 7484 4282 7512 5102
rect 7944 5080 7972 5630
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5234 8064 5510
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7944 5052 8064 5080
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 8036 3942 8064 5052
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 8128 3534 8156 6684
rect 8390 6352 8446 6361
rect 8390 6287 8446 6296
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 5250 8248 6190
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5370 8340 6054
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8220 5222 8340 5250
rect 8206 4720 8262 4729
rect 8206 4655 8262 4664
rect 8220 4078 8248 4655
rect 8312 4282 8340 5222
rect 8404 5166 8432 6287
rect 8496 5574 8524 7840
rect 8588 6254 8616 14894
rect 9232 14414 9260 14962
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13938 8892 14214
rect 9324 14006 9352 14350
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9312 14000 9364 14006
rect 9588 14000 9640 14006
rect 9364 13960 9444 13988
rect 9312 13942 9364 13948
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13841 8892 13874
rect 8850 13832 8906 13841
rect 8850 13767 8906 13776
rect 9218 13288 9274 13297
rect 9218 13223 9274 13232
rect 9232 12918 9260 13223
rect 9416 12918 9444 13960
rect 9588 13942 9640 13948
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11150 8708 11630
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8772 11082 8800 12106
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8864 10810 8892 11222
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8850 10432 8906 10441
rect 8850 10367 8906 10376
rect 8864 10266 8892 10367
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8758 10024 8814 10033
rect 8758 9959 8814 9968
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 8634 8708 9862
rect 8772 9178 8800 9959
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8588 5778 8616 6190
rect 8680 5846 8708 8570
rect 8864 8090 8892 10202
rect 8956 9382 8984 11698
rect 9416 11082 9444 12854
rect 9600 12374 9628 13942
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11898 9628 12310
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9692 10962 9720 14214
rect 9784 14074 9812 16510
rect 9954 16400 10010 16510
rect 13910 16538 13966 17200
rect 17866 16538 17922 17200
rect 13910 16510 14320 16538
rect 13910 16400 13966 16510
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10060 14346 10088 14826
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 10244 14074 10272 14214
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9876 13308 9904 13466
rect 10048 13320 10100 13326
rect 9876 13280 10048 13308
rect 10048 13262 10100 13268
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 11082 9812 13126
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 10336 12442 10364 14962
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11354 9996 11494
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10244 11150 10272 11630
rect 10336 11354 10364 12378
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9692 10934 9812 10962
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9218 10704 9274 10713
rect 9218 10639 9274 10648
rect 9232 10538 9260 10639
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 7342 8800 7890
rect 8956 7834 8984 9046
rect 9048 8809 9076 9318
rect 9034 8800 9090 8809
rect 9034 8735 9090 8744
rect 8956 7806 9076 7834
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 7336 8812 7342
rect 8864 7313 8892 7346
rect 8760 7278 8812 7284
rect 8850 7304 8906 7313
rect 8772 6934 8800 7278
rect 8850 7239 8906 7248
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8864 6458 8892 7239
rect 8956 6905 8984 7686
rect 8942 6896 8998 6905
rect 8942 6831 8998 6840
rect 8942 6760 8998 6769
rect 8942 6695 8998 6704
rect 8956 6662 8984 6695
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8760 6384 8812 6390
rect 8758 6352 8760 6361
rect 8812 6352 8814 6361
rect 8758 6287 8814 6296
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8496 4282 8524 5510
rect 8772 4826 8800 6287
rect 8864 5273 8892 6394
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5778 8984 6258
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8850 5264 8906 5273
rect 8850 5199 8906 5208
rect 9048 4826 9076 7806
rect 9140 6662 9168 10134
rect 9232 9586 9260 10474
rect 9416 9926 9444 10746
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9692 9518 9720 9998
rect 9784 9654 9812 10934
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 10244 10742 10272 11086
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10470 9996 10542
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 10060 9994 10088 10095
rect 10244 10062 10272 10678
rect 10428 10062 10456 14554
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10520 12434 10548 14282
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11426 13424 11482 13433
rect 11426 13359 11482 13368
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10520 12406 10640 12434
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10232 9920 10284 9926
rect 10230 9888 10232 9897
rect 10284 9888 10286 9897
rect 9846 9820 10154 9829
rect 10230 9823 10286 9832
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 10138 9688 10194 9697
rect 9772 9648 9824 9654
rect 10138 9623 10194 9632
rect 10232 9648 10284 9654
rect 9772 9590 9824 9596
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 7002 9352 7346
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6730 9352 6802
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9416 6497 9444 7278
rect 9508 6916 9536 7482
rect 9600 7342 9628 9114
rect 9692 8974 9720 9454
rect 10152 9450 10180 9623
rect 10232 9590 10284 9596
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8294 9720 8910
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9588 6928 9640 6934
rect 9508 6888 9588 6916
rect 9588 6870 9640 6876
rect 9402 6488 9458 6497
rect 9312 6452 9364 6458
rect 9600 6458 9628 6870
rect 9692 6866 9720 8026
rect 9784 7750 9812 9386
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9217 10088 9318
rect 10046 9208 10102 9217
rect 10046 9143 10102 9152
rect 10244 8922 10272 9590
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10336 9178 10364 9415
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10244 8894 10364 8922
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9876 8294 9904 8434
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7750 9904 8230
rect 10244 7818 10272 8774
rect 10336 7993 10364 8894
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9784 6798 9812 7142
rect 9772 6792 9824 6798
rect 10152 6769 10180 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9772 6734 9824 6740
rect 10138 6760 10194 6769
rect 10138 6695 10194 6704
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 9402 6423 9458 6432
rect 9588 6452 9640 6458
rect 9312 6394 9364 6400
rect 9324 5545 9352 6394
rect 9416 6304 9444 6423
rect 9588 6394 9640 6400
rect 10244 6322 10272 6938
rect 10336 6866 10364 7919
rect 10428 7562 10456 9998
rect 10520 8498 10548 10610
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10428 7534 10548 7562
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6458 10364 6598
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 9772 6316 9824 6322
rect 9416 6276 9772 6304
rect 9772 6258 9824 6264
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9496 5568 9548 5574
rect 9310 5536 9366 5545
rect 9496 5510 9548 5516
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9310 5471 9366 5480
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8772 4622 8800 4762
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3738 8248 4014
rect 8772 3738 8800 4558
rect 9048 3913 9076 4762
rect 9324 4622 9352 5471
rect 9508 4826 9536 5510
rect 9600 5370 9628 5510
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9692 5234 9720 5607
rect 9784 5273 9812 6258
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9876 5574 9904 6122
rect 9968 5914 9996 6190
rect 10428 6186 10456 7346
rect 10520 7342 10548 7534
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10520 6458 10548 7278
rect 10612 7274 10640 12406
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9897 10732 9930
rect 10690 9888 10746 9897
rect 10690 9823 10746 9832
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 8498 10732 9522
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10690 7984 10746 7993
rect 10690 7919 10746 7928
rect 10704 7449 10732 7919
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 10244 5370 10272 6054
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 9770 5264 9826 5273
rect 9680 5228 9732 5234
rect 10336 5234 10364 5578
rect 10416 5568 10468 5574
rect 10414 5536 10416 5545
rect 10508 5568 10560 5574
rect 10468 5536 10470 5545
rect 10508 5510 10560 5516
rect 10414 5471 10470 5480
rect 9770 5199 9826 5208
rect 10232 5228 10284 5234
rect 9680 5170 9732 5176
rect 10232 5170 10284 5176
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 9876 5030 9904 5102
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9416 4486 9444 4762
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9508 3942 9536 4558
rect 9600 4282 9628 4966
rect 10152 4690 10180 5102
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9496 3936 9548 3942
rect 9034 3904 9090 3913
rect 9496 3878 9548 3884
rect 9034 3839 9090 3848
rect 9048 3738 9076 3839
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7024 800 7052 2858
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 8036 1714 8064 3402
rect 8220 2378 8248 3674
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 7852 1686 8064 1714
rect 7852 800 7880 1686
rect 8680 800 8708 3538
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9508 800 9536 3402
rect 9692 3398 9720 4558
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 10244 4010 10272 5170
rect 10336 4729 10364 5170
rect 10428 5030 10456 5471
rect 10520 5302 10548 5510
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10520 5030 10548 5238
rect 10612 5098 10640 6394
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10322 4720 10378 4729
rect 10322 4655 10324 4664
rect 10376 4655 10378 4664
rect 10324 4626 10376 4632
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10336 3738 10364 4626
rect 10428 4214 10456 4966
rect 10520 4282 10548 4966
rect 10612 4690 10640 5034
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10704 4593 10732 6598
rect 10796 6254 10824 13223
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11762 11100 12174
rect 11164 11801 11192 12786
rect 11150 11792 11206 11801
rect 11060 11756 11112 11762
rect 11150 11727 11206 11736
rect 11060 11698 11112 11704
rect 10968 11552 11020 11558
rect 11060 11552 11112 11558
rect 10968 11494 11020 11500
rect 11058 11520 11060 11529
rect 11112 11520 11114 11529
rect 11256 11506 11284 13126
rect 11440 12434 11468 13359
rect 11532 12850 11560 14214
rect 11624 14074 11652 14758
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 12636 13938 12664 14894
rect 12900 14544 12952 14550
rect 12820 14492 12900 14498
rect 12820 14486 12952 14492
rect 12820 14470 12940 14486
rect 12820 14006 12848 14470
rect 13096 14414 13124 14894
rect 14292 14618 14320 16510
rect 17604 16510 17922 16538
rect 15014 15056 15070 15065
rect 15014 14991 15070 15000
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 12992 14408 13044 14414
rect 12912 14356 12992 14362
rect 12912 14350 13044 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12912 14334 13032 14350
rect 13452 14340 13504 14346
rect 12912 14006 12940 14334
rect 13452 14282 13504 14288
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12912 13870 12940 13942
rect 12900 13864 12952 13870
rect 11702 13832 11758 13841
rect 12900 13806 12952 13812
rect 11702 13767 11758 13776
rect 11716 13462 11744 13767
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12918 11652 13262
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10888 10062 10916 10678
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10874 9344 10930 9353
rect 10874 9279 10930 9288
rect 10888 8537 10916 9279
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10888 6100 10916 7822
rect 10796 6072 10916 6100
rect 10796 5137 10824 6072
rect 10980 5681 11008 11494
rect 11058 11455 11114 11464
rect 11164 11478 11284 11506
rect 11348 12406 11468 12434
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 8498 11100 10950
rect 11164 8974 11192 11478
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10888 5370 10916 5510
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10980 5302 11008 5510
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10782 5128 10838 5137
rect 10782 5063 10838 5072
rect 11072 4622 11100 8298
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11164 7546 11192 7958
rect 11256 7954 11284 11290
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11256 6866 11284 7890
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11164 6361 11192 6734
rect 11150 6352 11206 6361
rect 11150 6287 11206 6296
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11164 4690 11192 6122
rect 11256 5846 11284 6802
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11256 4690 11284 5607
rect 11348 4826 11376 12406
rect 11624 12238 11652 12854
rect 11612 12232 11664 12238
rect 11532 12180 11612 12186
rect 11532 12174 11664 12180
rect 11532 12158 11652 12174
rect 11532 11694 11560 12158
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11354 11560 11494
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10600 11480 10606
rect 11426 10568 11428 10577
rect 11480 10568 11482 10577
rect 11426 10503 11482 10512
rect 11532 10266 11560 10610
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11426 10160 11482 10169
rect 11426 10095 11482 10104
rect 11440 7886 11468 10095
rect 11624 9674 11652 11698
rect 11716 11558 11744 12038
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11704 11552 11756 11558
rect 11808 11529 11836 11698
rect 11704 11494 11756 11500
rect 11794 11520 11850 11529
rect 11794 11455 11850 11464
rect 11900 10810 11928 13670
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 12072 12436 12124 12442
rect 12452 12434 12480 13126
rect 12912 12850 12940 13806
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 13188 12646 13216 13466
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12452 12406 12572 12434
rect 12072 12378 12124 12384
rect 12084 12102 12112 12378
rect 12544 12102 12572 12406
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 11992 11830 12020 12038
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10810 12296 10950
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11624 9646 11744 9674
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11440 7002 11468 7278
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 6390 11468 6734
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11440 5370 11468 6190
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 10876 4616 10928 4622
rect 10690 4584 10746 4593
rect 11060 4616 11112 4622
rect 10928 4576 11008 4604
rect 10876 4558 10928 4564
rect 10690 4519 10746 4528
rect 10980 4486 11008 4576
rect 11060 4558 11112 4564
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3777 10548 3878
rect 10506 3768 10562 3777
rect 10324 3732 10376 3738
rect 10796 3738 10824 3975
rect 10506 3703 10562 3712
rect 10784 3732 10836 3738
rect 10324 3674 10376 3680
rect 10784 3674 10836 3680
rect 10796 3534 10824 3674
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 10888 3058 10916 4422
rect 11256 3942 11284 4626
rect 11532 4146 11560 7142
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11624 4078 11652 8842
rect 11716 7954 11744 9646
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9042 11836 9522
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11900 8974 11928 9862
rect 12452 9654 12480 11086
rect 12544 11014 12572 12038
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11702 7712 11758 7721
rect 11702 7647 11758 7656
rect 11716 7177 11744 7647
rect 11702 7168 11758 7177
rect 11702 7103 11758 7112
rect 11808 6390 11836 8298
rect 11900 7342 11928 8910
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8634 12296 8842
rect 12728 8634 12756 11018
rect 12820 9926 12848 12106
rect 12912 11558 12940 12106
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11257 12940 11494
rect 12898 11248 12954 11257
rect 12898 11183 12954 11192
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 8090 12020 8366
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12452 8090 12480 8434
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11888 6792 11940 6798
rect 11992 6780 12020 7822
rect 12084 7750 12112 7890
rect 12544 7886 12572 8366
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12084 7206 12112 7686
rect 12636 7478 12664 7686
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 12452 7002 12480 7142
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 11940 6752 12020 6780
rect 11888 6734 11940 6740
rect 11888 6656 11940 6662
rect 11886 6624 11888 6633
rect 11940 6624 11942 6633
rect 11886 6559 11942 6568
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11716 5642 11744 6258
rect 11900 5914 11928 6258
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11886 5808 11942 5817
rect 11886 5743 11942 5752
rect 11900 5710 11928 5743
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11992 5574 12020 6752
rect 12176 6390 12204 6870
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6497 12664 6598
rect 12622 6488 12678 6497
rect 12622 6423 12678 6432
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 12544 5778 12572 6054
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12530 5672 12586 5681
rect 11796 5568 11848 5574
rect 11716 5516 11796 5522
rect 11716 5510 11848 5516
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 11716 5494 11836 5510
rect 11716 4486 11744 5494
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11808 4282 11836 5170
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11992 5080 12020 5238
rect 12256 5092 12308 5098
rect 11992 5052 12256 5080
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 10336 800 10364 2858
rect 11164 800 11192 3062
rect 11900 3058 11928 5034
rect 11992 4554 12020 5052
rect 12256 5034 12308 5040
rect 12360 5012 12388 5510
rect 12452 5166 12480 5646
rect 12530 5607 12586 5616
rect 12544 5574 12572 5607
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12636 5250 12664 6190
rect 12728 5778 12756 7754
rect 12820 6866 12848 9862
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 13004 9042 13032 9551
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13004 8378 13032 8978
rect 13096 8566 13124 12582
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12912 8350 13032 8378
rect 12912 7857 12940 8350
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 7993 13032 8230
rect 12990 7984 13046 7993
rect 13188 7954 13216 12582
rect 13372 10266 13400 13194
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13266 9208 13322 9217
rect 13372 9178 13400 10202
rect 13464 9761 13492 14282
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13450 9752 13506 9761
rect 13450 9687 13506 9696
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9178 13492 9318
rect 13266 9143 13322 9152
rect 13360 9172 13412 9178
rect 12990 7919 13046 7928
rect 13176 7948 13228 7954
rect 12898 7848 12954 7857
rect 12898 7783 12954 7792
rect 12912 6866 12940 7783
rect 13004 7410 13032 7919
rect 13176 7890 13228 7896
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7546 13124 7686
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12820 6458 12848 6802
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12912 6322 12940 6666
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12820 5545 12848 5646
rect 12900 5568 12952 5574
rect 12806 5536 12862 5545
rect 12900 5510 12952 5516
rect 12806 5471 12862 5480
rect 12544 5222 12664 5250
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12544 5098 12572 5222
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12360 4984 12480 5012
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 12452 4826 12480 4984
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 12544 4282 12572 5034
rect 12636 4826 12664 5102
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12820 4690 12848 5471
rect 12912 4690 12940 5510
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 11980 4072 12032 4078
rect 12808 4072 12860 4078
rect 11980 4014 12032 4020
rect 12806 4040 12808 4049
rect 12860 4040 12862 4049
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11992 800 12020 4014
rect 12806 3975 12862 3984
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 12820 3670 12848 3975
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 13096 3534 13124 6598
rect 13188 4826 13216 6666
rect 13280 6322 13308 9143
rect 13360 9114 13412 9120
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13358 9072 13414 9081
rect 13358 9007 13414 9016
rect 13372 8974 13400 9007
rect 13360 8968 13412 8974
rect 13464 8945 13492 9114
rect 13360 8910 13412 8916
rect 13450 8936 13506 8945
rect 13372 8838 13400 8910
rect 13450 8871 13506 8880
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13450 8392 13506 8401
rect 13450 8327 13506 8336
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13280 5846 13308 6258
rect 13372 6254 13400 7278
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13280 5001 13308 5306
rect 13372 5098 13400 5510
rect 13464 5166 13492 8327
rect 13556 8022 13584 13466
rect 13832 11762 13860 14418
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13924 13297 13952 14214
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 14844 14074 14872 14350
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 13910 13288 13966 13297
rect 13910 13223 13966 13232
rect 14108 12434 14136 14010
rect 14936 13326 14964 14350
rect 15028 13977 15056 14991
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15304 14006 15332 14486
rect 15292 14000 15344 14006
rect 15014 13968 15070 13977
rect 15292 13942 15344 13948
rect 15948 13938 15976 14554
rect 15014 13903 15070 13912
rect 15936 13932 15988 13938
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 14936 12918 14964 13262
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14830 12744 14886 12753
rect 14830 12679 14886 12688
rect 14016 12406 14136 12434
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 11286 13860 11698
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13556 7478 13584 7958
rect 13648 7886 13676 10746
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13648 7342 13676 7822
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13556 6798 13584 7142
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13648 6662 13676 7142
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13740 5778 13768 10134
rect 13832 7478 13860 10202
rect 13924 9654 13952 10542
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13924 9042 13952 9590
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 14016 8974 14044 12406
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 9586 14136 11494
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14200 9466 14228 10406
rect 14568 10198 14596 10610
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14660 9674 14688 12038
rect 14568 9646 14688 9674
rect 14200 9438 14320 9466
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14002 8800 14058 8809
rect 14002 8735 14058 8744
rect 14016 7993 14044 8735
rect 14108 8514 14136 8978
rect 14108 8498 14145 8514
rect 14105 8492 14157 8498
rect 14105 8434 14157 8440
rect 14096 8016 14148 8022
rect 14002 7984 14058 7993
rect 14096 7958 14148 7964
rect 14002 7919 14058 7928
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13818 6624 13874 6633
rect 13818 6559 13874 6568
rect 13832 5914 13860 6559
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13452 5160 13504 5166
rect 13636 5160 13688 5166
rect 13452 5102 13504 5108
rect 13634 5128 13636 5137
rect 13688 5128 13690 5137
rect 13360 5092 13412 5098
rect 13634 5063 13690 5072
rect 13360 5034 13412 5040
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13188 4457 13216 4762
rect 13280 4486 13308 4927
rect 13740 4842 13768 5714
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13556 4826 13860 4842
rect 13556 4820 13872 4826
rect 13556 4814 13820 4820
rect 13268 4480 13320 4486
rect 13174 4448 13230 4457
rect 13268 4422 13320 4428
rect 13174 4383 13230 4392
rect 13556 4078 13584 4814
rect 13820 4762 13872 4768
rect 13726 4720 13782 4729
rect 13726 4655 13782 4664
rect 13740 4282 13768 4655
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13740 4185 13768 4218
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13740 3738 13768 4111
rect 13924 4010 13952 5170
rect 14016 4146 14044 6734
rect 14108 6458 14136 7958
rect 14200 7528 14228 9318
rect 14292 8922 14320 9438
rect 14568 9024 14596 9646
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14752 9364 14780 9522
rect 14844 9489 14872 12679
rect 15028 12434 15056 13903
rect 15936 13874 15988 13880
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15212 13297 15240 13466
rect 15474 13424 15530 13433
rect 15474 13359 15530 13368
rect 15198 13288 15254 13297
rect 15198 13223 15254 13232
rect 15382 12880 15438 12889
rect 15382 12815 15438 12824
rect 14936 12406 15056 12434
rect 14830 9480 14886 9489
rect 14830 9415 14886 9424
rect 14752 9336 14872 9364
rect 14568 8996 14780 9024
rect 14292 8906 14688 8922
rect 14280 8900 14688 8906
rect 14332 8894 14688 8900
rect 14280 8842 14332 8848
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14384 7970 14412 8230
rect 14462 7984 14518 7993
rect 14384 7942 14462 7970
rect 14568 7954 14596 8570
rect 14462 7919 14518 7928
rect 14556 7948 14608 7954
rect 14476 7886 14504 7919
rect 14556 7890 14608 7896
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14200 7500 14320 7528
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14108 5914 14136 6190
rect 14200 6186 14228 7278
rect 14292 6866 14320 7500
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 6866 14504 7142
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14568 6798 14596 7414
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14186 5808 14242 5817
rect 14186 5743 14242 5752
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5273 14136 5510
rect 14200 5284 14228 5743
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14280 5296 14332 5302
rect 14094 5264 14150 5273
rect 14094 5199 14150 5208
rect 14200 5256 14280 5284
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4282 14136 5102
rect 14200 4554 14228 5256
rect 14280 5238 14332 5244
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14476 4690 14504 5102
rect 14568 4758 14596 5170
rect 14660 5166 14688 8894
rect 14752 8566 14780 8996
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14752 7868 14780 8502
rect 14844 7970 14872 9336
rect 14936 8090 14964 12406
rect 15396 12209 15424 12815
rect 15382 12200 15438 12209
rect 15382 12135 15438 12144
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15014 10160 15070 10169
rect 15014 10095 15070 10104
rect 15028 8673 15056 10095
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 15120 8974 15148 9590
rect 15212 9178 15240 11018
rect 15290 10704 15346 10713
rect 15290 10639 15346 10648
rect 15304 9625 15332 10639
rect 15290 9616 15346 9625
rect 15290 9551 15346 9560
rect 15396 9353 15424 12135
rect 15382 9344 15438 9353
rect 15382 9279 15438 9288
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14844 7942 14964 7970
rect 14752 7840 14872 7868
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7546 14780 7686
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14738 7440 14794 7449
rect 14738 7375 14794 7384
rect 14752 7274 14780 7375
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14844 6866 14872 7840
rect 14936 7274 14964 7942
rect 15028 7750 15056 8502
rect 15120 7886 15148 8910
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15212 8265 15240 8434
rect 15396 8401 15424 8774
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 15488 8294 15516 13359
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 9466 15608 12786
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 11830 15700 12310
rect 15764 12170 15792 13126
rect 15856 12646 15884 13670
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15658 10024 15714 10033
rect 15658 9959 15660 9968
rect 15712 9959 15714 9968
rect 15660 9930 15712 9936
rect 15580 9438 15700 9466
rect 15580 9217 15608 9438
rect 15672 9382 15700 9438
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15566 9208 15622 9217
rect 15566 9143 15622 9152
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15476 8288 15528 8294
rect 15198 8256 15254 8265
rect 15476 8230 15528 8236
rect 15198 8191 15254 8200
rect 15580 8106 15608 8298
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15488 8078 15608 8106
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 15028 6934 15056 7686
rect 15212 7342 15240 7686
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14568 4570 14596 4694
rect 14188 4548 14240 4554
rect 14568 4542 14688 4570
rect 14188 4490 14240 4496
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 14016 3534 14044 4082
rect 14200 3738 14228 4490
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14660 4162 14688 4542
rect 14568 4134 14688 4162
rect 14568 3738 14596 4134
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 12820 800 12848 3402
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 14660 3126 14688 3878
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14752 3058 14780 6054
rect 14844 3058 14872 6598
rect 15212 6458 15240 6598
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14936 5778 14964 6122
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14924 5568 14976 5574
rect 14922 5536 14924 5545
rect 14976 5536 14978 5545
rect 14922 5471 14978 5480
rect 14936 4457 14964 5471
rect 15028 4554 15056 6394
rect 15304 6254 15332 7890
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5370 15148 6054
rect 15396 5914 15424 6598
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15200 5568 15252 5574
rect 15488 5545 15516 8078
rect 15566 7576 15622 7585
rect 15566 7511 15622 7520
rect 15200 5510 15252 5516
rect 15474 5536 15530 5545
rect 15212 5409 15240 5510
rect 15474 5471 15530 5480
rect 15198 5400 15254 5409
rect 15108 5364 15160 5370
rect 15198 5335 15254 5344
rect 15292 5364 15344 5370
rect 15108 5306 15160 5312
rect 15292 5306 15344 5312
rect 15304 5273 15332 5306
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 15292 5160 15344 5166
rect 15198 5128 15254 5137
rect 15292 5102 15344 5108
rect 15198 5063 15200 5072
rect 15252 5063 15254 5072
rect 15200 5034 15252 5040
rect 15108 5024 15160 5030
rect 15160 4972 15240 4978
rect 15108 4966 15240 4972
rect 15120 4950 15240 4966
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14922 4448 14978 4457
rect 14922 4383 14978 4392
rect 14936 4282 14964 4383
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14936 3126 14964 4218
rect 15028 4078 15056 4490
rect 15120 4282 15148 4694
rect 15212 4486 15240 4950
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15028 3738 15056 4014
rect 15212 3738 15240 4422
rect 15304 3913 15332 5102
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15488 4826 15516 5034
rect 15580 5001 15608 7511
rect 15672 6118 15700 8230
rect 15764 6866 15792 12106
rect 15856 11665 15884 12378
rect 15948 11898 15976 13874
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15842 11656 15898 11665
rect 15842 11591 15898 11600
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11150 15884 11494
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15948 11257 15976 11290
rect 15934 11248 15990 11257
rect 15934 11183 15990 11192
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10742 15884 11086
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15856 10062 15884 10678
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15934 9888 15990 9897
rect 15934 9823 15990 9832
rect 15844 7200 15896 7206
rect 15948 7188 15976 9823
rect 16040 8634 16068 13194
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16592 12753 16620 12786
rect 16578 12744 16634 12753
rect 16578 12679 16634 12688
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11830 16160 12038
rect 16120 11824 16172 11830
rect 16172 11784 16344 11812
rect 16120 11766 16172 11772
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16132 7818 16160 10950
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15896 7160 15976 7188
rect 15844 7142 15896 7148
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15764 6118 15792 6802
rect 15856 6633 15884 7142
rect 16040 7002 16068 7754
rect 16118 7712 16174 7721
rect 16118 7647 16174 7656
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15842 6624 15898 6633
rect 15842 6559 15898 6568
rect 15856 6390 15884 6559
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15658 5808 15714 5817
rect 15764 5778 15792 6054
rect 15658 5743 15714 5752
rect 15752 5772 15804 5778
rect 15672 5574 15700 5743
rect 15752 5714 15804 5720
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15752 5160 15804 5166
rect 15856 5148 15884 6326
rect 15948 6322 15976 6734
rect 16132 6338 16160 7647
rect 16224 6798 16252 8366
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16040 6310 16160 6338
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15804 5120 15884 5148
rect 15752 5102 15804 5108
rect 15566 4992 15622 5001
rect 15566 4927 15622 4936
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15384 4072 15436 4078
rect 15382 4040 15384 4049
rect 15436 4040 15438 4049
rect 15382 3975 15438 3984
rect 15476 3936 15528 3942
rect 15290 3904 15346 3913
rect 15580 3924 15608 4927
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15528 3896 15608 3924
rect 15476 3878 15528 3884
rect 15290 3839 15346 3848
rect 15304 3738 15332 3839
rect 15672 3738 15700 4082
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15028 3534 15056 3674
rect 15304 3618 15332 3674
rect 15476 3664 15528 3670
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15212 3590 15332 3618
rect 15474 3632 15476 3641
rect 15528 3632 15530 3641
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 13648 800 13676 2926
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14660 1578 14688 2926
rect 15120 2530 15148 3538
rect 15212 3233 15240 3590
rect 15474 3567 15530 3576
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15580 3398 15608 3538
rect 15764 3398 15792 5102
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15198 3224 15254 3233
rect 15198 3159 15254 3168
rect 15212 2650 15240 3159
rect 15382 3088 15438 3097
rect 15382 3023 15384 3032
rect 15436 3023 15438 3032
rect 15384 2994 15436 3000
rect 15580 2922 15608 3334
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15198 2544 15254 2553
rect 15016 2508 15068 2514
rect 15120 2502 15198 2530
rect 15198 2479 15254 2488
rect 15016 2450 15068 2456
rect 15028 2417 15056 2450
rect 15014 2408 15070 2417
rect 15014 2343 15070 2352
rect 14476 1550 14688 1578
rect 14476 800 14504 1550
rect 15304 800 15332 2790
rect 15672 2650 15700 3062
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 15856 762 15884 4558
rect 15948 4282 15976 5782
rect 16040 5658 16068 6310
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16132 5914 16160 6190
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16040 5630 16160 5658
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16040 4162 16068 5510
rect 16132 5302 16160 5630
rect 16224 5370 16252 6734
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4622 16160 4966
rect 16316 4690 16344 11784
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16868 11082 16896 13194
rect 16960 12714 16988 14826
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10810 16620 10950
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16408 7970 16436 8570
rect 16868 8430 16896 11018
rect 16960 9178 16988 12106
rect 17052 12102 17080 14214
rect 17604 14006 17632 16510
rect 17866 16400 17922 16510
rect 18878 14920 18934 14929
rect 18878 14855 18934 14864
rect 17958 14512 18014 14521
rect 17958 14447 18014 14456
rect 17972 14113 18000 14447
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17958 14104 18014 14113
rect 17958 14039 18014 14048
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 18064 13870 18092 14350
rect 18420 14340 18472 14346
rect 18420 14282 18472 14288
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13326 18092 13806
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17788 12617 17816 12922
rect 18064 12850 18092 13262
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17774 12608 17830 12617
rect 17774 12543 17830 12552
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16960 8786 16988 9114
rect 17052 8888 17080 12038
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 9994 17172 11630
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11150 17356 11494
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17314 10976 17370 10985
rect 17314 10911 17370 10920
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17144 9625 17172 9930
rect 17130 9616 17186 9625
rect 17130 9551 17186 9560
rect 17052 8860 17264 8888
rect 16960 8758 17080 8786
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 8537 16988 8570
rect 16946 8528 17002 8537
rect 16946 8463 17002 8472
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16408 7954 16620 7970
rect 16408 7948 16632 7954
rect 16408 7942 16580 7948
rect 16580 7890 16632 7896
rect 16578 7848 16634 7857
rect 16578 7783 16634 7792
rect 16856 7812 16908 7818
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16486 7712 16542 7721
rect 16408 5778 16436 7686
rect 16486 7647 16542 7656
rect 16500 7274 16528 7647
rect 16592 7410 16620 7783
rect 16856 7754 16908 7760
rect 16868 7585 16896 7754
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16854 7576 16910 7585
rect 16854 7511 16910 7520
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16684 7274 16712 7414
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16776 7188 16804 7278
rect 16960 7274 16988 7686
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16776 7160 16896 7188
rect 16868 7154 16896 7160
rect 16868 7126 16988 7154
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16960 7002 16988 7126
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17052 6882 17080 8758
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7886 17172 8230
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17052 6866 17172 6882
rect 17052 6860 17184 6866
rect 17052 6854 17132 6860
rect 17132 6802 17184 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16762 6760 16818 6769
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6497 16528 6598
rect 16486 6488 16542 6497
rect 16486 6423 16542 6432
rect 16684 6254 16712 6734
rect 16762 6695 16818 6704
rect 16776 6390 16804 6695
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16764 6384 16816 6390
rect 16762 6352 16764 6361
rect 16816 6352 16818 6361
rect 16762 6287 16818 6296
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16120 4616 16172 4622
rect 16316 4570 16344 4626
rect 16120 4558 16172 4564
rect 15948 4134 16068 4162
rect 16224 4542 16344 4570
rect 15948 3942 15976 4134
rect 16224 4078 16252 4542
rect 16408 4146 16436 4966
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16304 4072 16356 4078
rect 16592 4026 16620 4558
rect 16764 4480 16816 4486
rect 16762 4448 16764 4457
rect 16816 4448 16818 4457
rect 16762 4383 16818 4392
rect 16868 4298 16896 5238
rect 16960 5166 16988 6598
rect 17144 6186 17172 6802
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17236 5846 17264 8860
rect 17328 6730 17356 10911
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 9648 17460 9654
rect 17406 9616 17408 9625
rect 17460 9616 17462 9625
rect 17406 9551 17462 9560
rect 17420 7818 17448 9551
rect 17512 9353 17540 10406
rect 17788 10130 17816 12543
rect 18156 12442 18184 13126
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11082 17908 12038
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17880 10062 17908 11018
rect 17868 10056 17920 10062
rect 17774 10024 17830 10033
rect 17868 9998 17920 10004
rect 17774 9959 17830 9968
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17498 9344 17554 9353
rect 17498 9279 17554 9288
rect 17512 8634 17540 9279
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17512 7993 17540 8570
rect 17604 8090 17632 9522
rect 17696 9382 17724 9522
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 8430 17724 9318
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17498 7984 17554 7993
rect 17498 7919 17554 7928
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17316 6724 17368 6730
rect 17316 6666 17368 6672
rect 17420 6186 17448 7346
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17314 5944 17370 5953
rect 17314 5879 17370 5888
rect 17408 5908 17460 5914
rect 17328 5846 17356 5879
rect 17408 5850 17460 5856
rect 17224 5840 17276 5846
rect 17038 5808 17094 5817
rect 17224 5782 17276 5788
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17038 5743 17094 5752
rect 17052 5710 17080 5743
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17236 5370 17264 5510
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4570 16988 5102
rect 16960 4542 17080 4570
rect 16946 4448 17002 4457
rect 16946 4383 17002 4392
rect 16304 4014 16356 4020
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 2417 15976 3878
rect 16040 3602 16068 3946
rect 16118 3632 16174 3641
rect 16028 3596 16080 3602
rect 16118 3567 16120 3576
rect 16028 3538 16080 3544
rect 16172 3567 16174 3576
rect 16120 3538 16172 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 3194 16252 3470
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16316 3097 16344 4014
rect 16408 3998 16620 4026
rect 16776 4270 16896 4298
rect 16776 4010 16804 4270
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16764 4004 16816 4010
rect 16408 3738 16436 3998
rect 16764 3946 16816 3952
rect 16868 3942 16896 4150
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16578 3632 16634 3641
rect 16396 3596 16448 3602
rect 16578 3567 16634 3576
rect 16396 3538 16448 3544
rect 16302 3088 16358 3097
rect 16302 3023 16358 3032
rect 16210 2680 16266 2689
rect 16408 2650 16436 3538
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16500 2854 16528 3334
rect 16592 3126 16620 3567
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 16210 2615 16212 2624
rect 16264 2615 16266 2624
rect 16396 2644 16448 2650
rect 16212 2586 16264 2592
rect 16396 2586 16448 2592
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16684 2446 16712 2518
rect 16580 2440 16632 2446
rect 15934 2408 15990 2417
rect 16580 2382 16632 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 15934 2343 15990 2352
rect 16592 2310 16620 2382
rect 16868 2310 16896 3878
rect 16960 3738 16988 4383
rect 17052 4214 17080 4542
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17052 3194 17080 3946
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16946 2952 17002 2961
rect 16946 2887 17002 2896
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16040 1834 16068 2246
rect 16028 1828 16080 1834
rect 16028 1770 16080 1776
rect 16040 870 16160 898
rect 16040 762 16068 870
rect 16132 800 16160 870
rect 16960 800 16988 2887
rect 17144 2774 17172 5238
rect 17328 5166 17356 5510
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17222 4856 17278 4865
rect 17222 4791 17278 4800
rect 17236 4554 17264 4791
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17420 4282 17448 5850
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17314 4176 17370 4185
rect 17224 4140 17276 4146
rect 17314 4111 17370 4120
rect 17224 4082 17276 4088
rect 17236 3670 17264 4082
rect 17328 3738 17356 4111
rect 17406 3904 17462 3913
rect 17406 3839 17462 3848
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17420 3194 17448 3839
rect 17512 3670 17540 7822
rect 17604 7410 17632 8026
rect 17696 7750 17724 8366
rect 17788 7834 17816 9959
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9722 17908 9862
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17880 8498 17908 9658
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17960 8832 18012 8838
rect 18064 8809 18092 9318
rect 17960 8774 18012 8780
rect 18050 8800 18106 8809
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 8090 17908 8230
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17788 7806 17908 7834
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17696 7449 17724 7686
rect 17682 7440 17738 7449
rect 17592 7404 17644 7410
rect 17682 7375 17738 7384
rect 17592 7346 17644 7352
rect 17788 7313 17816 7686
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17880 6984 17908 7806
rect 17696 6956 17908 6984
rect 17592 6452 17644 6458
rect 17696 6440 17724 6956
rect 17866 6896 17922 6905
rect 17866 6831 17922 6840
rect 17880 6730 17908 6831
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17776 6656 17828 6662
rect 17774 6624 17776 6633
rect 17828 6624 17830 6633
rect 17774 6559 17830 6568
rect 17696 6412 17816 6440
rect 17592 6394 17644 6400
rect 17604 4622 17632 6394
rect 17682 6352 17738 6361
rect 17788 6322 17816 6412
rect 17682 6287 17738 6296
rect 17776 6316 17828 6322
rect 17696 4826 17724 6287
rect 17776 6258 17828 6264
rect 17880 5914 17908 6666
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17774 5400 17830 5409
rect 17774 5335 17830 5344
rect 17788 5234 17816 5335
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17774 4720 17830 4729
rect 17880 4706 17908 5646
rect 17830 4678 17908 4706
rect 17972 4690 18000 8774
rect 18050 8735 18106 8744
rect 18156 8480 18184 12378
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18064 8452 18184 8480
rect 18064 7954 18092 8452
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 8265 18184 8298
rect 18142 8256 18198 8265
rect 18142 8191 18198 8200
rect 18248 8106 18276 10406
rect 18326 9072 18382 9081
rect 18326 9007 18382 9016
rect 18156 8078 18276 8106
rect 18340 8090 18368 9007
rect 18432 8838 18460 14282
rect 18694 14240 18750 14249
rect 18694 14175 18750 14184
rect 18510 12064 18566 12073
rect 18510 11999 18566 12008
rect 18524 10470 18552 11999
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18328 8084 18380 8090
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18156 7886 18184 8078
rect 18328 8026 18380 8032
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18418 7984 18474 7993
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18064 5914 18092 7375
rect 18156 6934 18184 7822
rect 18248 7546 18276 7958
rect 18328 7948 18380 7954
rect 18418 7919 18474 7928
rect 18328 7890 18380 7896
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 7410 18368 7890
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18340 6934 18368 7346
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18144 6792 18196 6798
rect 18328 6792 18380 6798
rect 18144 6734 18196 6740
rect 18326 6760 18328 6769
rect 18380 6760 18382 6769
rect 18156 6202 18184 6734
rect 18326 6695 18382 6704
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6322 18368 6598
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18156 6174 18368 6202
rect 18340 6118 18368 6174
rect 18328 6112 18380 6118
rect 18142 6080 18198 6089
rect 18328 6054 18380 6060
rect 18142 6015 18198 6024
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17960 4684 18012 4690
rect 17774 4655 17830 4664
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17500 3664 17552 3670
rect 17696 3618 17724 4082
rect 17500 3606 17552 3612
rect 17604 3590 17724 3618
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17512 3058 17540 3470
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17144 2746 17264 2774
rect 17038 2680 17094 2689
rect 17038 2615 17094 2624
rect 17052 2582 17080 2615
rect 17236 2582 17264 2746
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 17224 2576 17276 2582
rect 17512 2530 17540 2994
rect 17224 2518 17276 2524
rect 17328 2502 17540 2530
rect 17328 2446 17356 2502
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17604 2378 17632 3590
rect 17788 3482 17816 4655
rect 17960 4626 18012 4632
rect 17868 4616 17920 4622
rect 17866 4584 17868 4593
rect 17920 4584 17922 4593
rect 17866 4519 17922 4528
rect 17960 4548 18012 4554
rect 17880 4162 17908 4519
rect 17960 4490 18012 4496
rect 17972 4321 18000 4490
rect 17958 4312 18014 4321
rect 17958 4247 18014 4256
rect 17880 4134 18000 4162
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17696 3454 17816 3482
rect 17696 3126 17724 3454
rect 17776 3392 17828 3398
rect 17880 3369 17908 4014
rect 17776 3334 17828 3340
rect 17866 3360 17922 3369
rect 17684 3120 17736 3126
rect 17788 3097 17816 3334
rect 17866 3295 17922 3304
rect 17972 3210 18000 4134
rect 18064 3641 18092 5102
rect 18156 4010 18184 6015
rect 18234 5808 18290 5817
rect 18234 5743 18290 5752
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18248 3738 18276 5743
rect 18340 5658 18368 6054
rect 18432 5914 18460 7919
rect 18524 7750 18552 10406
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18510 7168 18566 7177
rect 18510 7103 18566 7112
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18340 5630 18460 5658
rect 18326 5536 18382 5545
rect 18326 5471 18382 5480
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18050 3632 18106 3641
rect 18050 3567 18106 3576
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 17880 3182 18000 3210
rect 17684 3062 17736 3068
rect 17774 3088 17830 3097
rect 17774 3023 17830 3032
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17696 1578 17724 2926
rect 17880 2650 17908 3182
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17972 2582 18000 3062
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 18064 2514 18092 3470
rect 18142 3224 18198 3233
rect 18340 3194 18368 5471
rect 18142 3159 18198 3168
rect 18328 3188 18380 3194
rect 18156 3058 18184 3159
rect 18328 3130 18380 3136
rect 18432 3058 18460 5630
rect 18524 4826 18552 7103
rect 18616 6633 18644 9318
rect 18708 7041 18736 14175
rect 18786 11792 18842 11801
rect 18786 11727 18842 11736
rect 18800 11082 18828 11727
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18694 7032 18750 7041
rect 18694 6967 18750 6976
rect 18694 6896 18750 6905
rect 18694 6831 18750 6840
rect 18602 6624 18658 6633
rect 18602 6559 18658 6568
rect 18604 5704 18656 5710
rect 18602 5672 18604 5681
rect 18656 5672 18658 5681
rect 18602 5607 18658 5616
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18510 4720 18566 4729
rect 18510 4655 18566 4664
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18156 2582 18184 2858
rect 18524 2650 18552 4655
rect 18616 4604 18644 5607
rect 18708 4758 18736 6831
rect 18800 6730 18828 9386
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18786 6488 18842 6497
rect 18786 6423 18842 6432
rect 18800 5370 18828 6423
rect 18892 5409 18920 14855
rect 18970 14376 19026 14385
rect 18970 14311 19026 14320
rect 18878 5400 18934 5409
rect 18788 5364 18840 5370
rect 18878 5335 18934 5344
rect 18788 5306 18840 5312
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18616 4576 18736 4604
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17868 2440 17920 2446
rect 17866 2408 17868 2417
rect 17920 2408 17922 2417
rect 17866 2343 17922 2352
rect 17696 1550 17816 1578
rect 17788 800 17816 1550
rect 18616 800 18644 2926
rect 18708 2378 18736 4576
rect 18984 3602 19012 14311
rect 19062 14104 19118 14113
rect 19062 14039 19118 14048
rect 19076 4078 19104 14039
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19168 5370 19196 11018
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19260 3738 19288 6734
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 19352 2582 19380 6394
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 15856 734 16068 762
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< via2 >>
rect 2134 14320 2190 14376
rect 1582 14048 1638 14104
rect 1858 13504 1914 13560
rect 1858 13252 1914 13288
rect 1858 13232 1860 13252
rect 1860 13232 1912 13252
rect 1912 13232 1914 13252
rect 2410 13812 2412 13832
rect 2412 13812 2464 13832
rect 2464 13812 2466 13832
rect 2410 13776 2466 13812
rect 2410 12960 2466 13016
rect 2502 12688 2558 12744
rect 2870 15408 2926 15464
rect 2778 15136 2834 15192
rect 3054 14864 3110 14920
rect 2962 14592 3018 14648
rect 2962 14320 3018 14376
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 3606 13640 3662 13696
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 5998 13368 6054 13424
rect 2686 13268 2688 13288
rect 2688 13268 2740 13288
rect 2740 13268 2742 13288
rect 2686 13232 2742 13268
rect 1766 11328 1822 11384
rect 1582 9696 1638 9752
rect 1306 7248 1362 7304
rect 1306 6976 1362 7032
rect 1306 6568 1362 6624
rect 1582 6840 1638 6896
rect 1950 8880 2006 8936
rect 2318 10376 2374 10432
rect 2778 12416 2834 12472
rect 2594 10512 2650 10568
rect 1674 6704 1730 6760
rect 1582 6160 1638 6216
rect 1398 4800 1454 4856
rect 1950 6316 2006 6352
rect 1950 6296 1952 6316
rect 1952 6296 2004 6316
rect 2004 6296 2006 6316
rect 2410 7520 2466 7576
rect 2594 9832 2650 9888
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 3514 12280 3570 12336
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 2962 10648 3018 10704
rect 2962 10376 3018 10432
rect 2962 9696 3018 9752
rect 2962 9152 3018 9208
rect 2686 8744 2742 8800
rect 2042 6160 2098 6216
rect 1858 5616 1914 5672
rect 1858 4528 1914 4584
rect 1214 3032 1270 3088
rect 2042 4936 2098 4992
rect 2226 4256 2282 4312
rect 2042 3848 2098 3904
rect 1490 2624 1546 2680
rect 1858 2080 1914 2136
rect 1674 1536 1730 1592
rect 2134 3576 2190 3632
rect 2962 8336 3018 8392
rect 2870 8064 2926 8120
rect 2686 7948 2742 7984
rect 2686 7928 2688 7948
rect 2688 7928 2740 7948
rect 2740 7928 2742 7948
rect 2410 3732 2466 3768
rect 2410 3712 2412 3732
rect 2412 3712 2464 3732
rect 2464 3712 2466 3732
rect 2870 7384 2926 7440
rect 2778 5888 2834 5944
rect 3514 10648 3570 10704
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3514 9696 3570 9752
rect 3790 11600 3846 11656
rect 4066 12180 4068 12200
rect 4068 12180 4120 12200
rect 4120 12180 4122 12200
rect 4066 12144 4122 12180
rect 4710 12144 4766 12200
rect 4158 11736 4214 11792
rect 4066 11464 4122 11520
rect 4066 10784 4122 10840
rect 3974 10648 4030 10704
rect 3698 9560 3754 9616
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3054 7384 3110 7440
rect 3422 7928 3478 7984
rect 4066 9988 4122 10024
rect 4066 9968 4068 9988
rect 4068 9968 4120 9988
rect 4120 9968 4122 9988
rect 3882 9016 3938 9072
rect 3698 8336 3754 8392
rect 4066 9152 4122 9208
rect 3514 7792 3570 7848
rect 3238 7248 3294 7304
rect 2962 6296 3018 6352
rect 2778 5228 2834 5264
rect 2778 5208 2780 5228
rect 2780 5208 2832 5228
rect 2832 5208 2834 5228
rect 2778 5092 2834 5128
rect 2778 5072 2780 5092
rect 2780 5072 2832 5092
rect 2832 5072 2834 5092
rect 2778 4004 2834 4040
rect 2778 3984 2780 4004
rect 2780 3984 2832 4004
rect 2832 3984 2834 4004
rect 2594 2352 2650 2408
rect 2870 2896 2926 2952
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3146 6860 3202 6896
rect 3146 6840 3148 6860
rect 3148 6840 3200 6860
rect 3200 6840 3202 6860
rect 3606 7520 3662 7576
rect 3606 7112 3662 7168
rect 3882 7812 3938 7848
rect 3882 7792 3884 7812
rect 3884 7792 3936 7812
rect 3936 7792 3938 7812
rect 3882 7284 3884 7304
rect 3884 7284 3936 7304
rect 3936 7284 3938 7304
rect 3882 7248 3938 7284
rect 3790 6976 3846 7032
rect 3882 6840 3938 6896
rect 4066 8608 4122 8664
rect 4158 8472 4214 8528
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 3330 5244 3332 5264
rect 3332 5244 3384 5264
rect 3384 5244 3386 5264
rect 3330 5208 3386 5244
rect 3422 5108 3424 5128
rect 3424 5108 3476 5128
rect 3476 5108 3478 5128
rect 3422 5072 3478 5108
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 3146 4528 3202 4584
rect 3514 4120 3570 4176
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3054 3440 3110 3496
rect 4158 7248 4214 7304
rect 4066 5364 4122 5400
rect 4066 5344 4068 5364
rect 4068 5344 4120 5364
rect 4120 5344 4122 5364
rect 3974 4528 4030 4584
rect 3882 3168 3938 3224
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 2778 1808 2834 1864
rect 4710 11736 4766 11792
rect 4434 8880 4490 8936
rect 4342 8336 4398 8392
rect 4618 9424 4674 9480
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 4894 11636 4896 11656
rect 4896 11636 4948 11656
rect 4948 11636 4950 11656
rect 4894 11600 4950 11636
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5078 8744 5134 8800
rect 4986 8336 5042 8392
rect 5906 9036 5962 9072
rect 5906 9016 5908 9036
rect 5908 9016 5960 9036
rect 5960 9016 5962 9036
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5078 7520 5134 7576
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5262 6568 5318 6624
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5814 6432 5870 6488
rect 4986 5616 5042 5672
rect 5538 5652 5540 5672
rect 5540 5652 5592 5672
rect 5592 5652 5594 5672
rect 5538 5616 5594 5652
rect 6734 11192 6790 11248
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 6182 10104 6238 10160
rect 6182 9424 6238 9480
rect 6182 8472 6238 8528
rect 6182 7112 6238 7168
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 6550 8880 6606 8936
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 6918 13912 6974 13968
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 6734 9968 6790 10024
rect 6826 8744 6882 8800
rect 6734 8472 6790 8528
rect 6550 7248 6606 7304
rect 6458 6296 6514 6352
rect 6734 5636 6790 5672
rect 6734 5616 6736 5636
rect 6736 5616 6788 5636
rect 6788 5616 6790 5636
rect 6826 5480 6882 5536
rect 7010 7248 7066 7304
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 8022 11056 8078 11112
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7194 6976 7250 7032
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 8390 10512 8446 10568
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7838 7948 7894 7984
rect 7838 7928 7840 7948
rect 7840 7928 7892 7948
rect 7892 7928 7894 7948
rect 7562 7520 7618 7576
rect 8114 8064 8170 8120
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7286 5344 7342 5400
rect 7010 4664 7066 4720
rect 7746 6568 7802 6624
rect 8022 6452 8078 6488
rect 8022 6432 8024 6452
rect 8024 6432 8076 6452
rect 8076 6432 8078 6452
rect 7746 6196 7748 6216
rect 7748 6196 7800 6216
rect 7800 6196 7802 6216
rect 7746 6160 7802 6196
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7562 5344 7618 5400
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 8390 6296 8446 6352
rect 8206 4664 8262 4720
rect 8850 13776 8906 13832
rect 9218 13232 9274 13288
rect 8850 10376 8906 10432
rect 8758 9968 8814 10024
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9218 10648 9274 10704
rect 9034 8744 9090 8800
rect 8850 7248 8906 7304
rect 8942 6840 8998 6896
rect 8942 6704 8998 6760
rect 8758 6332 8760 6352
rect 8760 6332 8812 6352
rect 8812 6332 8814 6352
rect 8758 6296 8814 6332
rect 8850 5208 8906 5264
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10046 10104 10102 10160
rect 11426 13368 11482 13424
rect 10782 13232 10838 13288
rect 10230 9868 10232 9888
rect 10232 9868 10284 9888
rect 10284 9868 10286 9888
rect 10230 9832 10286 9868
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10138 9632 10194 9688
rect 9402 6432 9458 6488
rect 10046 9152 10102 9208
rect 10322 9424 10378 9480
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10322 7928 10378 7984
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10138 6704 10194 6760
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9678 5616 9734 5672
rect 9310 5480 9366 5536
rect 10690 9832 10746 9888
rect 10690 7928 10746 7984
rect 10690 7384 10746 7440
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9770 5208 9826 5264
rect 10414 5516 10416 5536
rect 10416 5516 10468 5536
rect 10468 5516 10470 5536
rect 10414 5480 10470 5516
rect 9034 3848 9090 3904
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10322 4684 10378 4720
rect 10322 4664 10324 4684
rect 10324 4664 10376 4684
rect 10376 4664 10378 4684
rect 11150 11736 11206 11792
rect 11058 11500 11060 11520
rect 11060 11500 11112 11520
rect 11112 11500 11114 11520
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 15014 15000 15070 15056
rect 11702 13776 11758 13832
rect 10874 9288 10930 9344
rect 10874 8472 10930 8528
rect 11058 11464 11114 11500
rect 10966 5616 11022 5672
rect 10782 5072 10838 5128
rect 11150 6296 11206 6352
rect 11242 5616 11298 5672
rect 11426 10548 11428 10568
rect 11428 10548 11480 10568
rect 11480 10548 11482 10568
rect 11426 10512 11482 10548
rect 11426 10104 11482 10160
rect 11794 11464 11850 11520
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 10690 4528 10746 4584
rect 10782 3984 10838 4040
rect 10506 3712 10562 3768
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 11702 7656 11758 7712
rect 11702 7112 11758 7168
rect 12898 11192 12954 11248
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 11886 6604 11888 6624
rect 11888 6604 11940 6624
rect 11940 6604 11942 6624
rect 11886 6568 11942 6604
rect 11886 5752 11942 5808
rect 12622 6432 12678 6488
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12530 5616 12586 5672
rect 12990 9560 13046 9616
rect 12990 7928 13046 7984
rect 13266 9152 13322 9208
rect 13450 9696 13506 9752
rect 12898 7792 12954 7848
rect 12806 5480 12862 5536
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 12806 4020 12808 4040
rect 12808 4020 12860 4040
rect 12860 4020 12862 4040
rect 12806 3984 12862 4020
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 13358 9016 13414 9072
rect 13450 8880 13506 8936
rect 13450 8336 13506 8392
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 13910 13232 13966 13288
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 15014 13912 15070 13968
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14830 12688 14886 12744
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 14002 8744 14058 8800
rect 14002 7928 14058 7984
rect 13818 6568 13874 6624
rect 13634 5108 13636 5128
rect 13636 5108 13688 5128
rect 13688 5108 13690 5128
rect 13634 5072 13690 5108
rect 13266 4936 13322 4992
rect 13174 4392 13230 4448
rect 13726 4664 13782 4720
rect 13726 4120 13782 4176
rect 15474 13368 15530 13424
rect 15198 13232 15254 13288
rect 15382 12824 15438 12880
rect 14830 9424 14886 9480
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14462 7928 14518 7984
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14186 5752 14242 5808
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14094 5208 14150 5264
rect 15382 12144 15438 12200
rect 15014 10104 15070 10160
rect 15290 10648 15346 10704
rect 15290 9560 15346 9616
rect 15382 9288 15438 9344
rect 15014 8608 15070 8664
rect 14738 7384 14794 7440
rect 15382 8336 15438 8392
rect 15658 9988 15714 10024
rect 15658 9968 15660 9988
rect 15660 9968 15712 9988
rect 15712 9968 15714 9988
rect 15566 9152 15622 9208
rect 15198 8200 15254 8256
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14922 5516 14924 5536
rect 14924 5516 14976 5536
rect 14976 5516 14978 5536
rect 14922 5480 14978 5516
rect 15566 7520 15622 7576
rect 15474 5480 15530 5536
rect 15198 5344 15254 5400
rect 15290 5208 15346 5264
rect 15198 5092 15254 5128
rect 15198 5072 15200 5092
rect 15200 5072 15252 5092
rect 15252 5072 15254 5092
rect 14922 4392 14978 4448
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 15842 11600 15898 11656
rect 15934 11192 15990 11248
rect 15934 9832 15990 9888
rect 16578 12688 16634 12744
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16118 7656 16174 7712
rect 15842 6568 15898 6624
rect 15658 5752 15714 5808
rect 15566 4936 15622 4992
rect 15382 4020 15384 4040
rect 15384 4020 15436 4040
rect 15436 4020 15438 4040
rect 15382 3984 15438 4020
rect 15290 3848 15346 3904
rect 15474 3612 15476 3632
rect 15476 3612 15528 3632
rect 15528 3612 15530 3632
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 15474 3576 15530 3612
rect 15198 3168 15254 3224
rect 15382 3052 15438 3088
rect 15382 3032 15384 3052
rect 15384 3032 15436 3052
rect 15436 3032 15438 3052
rect 15198 2488 15254 2544
rect 15014 2352 15070 2408
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 18878 14864 18934 14920
rect 17958 14456 18014 14512
rect 17958 14048 18014 14104
rect 17774 12552 17830 12608
rect 17314 10920 17370 10976
rect 17130 9560 17186 9616
rect 16946 8472 17002 8528
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16578 7792 16634 7848
rect 16486 7656 16542 7712
rect 16854 7520 16910 7576
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16486 6432 16542 6488
rect 16762 6704 16818 6760
rect 16762 6332 16764 6352
rect 16764 6332 16816 6352
rect 16816 6332 16818 6352
rect 16762 6296 16818 6332
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16762 4428 16764 4448
rect 16764 4428 16816 4448
rect 16816 4428 16818 4448
rect 16762 4392 16818 4428
rect 17406 9596 17408 9616
rect 17408 9596 17460 9616
rect 17460 9596 17462 9616
rect 17406 9560 17462 9596
rect 17774 9968 17830 10024
rect 17498 9288 17554 9344
rect 17498 7928 17554 7984
rect 17314 5888 17370 5944
rect 17038 5752 17094 5808
rect 16946 4392 17002 4448
rect 16118 3596 16174 3632
rect 16118 3576 16120 3596
rect 16120 3576 16172 3596
rect 16172 3576 16174 3596
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16578 3576 16634 3632
rect 16302 3032 16358 3088
rect 16210 2644 16266 2680
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 16210 2624 16212 2644
rect 16212 2624 16264 2644
rect 16264 2624 16266 2644
rect 15934 2352 15990 2408
rect 16946 2896 17002 2952
rect 17222 4800 17278 4856
rect 17314 4120 17370 4176
rect 17406 3848 17462 3904
rect 17682 7384 17738 7440
rect 17774 7248 17830 7304
rect 17866 6840 17922 6896
rect 17774 6604 17776 6624
rect 17776 6604 17828 6624
rect 17828 6604 17830 6624
rect 17774 6568 17830 6604
rect 17682 6296 17738 6352
rect 17774 5344 17830 5400
rect 17774 4664 17830 4720
rect 18050 8744 18106 8800
rect 18142 8200 18198 8256
rect 18326 9016 18382 9072
rect 18694 14184 18750 14240
rect 18510 12008 18566 12064
rect 18050 7384 18106 7440
rect 18418 7928 18474 7984
rect 18326 6740 18328 6760
rect 18328 6740 18380 6760
rect 18380 6740 18382 6760
rect 18326 6704 18382 6740
rect 18142 6024 18198 6080
rect 17038 2624 17094 2680
rect 17866 4564 17868 4584
rect 17868 4564 17920 4584
rect 17920 4564 17922 4584
rect 17866 4528 17922 4564
rect 17958 4256 18014 4312
rect 17866 3304 17922 3360
rect 18234 5752 18290 5808
rect 18510 7112 18566 7168
rect 18326 5480 18382 5536
rect 18050 3576 18106 3632
rect 17774 3032 17830 3088
rect 18142 3168 18198 3224
rect 18786 11736 18842 11792
rect 18694 6976 18750 7032
rect 18694 6840 18750 6896
rect 18602 6568 18658 6624
rect 18602 5652 18604 5672
rect 18604 5652 18656 5672
rect 18656 5652 18658 5672
rect 18602 5616 18658 5652
rect 18510 4664 18566 4720
rect 18786 6432 18842 6488
rect 18970 14320 19026 14376
rect 18878 5344 18934 5400
rect 17866 2388 17868 2408
rect 17868 2388 17920 2408
rect 17920 2388 17922 2408
rect 17866 2352 17922 2388
rect 19062 14048 19118 14104
<< metal3 >>
rect 0 15466 800 15496
rect 2865 15466 2931 15469
rect 0 15464 2931 15466
rect 0 15408 2870 15464
rect 2926 15408 2931 15464
rect 0 15406 2931 15408
rect 0 15376 800 15406
rect 2865 15403 2931 15406
rect 0 15194 800 15224
rect 2773 15194 2839 15197
rect 0 15192 12450 15194
rect 0 15136 2778 15192
rect 2834 15136 12450 15192
rect 0 15134 12450 15136
rect 0 15104 800 15134
rect 2773 15131 2839 15134
rect 0 14922 800 14952
rect 3049 14922 3115 14925
rect 9070 14922 9076 14924
rect 0 14862 2698 14922
rect 2922 14920 9076 14922
rect 2922 14864 3054 14920
rect 3110 14864 9076 14920
rect 2922 14862 9076 14864
rect 0 14832 800 14862
rect 2638 14786 2698 14862
rect 3006 14859 3115 14862
rect 9070 14860 9076 14862
rect 9140 14860 9146 14924
rect 12390 14922 12450 15134
rect 15009 15058 15075 15061
rect 15009 15056 19074 15058
rect 15009 15000 15014 15056
rect 15070 15000 19074 15056
rect 15009 14998 19074 15000
rect 15009 14995 15075 14998
rect 18873 14922 18939 14925
rect 12390 14920 18939 14922
rect 12390 14864 18878 14920
rect 18934 14864 18939 14920
rect 12390 14862 18939 14864
rect 18873 14859 18939 14862
rect 3006 14786 3066 14859
rect 2638 14726 3066 14786
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 17953 14514 18019 14517
rect 2730 14512 18019 14514
rect 2730 14456 17958 14512
rect 18014 14456 18019 14512
rect 2730 14454 18019 14456
rect 19014 14514 19074 14998
rect 19200 14514 20000 14544
rect 19014 14454 20000 14514
rect 0 14378 800 14408
rect 2129 14378 2195 14381
rect 2730 14378 2790 14454
rect 17953 14451 18019 14454
rect 19200 14424 20000 14454
rect 0 14376 2790 14378
rect 0 14320 2134 14376
rect 2190 14320 2790 14376
rect 0 14318 2790 14320
rect 2957 14378 3023 14381
rect 18965 14378 19031 14381
rect 2957 14376 19031 14378
rect 2957 14320 2962 14376
rect 3018 14320 18970 14376
rect 19026 14320 19031 14376
rect 2957 14318 19031 14320
rect 0 14288 800 14318
rect 2129 14315 2195 14318
rect 2957 14315 3023 14318
rect 18965 14315 19031 14318
rect 18689 14242 18755 14245
rect 19200 14242 20000 14272
rect 18689 14240 20000 14242
rect 18689 14184 18694 14240
rect 18750 14184 20000 14240
rect 18689 14182 20000 14184
rect 18689 14179 18755 14182
rect 5394 14176 5710 14177
rect 0 14106 800 14136
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 19200 14152 20000 14182
rect 14290 14111 14606 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 800 14046
rect 1577 14043 1643 14046
rect 17953 14106 18019 14109
rect 19057 14106 19123 14109
rect 17953 14104 19123 14106
rect 17953 14048 17958 14104
rect 18014 14048 19062 14104
rect 19118 14048 19123 14104
rect 17953 14046 19123 14048
rect 17953 14043 18019 14046
rect 19057 14043 19123 14046
rect 6913 13970 6979 13973
rect 15009 13970 15075 13973
rect 6913 13968 15075 13970
rect 6913 13912 6918 13968
rect 6974 13912 15014 13968
rect 15070 13912 15075 13968
rect 6913 13910 15075 13912
rect 6913 13907 6979 13910
rect 15009 13907 15075 13910
rect 15694 13908 15700 13972
rect 15764 13970 15770 13972
rect 19200 13970 20000 14000
rect 15764 13910 20000 13970
rect 15764 13908 15770 13910
rect 19200 13880 20000 13910
rect 0 13834 800 13864
rect 2405 13834 2471 13837
rect 0 13832 2471 13834
rect 0 13776 2410 13832
rect 2466 13776 2471 13832
rect 0 13774 2471 13776
rect 0 13744 800 13774
rect 2405 13771 2471 13774
rect 8845 13834 8911 13837
rect 11697 13834 11763 13837
rect 8845 13832 11763 13834
rect 8845 13776 8850 13832
rect 8906 13776 11702 13832
rect 11758 13776 11763 13832
rect 8845 13774 11763 13776
rect 8845 13771 8911 13774
rect 11697 13771 11763 13774
rect 3601 13698 3667 13701
rect 6310 13698 6316 13700
rect 3601 13696 6316 13698
rect 3601 13640 3606 13696
rect 3662 13640 6316 13696
rect 3601 13638 6316 13640
rect 3601 13635 3667 13638
rect 6310 13636 6316 13638
rect 6380 13636 6386 13700
rect 19200 13698 20000 13728
rect 17358 13638 20000 13698
rect 3170 13632 3486 13633
rect 0 13562 800 13592
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 16514 13567 16830 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 800 13502
rect 1853 13499 1919 13502
rect 5993 13426 6059 13429
rect 11421 13426 11487 13429
rect 5993 13424 11487 13426
rect 5993 13368 5998 13424
rect 6054 13368 11426 13424
rect 11482 13368 11487 13424
rect 5993 13366 11487 13368
rect 5993 13363 6059 13366
rect 11421 13363 11487 13366
rect 15469 13426 15535 13429
rect 17358 13426 17418 13638
rect 19200 13608 20000 13638
rect 19200 13426 20000 13456
rect 15469 13424 17418 13426
rect 15469 13368 15474 13424
rect 15530 13368 17418 13424
rect 15469 13366 17418 13368
rect 17542 13366 20000 13426
rect 15469 13363 15535 13366
rect 0 13290 800 13320
rect 1853 13290 1919 13293
rect 0 13288 1919 13290
rect 0 13232 1858 13288
rect 1914 13232 1919 13288
rect 0 13230 1919 13232
rect 0 13200 800 13230
rect 1853 13227 1919 13230
rect 2681 13290 2747 13293
rect 4102 13290 4108 13292
rect 2681 13288 4108 13290
rect 2681 13232 2686 13288
rect 2742 13232 4108 13288
rect 2681 13230 4108 13232
rect 2681 13227 2747 13230
rect 4102 13228 4108 13230
rect 4172 13228 4178 13292
rect 9213 13290 9279 13293
rect 10777 13290 10843 13293
rect 13905 13290 13971 13293
rect 9213 13288 13971 13290
rect 9213 13232 9218 13288
rect 9274 13232 10782 13288
rect 10838 13232 13910 13288
rect 13966 13232 13971 13288
rect 9213 13230 13971 13232
rect 9213 13227 9279 13230
rect 10777 13227 10843 13230
rect 13905 13227 13971 13230
rect 15193 13290 15259 13293
rect 17542 13290 17602 13366
rect 19200 13336 20000 13366
rect 15193 13288 17602 13290
rect 15193 13232 15198 13288
rect 15254 13232 17602 13288
rect 15193 13230 17602 13232
rect 15193 13227 15259 13230
rect 16246 13092 16252 13156
rect 16316 13154 16322 13156
rect 19200 13154 20000 13184
rect 16316 13094 20000 13154
rect 16316 13092 16322 13094
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 19200 13064 20000 13094
rect 14290 13023 14606 13024
rect 2405 13018 2471 13021
rect 0 13016 2471 13018
rect 0 12960 2410 13016
rect 2466 12960 2471 13016
rect 0 12958 2471 12960
rect 0 12928 800 12958
rect 2405 12955 2471 12958
rect 15377 12882 15443 12885
rect 19200 12882 20000 12912
rect 15377 12880 20000 12882
rect 15377 12824 15382 12880
rect 15438 12824 20000 12880
rect 15377 12822 20000 12824
rect 15377 12819 15443 12822
rect 19200 12792 20000 12822
rect 0 12746 800 12776
rect 2497 12746 2563 12749
rect 0 12744 2563 12746
rect 0 12688 2502 12744
rect 2558 12688 2563 12744
rect 0 12686 2563 12688
rect 0 12656 800 12686
rect 2497 12683 2563 12686
rect 14825 12746 14891 12749
rect 16573 12746 16639 12749
rect 14825 12744 16639 12746
rect 14825 12688 14830 12744
rect 14886 12688 16578 12744
rect 16634 12688 16639 12744
rect 14825 12686 16639 12688
rect 14825 12683 14891 12686
rect 16573 12683 16639 12686
rect 17769 12610 17835 12613
rect 19200 12610 20000 12640
rect 17769 12608 20000 12610
rect 17769 12552 17774 12608
rect 17830 12552 20000 12608
rect 17769 12550 20000 12552
rect 17769 12547 17835 12550
rect 3170 12544 3486 12545
rect 0 12474 800 12504
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 19200 12520 20000 12550
rect 16514 12479 16830 12480
rect 2773 12474 2839 12477
rect 0 12472 2839 12474
rect 0 12416 2778 12472
rect 2834 12416 2839 12472
rect 0 12414 2839 12416
rect 0 12384 800 12414
rect 2773 12411 2839 12414
rect 3509 12338 3575 12341
rect 12566 12338 12572 12340
rect 3509 12336 12572 12338
rect 3509 12280 3514 12336
rect 3570 12280 12572 12336
rect 3509 12278 12572 12280
rect 3509 12275 3575 12278
rect 12566 12276 12572 12278
rect 12636 12276 12642 12340
rect 19200 12338 20000 12368
rect 15518 12278 20000 12338
rect 0 12202 800 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 800 12142
rect 4061 12139 4127 12142
rect 4705 12202 4771 12205
rect 15377 12202 15443 12205
rect 4705 12200 15443 12202
rect 4705 12144 4710 12200
rect 4766 12144 15382 12200
rect 15438 12144 15443 12200
rect 4705 12142 15443 12144
rect 4705 12139 4771 12142
rect 15377 12139 15443 12142
rect 5394 12000 5710 12001
rect 0 11930 800 11960
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 14290 11935 14606 11936
rect 0 11870 2790 11930
rect 0 11840 800 11870
rect 2730 11794 2790 11870
rect 4153 11794 4219 11797
rect 4705 11794 4771 11797
rect 11145 11794 11211 11797
rect 13854 11794 13860 11796
rect 2730 11734 3986 11794
rect 0 11658 800 11688
rect 3785 11658 3851 11661
rect 0 11656 3851 11658
rect 0 11600 3790 11656
rect 3846 11600 3851 11656
rect 0 11598 3851 11600
rect 0 11568 800 11598
rect 3785 11595 3851 11598
rect 3926 11522 3986 11734
rect 4153 11792 11211 11794
rect 4153 11736 4158 11792
rect 4214 11736 4710 11792
rect 4766 11736 11150 11792
rect 11206 11736 11211 11792
rect 4153 11734 11211 11736
rect 4153 11731 4219 11734
rect 4705 11731 4771 11734
rect 11145 11731 11211 11734
rect 12390 11734 13860 11794
rect 4889 11658 4955 11661
rect 12390 11658 12450 11734
rect 13854 11732 13860 11734
rect 13924 11794 13930 11796
rect 15518 11794 15578 12278
rect 19200 12248 20000 12278
rect 18505 12066 18571 12069
rect 19200 12066 20000 12096
rect 18505 12064 20000 12066
rect 18505 12008 18510 12064
rect 18566 12008 20000 12064
rect 18505 12006 20000 12008
rect 18505 12003 18571 12006
rect 19200 11976 20000 12006
rect 13924 11734 15578 11794
rect 18781 11794 18847 11797
rect 19200 11794 20000 11824
rect 18781 11792 20000 11794
rect 18781 11736 18786 11792
rect 18842 11736 20000 11792
rect 18781 11734 20000 11736
rect 13924 11732 13930 11734
rect 18781 11731 18847 11734
rect 19200 11704 20000 11734
rect 4889 11656 12450 11658
rect 4889 11600 4894 11656
rect 4950 11600 12450 11656
rect 4889 11598 12450 11600
rect 15837 11658 15903 11661
rect 15837 11656 17050 11658
rect 15837 11600 15842 11656
rect 15898 11600 17050 11656
rect 15837 11598 17050 11600
rect 4889 11595 4955 11598
rect 15837 11595 15903 11598
rect 4061 11522 4127 11525
rect 11053 11524 11119 11525
rect 11053 11522 11100 11524
rect 3926 11520 4127 11522
rect 3926 11464 4066 11520
rect 4122 11464 4127 11520
rect 3926 11462 4127 11464
rect 11008 11520 11100 11522
rect 11164 11522 11170 11524
rect 11789 11522 11855 11525
rect 11164 11520 11855 11522
rect 11008 11464 11058 11520
rect 11164 11464 11794 11520
rect 11850 11464 11855 11520
rect 11008 11462 11100 11464
rect 4061 11459 4127 11462
rect 11053 11460 11100 11462
rect 11164 11462 11855 11464
rect 16990 11522 17050 11598
rect 19200 11522 20000 11552
rect 16990 11462 20000 11522
rect 11164 11460 11170 11462
rect 11053 11459 11119 11460
rect 11789 11459 11855 11462
rect 3170 11456 3486 11457
rect 0 11386 800 11416
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 19200 11432 20000 11462
rect 16514 11391 16830 11392
rect 1761 11386 1827 11389
rect 0 11384 1827 11386
rect 0 11328 1766 11384
rect 1822 11328 1827 11384
rect 0 11326 1827 11328
rect 0 11296 800 11326
rect 1761 11323 1827 11326
rect 6729 11250 6795 11253
rect 12893 11250 12959 11253
rect 6729 11248 12959 11250
rect 6729 11192 6734 11248
rect 6790 11192 12898 11248
rect 12954 11192 12959 11248
rect 6729 11190 12959 11192
rect 6729 11187 6795 11190
rect 12893 11187 12959 11190
rect 15929 11250 15995 11253
rect 19200 11250 20000 11280
rect 15929 11248 20000 11250
rect 15929 11192 15934 11248
rect 15990 11192 20000 11248
rect 15929 11190 20000 11192
rect 15929 11187 15995 11190
rect 19200 11160 20000 11190
rect 0 11114 800 11144
rect 8017 11114 8083 11117
rect 0 11112 8083 11114
rect 0 11056 8022 11112
rect 8078 11056 8083 11112
rect 0 11054 8083 11056
rect 0 11024 800 11054
rect 8017 11051 8083 11054
rect 17309 10978 17375 10981
rect 19200 10978 20000 11008
rect 17309 10976 20000 10978
rect 17309 10920 17314 10976
rect 17370 10920 20000 10976
rect 17309 10918 20000 10920
rect 17309 10915 17375 10918
rect 5394 10912 5710 10913
rect 0 10842 800 10872
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 19200 10888 20000 10918
rect 14290 10847 14606 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 2957 10706 3023 10709
rect 3509 10706 3575 10709
rect 1350 10704 3575 10706
rect 1350 10648 2962 10704
rect 3018 10648 3514 10704
rect 3570 10648 3575 10704
rect 1350 10646 3575 10648
rect 0 10570 800 10600
rect 1350 10570 1410 10646
rect 2957 10643 3023 10646
rect 3509 10643 3575 10646
rect 3969 10706 4035 10709
rect 9213 10706 9279 10709
rect 3969 10704 9279 10706
rect 3969 10648 3974 10704
rect 4030 10648 9218 10704
rect 9274 10648 9279 10704
rect 3969 10646 9279 10648
rect 3969 10643 4035 10646
rect 9213 10643 9279 10646
rect 15285 10706 15351 10709
rect 19200 10706 20000 10736
rect 15285 10704 20000 10706
rect 15285 10648 15290 10704
rect 15346 10648 20000 10704
rect 15285 10646 20000 10648
rect 15285 10643 15351 10646
rect 19200 10616 20000 10646
rect 0 10510 1410 10570
rect 2589 10570 2655 10573
rect 8385 10570 8451 10573
rect 11421 10570 11487 10573
rect 2589 10568 8080 10570
rect 2589 10512 2594 10568
rect 2650 10512 8080 10568
rect 2589 10510 8080 10512
rect 0 10480 800 10510
rect 2589 10507 2655 10510
rect 2313 10434 2379 10437
rect 2957 10434 3023 10437
rect 2313 10432 3023 10434
rect 2313 10376 2318 10432
rect 2374 10376 2962 10432
rect 3018 10376 3023 10432
rect 2313 10374 3023 10376
rect 8020 10434 8080 10510
rect 8385 10568 11487 10570
rect 8385 10512 8390 10568
rect 8446 10512 11426 10568
rect 11482 10512 11487 10568
rect 8385 10510 11487 10512
rect 8385 10507 8451 10510
rect 11421 10507 11487 10510
rect 8845 10434 8911 10437
rect 19200 10434 20000 10464
rect 8020 10432 8911 10434
rect 8020 10376 8850 10432
rect 8906 10376 8911 10432
rect 8020 10374 8911 10376
rect 2313 10371 2379 10374
rect 2957 10371 3023 10374
rect 8845 10371 8911 10374
rect 16990 10374 20000 10434
rect 3170 10368 3486 10369
rect 0 10298 800 10328
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 16514 10303 16830 10304
rect 0 10238 2790 10298
rect 0 10208 800 10238
rect 2730 10162 2790 10238
rect 6177 10162 6243 10165
rect 2730 10160 6243 10162
rect 2730 10104 6182 10160
rect 6238 10104 6243 10160
rect 2730 10102 6243 10104
rect 6177 10099 6243 10102
rect 10041 10162 10107 10165
rect 11421 10162 11487 10165
rect 10041 10160 11487 10162
rect 10041 10104 10046 10160
rect 10102 10104 11426 10160
rect 11482 10104 11487 10160
rect 10041 10102 11487 10104
rect 10041 10099 10107 10102
rect 11421 10099 11487 10102
rect 15009 10162 15075 10165
rect 16990 10162 17050 10374
rect 19200 10344 20000 10374
rect 19200 10162 20000 10192
rect 15009 10160 17050 10162
rect 15009 10104 15014 10160
rect 15070 10104 17050 10160
rect 15009 10102 17050 10104
rect 17772 10102 20000 10162
rect 15009 10099 15075 10102
rect 0 10026 800 10056
rect 17772 10029 17832 10102
rect 19200 10072 20000 10102
rect 4061 10026 4127 10029
rect 6729 10026 6795 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 800 9966
rect 4061 9963 4127 9966
rect 5214 10024 6795 10026
rect 5214 9968 6734 10024
rect 6790 9968 6795 10024
rect 5214 9966 6795 9968
rect 2589 9890 2655 9893
rect 5214 9890 5274 9966
rect 6729 9963 6795 9966
rect 8753 10026 8819 10029
rect 13670 10026 13676 10028
rect 8753 10024 13676 10026
rect 8753 9968 8758 10024
rect 8814 9968 13676 10024
rect 8753 9966 13676 9968
rect 8753 9963 8819 9966
rect 13670 9964 13676 9966
rect 13740 10026 13746 10028
rect 15653 10026 15719 10029
rect 13740 10024 15719 10026
rect 13740 9968 15658 10024
rect 15714 9968 15719 10024
rect 13740 9966 15719 9968
rect 13740 9964 13746 9966
rect 15653 9963 15719 9966
rect 17769 10024 17835 10029
rect 17769 9968 17774 10024
rect 17830 9968 17835 10024
rect 17769 9963 17835 9968
rect 2589 9888 5274 9890
rect 2589 9832 2594 9888
rect 2650 9832 5274 9888
rect 2589 9830 5274 9832
rect 10225 9890 10291 9893
rect 10685 9890 10751 9893
rect 10225 9888 10751 9890
rect 10225 9832 10230 9888
rect 10286 9832 10690 9888
rect 10746 9832 10751 9888
rect 10225 9830 10751 9832
rect 2589 9827 2655 9830
rect 10225 9827 10291 9830
rect 10685 9827 10751 9830
rect 15929 9890 15995 9893
rect 19200 9890 20000 9920
rect 15929 9888 20000 9890
rect 15929 9832 15934 9888
rect 15990 9832 20000 9888
rect 15929 9830 20000 9832
rect 15929 9827 15995 9830
rect 5394 9824 5710 9825
rect 0 9754 800 9784
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 19200 9800 20000 9830
rect 14290 9759 14606 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 2957 9754 3023 9757
rect 3509 9754 3575 9757
rect 13445 9754 13511 9757
rect 2957 9752 3575 9754
rect 2957 9696 2962 9752
rect 3018 9696 3514 9752
rect 3570 9696 3575 9752
rect 2957 9694 3575 9696
rect 2957 9691 3023 9694
rect 3509 9691 3575 9694
rect 10320 9752 13511 9754
rect 10320 9696 13450 9752
rect 13506 9696 13511 9752
rect 10320 9694 13511 9696
rect 10133 9690 10199 9693
rect 10320 9690 10380 9694
rect 13445 9691 13511 9694
rect 10133 9688 10380 9690
rect 10133 9632 10138 9688
rect 10194 9632 10380 9688
rect 10133 9630 10380 9632
rect 10133 9627 10199 9630
rect 2078 9556 2084 9620
rect 2148 9618 2154 9620
rect 3693 9618 3759 9621
rect 2148 9616 3759 9618
rect 2148 9560 3698 9616
rect 3754 9560 3759 9616
rect 2148 9558 3759 9560
rect 2148 9556 2154 9558
rect 3693 9555 3759 9558
rect 12985 9618 13051 9621
rect 15285 9618 15351 9621
rect 12985 9616 15351 9618
rect 12985 9560 12990 9616
rect 13046 9560 15290 9616
rect 15346 9560 15351 9616
rect 12985 9558 15351 9560
rect 12985 9555 13051 9558
rect 15285 9555 15351 9558
rect 16982 9556 16988 9620
rect 17052 9618 17058 9620
rect 17125 9618 17191 9621
rect 17052 9616 17191 9618
rect 17052 9560 17130 9616
rect 17186 9560 17191 9616
rect 17052 9558 17191 9560
rect 17052 9556 17058 9558
rect 17125 9555 17191 9558
rect 17401 9618 17467 9621
rect 19200 9618 20000 9648
rect 17401 9616 20000 9618
rect 17401 9560 17406 9616
rect 17462 9560 20000 9616
rect 17401 9558 20000 9560
rect 17401 9555 17467 9558
rect 19200 9528 20000 9558
rect 0 9482 800 9512
rect 4613 9482 4679 9485
rect 0 9480 4679 9482
rect 0 9424 4618 9480
rect 4674 9424 4679 9480
rect 0 9422 4679 9424
rect 0 9392 800 9422
rect 4613 9419 4679 9422
rect 6177 9482 6243 9485
rect 10317 9482 10383 9485
rect 14825 9482 14891 9485
rect 6177 9480 8218 9482
rect 6177 9424 6182 9480
rect 6238 9424 8218 9480
rect 6177 9422 8218 9424
rect 6177 9419 6243 9422
rect 8158 9346 8218 9422
rect 10317 9480 14891 9482
rect 10317 9424 10322 9480
rect 10378 9424 14830 9480
rect 14886 9424 14891 9480
rect 10317 9422 14891 9424
rect 10317 9419 10383 9422
rect 14825 9419 14891 9422
rect 10869 9346 10935 9349
rect 8158 9344 10935 9346
rect 8158 9288 10874 9344
rect 10930 9288 10935 9344
rect 8158 9286 10935 9288
rect 10869 9283 10935 9286
rect 12934 9284 12940 9348
rect 13004 9346 13010 9348
rect 15377 9346 15443 9349
rect 13004 9344 15443 9346
rect 13004 9288 15382 9344
rect 15438 9288 15443 9344
rect 13004 9286 15443 9288
rect 13004 9284 13010 9286
rect 15377 9283 15443 9286
rect 17493 9346 17559 9349
rect 19200 9346 20000 9376
rect 17493 9344 20000 9346
rect 17493 9288 17498 9344
rect 17554 9288 20000 9344
rect 17493 9286 20000 9288
rect 17493 9283 17559 9286
rect 3170 9280 3486 9281
rect 0 9210 800 9240
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 19200 9256 20000 9286
rect 16514 9215 16830 9216
rect 2957 9210 3023 9213
rect 4061 9210 4127 9213
rect 0 9208 3023 9210
rect 0 9152 2962 9208
rect 3018 9152 3023 9208
rect 0 9150 3023 9152
rect 0 9120 800 9150
rect 2957 9147 3023 9150
rect 3926 9208 4127 9210
rect 3926 9152 4066 9208
rect 4122 9152 4127 9208
rect 3926 9150 4127 9152
rect 3926 9077 3986 9150
rect 4061 9147 4127 9150
rect 10041 9210 10107 9213
rect 10358 9210 10364 9212
rect 10041 9208 10364 9210
rect 10041 9152 10046 9208
rect 10102 9152 10364 9208
rect 10041 9150 10364 9152
rect 10041 9147 10107 9150
rect 10358 9148 10364 9150
rect 10428 9148 10434 9212
rect 13261 9210 13327 9213
rect 15561 9210 15627 9213
rect 13261 9208 15627 9210
rect 13261 9152 13266 9208
rect 13322 9152 15566 9208
rect 15622 9152 15627 9208
rect 13261 9150 15627 9152
rect 13261 9147 13327 9150
rect 15561 9147 15627 9150
rect 3877 9072 3986 9077
rect 3877 9016 3882 9072
rect 3938 9016 3986 9072
rect 3877 9014 3986 9016
rect 5901 9074 5967 9077
rect 13353 9074 13419 9077
rect 5901 9072 13419 9074
rect 5901 9016 5906 9072
rect 5962 9016 13358 9072
rect 13414 9016 13419 9072
rect 5901 9014 13419 9016
rect 3877 9011 3943 9014
rect 5901 9011 5967 9014
rect 13353 9011 13419 9014
rect 18321 9074 18387 9077
rect 19200 9074 20000 9104
rect 18321 9072 20000 9074
rect 18321 9016 18326 9072
rect 18382 9016 20000 9072
rect 18321 9014 20000 9016
rect 18321 9011 18387 9014
rect 19200 8984 20000 9014
rect 0 8938 800 8968
rect 1945 8938 2011 8941
rect 0 8936 2011 8938
rect 0 8880 1950 8936
rect 2006 8880 2011 8936
rect 0 8878 2011 8880
rect 0 8848 800 8878
rect 1945 8875 2011 8878
rect 2262 8876 2268 8940
rect 2332 8938 2338 8940
rect 4429 8938 4495 8941
rect 2332 8936 4495 8938
rect 2332 8880 4434 8936
rect 4490 8880 4495 8936
rect 2332 8878 4495 8880
rect 2332 8876 2338 8878
rect 4429 8875 4495 8878
rect 6545 8938 6611 8941
rect 13445 8938 13511 8941
rect 6545 8936 13511 8938
rect 6545 8880 6550 8936
rect 6606 8880 13450 8936
rect 13506 8880 13511 8936
rect 6545 8878 13511 8880
rect 6545 8875 6611 8878
rect 13445 8875 13511 8878
rect 2681 8802 2747 8805
rect 5073 8802 5139 8805
rect 2681 8800 5139 8802
rect 2681 8744 2686 8800
rect 2742 8744 5078 8800
rect 5134 8744 5139 8800
rect 2681 8742 5139 8744
rect 2681 8739 2747 8742
rect 5073 8739 5139 8742
rect 6821 8802 6887 8805
rect 9029 8802 9095 8805
rect 13997 8802 14063 8805
rect 6821 8800 9095 8802
rect 6821 8744 6826 8800
rect 6882 8744 9034 8800
rect 9090 8744 9095 8800
rect 6821 8742 9095 8744
rect 6821 8739 6887 8742
rect 9029 8739 9095 8742
rect 12390 8800 14063 8802
rect 12390 8744 14002 8800
rect 14058 8744 14063 8800
rect 12390 8742 14063 8744
rect 5394 8736 5710 8737
rect 0 8666 800 8696
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 4061 8666 4127 8669
rect 12390 8666 12450 8742
rect 13997 8739 14063 8742
rect 18045 8802 18111 8805
rect 19200 8802 20000 8832
rect 18045 8800 20000 8802
rect 18045 8744 18050 8800
rect 18106 8744 20000 8800
rect 18045 8742 20000 8744
rect 18045 8739 18111 8742
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 15009 8666 15075 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 800 8606
rect 4061 8603 4127 8606
rect 10366 8606 12450 8666
rect 14966 8664 15075 8666
rect 14966 8608 15014 8664
rect 15070 8608 15075 8664
rect 4153 8530 4219 8533
rect 6177 8530 6243 8533
rect 4153 8528 6243 8530
rect 4153 8472 4158 8528
rect 4214 8472 6182 8528
rect 6238 8472 6243 8528
rect 4153 8470 6243 8472
rect 4153 8467 4219 8470
rect 6177 8467 6243 8470
rect 6729 8530 6795 8533
rect 10366 8530 10426 8606
rect 14966 8603 15075 8608
rect 6729 8528 10426 8530
rect 6729 8472 6734 8528
rect 6790 8472 10426 8528
rect 6729 8470 10426 8472
rect 10869 8530 10935 8533
rect 14966 8530 15026 8603
rect 10869 8528 15026 8530
rect 10869 8472 10874 8528
rect 10930 8472 15026 8528
rect 10869 8470 15026 8472
rect 16941 8530 17007 8533
rect 19200 8530 20000 8560
rect 16941 8528 20000 8530
rect 16941 8472 16946 8528
rect 17002 8472 20000 8528
rect 16941 8470 20000 8472
rect 6729 8467 6795 8470
rect 10869 8467 10935 8470
rect 16941 8467 17007 8470
rect 19200 8440 20000 8470
rect 0 8394 800 8424
rect 2957 8394 3023 8397
rect 0 8392 3023 8394
rect 0 8336 2962 8392
rect 3018 8336 3023 8392
rect 0 8334 3023 8336
rect 0 8304 800 8334
rect 2957 8331 3023 8334
rect 3693 8394 3759 8397
rect 4102 8394 4108 8396
rect 3693 8392 4108 8394
rect 3693 8336 3698 8392
rect 3754 8336 4108 8392
rect 3693 8334 4108 8336
rect 3693 8331 3759 8334
rect 4102 8332 4108 8334
rect 4172 8332 4178 8396
rect 4337 8394 4403 8397
rect 4981 8394 5047 8397
rect 13445 8394 13511 8397
rect 15377 8394 15443 8397
rect 4337 8392 13370 8394
rect 4337 8336 4342 8392
rect 4398 8336 4986 8392
rect 5042 8336 13370 8392
rect 4337 8334 13370 8336
rect 4337 8331 4403 8334
rect 4981 8331 5047 8334
rect 13310 8258 13370 8334
rect 13445 8392 15443 8394
rect 13445 8336 13450 8392
rect 13506 8336 15382 8392
rect 15438 8336 15443 8392
rect 13445 8334 15443 8336
rect 13445 8331 13511 8334
rect 15377 8331 15443 8334
rect 15193 8258 15259 8261
rect 13310 8256 15259 8258
rect 13310 8200 15198 8256
rect 15254 8200 15259 8256
rect 13310 8198 15259 8200
rect 15193 8195 15259 8198
rect 18137 8258 18203 8261
rect 19200 8258 20000 8288
rect 18137 8256 20000 8258
rect 18137 8200 18142 8256
rect 18198 8200 20000 8256
rect 18137 8198 20000 8200
rect 18137 8195 18203 8198
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 19200 8168 20000 8198
rect 16514 8127 16830 8128
rect 2865 8122 2931 8125
rect 0 8120 2931 8122
rect 0 8064 2870 8120
rect 2926 8064 2931 8120
rect 0 8062 2931 8064
rect 0 8032 800 8062
rect 2865 8059 2931 8062
rect 8109 8124 8175 8125
rect 8109 8120 8156 8124
rect 8220 8122 8226 8124
rect 8109 8064 8114 8120
rect 8109 8060 8156 8064
rect 8220 8062 8266 8122
rect 8220 8060 8226 8062
rect 8109 8059 8175 8060
rect 2681 7986 2747 7989
rect 2814 7986 2820 7988
rect 2681 7984 2820 7986
rect 2681 7928 2686 7984
rect 2742 7928 2820 7984
rect 2681 7926 2820 7928
rect 2681 7923 2747 7926
rect 2814 7924 2820 7926
rect 2884 7986 2890 7988
rect 3417 7986 3483 7989
rect 2884 7984 3483 7986
rect 2884 7928 3422 7984
rect 3478 7928 3483 7984
rect 2884 7926 3483 7928
rect 2884 7924 2890 7926
rect 3417 7923 3483 7926
rect 7833 7986 7899 7989
rect 10317 7986 10383 7989
rect 7833 7984 10383 7986
rect 7833 7928 7838 7984
rect 7894 7928 10322 7984
rect 10378 7928 10383 7984
rect 7833 7926 10383 7928
rect 7833 7923 7899 7926
rect 10317 7923 10383 7926
rect 10685 7986 10751 7989
rect 12985 7986 13051 7989
rect 10685 7984 13051 7986
rect 10685 7928 10690 7984
rect 10746 7928 12990 7984
rect 13046 7928 13051 7984
rect 10685 7926 13051 7928
rect 10685 7923 10751 7926
rect 12985 7923 13051 7926
rect 13997 7986 14063 7989
rect 14457 7986 14523 7989
rect 15142 7986 15148 7988
rect 13997 7984 15148 7986
rect 13997 7928 14002 7984
rect 14058 7928 14462 7984
rect 14518 7928 15148 7984
rect 13997 7926 15148 7928
rect 13997 7923 14063 7926
rect 14457 7923 14523 7926
rect 15142 7924 15148 7926
rect 15212 7924 15218 7988
rect 17350 7924 17356 7988
rect 17420 7986 17426 7988
rect 17493 7986 17559 7989
rect 17420 7984 17559 7986
rect 17420 7928 17498 7984
rect 17554 7928 17559 7984
rect 17420 7926 17559 7928
rect 17420 7924 17426 7926
rect 17493 7923 17559 7926
rect 18413 7986 18479 7989
rect 19200 7986 20000 8016
rect 18413 7984 20000 7986
rect 18413 7928 18418 7984
rect 18474 7928 20000 7984
rect 18413 7926 20000 7928
rect 18413 7923 18479 7926
rect 19200 7896 20000 7926
rect 0 7850 800 7880
rect 3509 7850 3575 7853
rect 0 7848 3575 7850
rect 0 7792 3514 7848
rect 3570 7792 3575 7848
rect 0 7790 3575 7792
rect 0 7760 800 7790
rect 3509 7787 3575 7790
rect 3877 7850 3943 7853
rect 12893 7850 12959 7853
rect 16573 7850 16639 7853
rect 3877 7848 12959 7850
rect 3877 7792 3882 7848
rect 3938 7792 12898 7848
rect 12954 7792 12959 7848
rect 3877 7790 12959 7792
rect 3877 7787 3943 7790
rect 12893 7787 12959 7790
rect 14046 7848 16639 7850
rect 14046 7792 16578 7848
rect 16634 7792 16639 7848
rect 14046 7790 16639 7792
rect 11697 7714 11763 7717
rect 14046 7714 14106 7790
rect 16116 7717 16176 7790
rect 16573 7787 16639 7790
rect 11697 7712 14106 7714
rect 11697 7656 11702 7712
rect 11758 7656 14106 7712
rect 11697 7654 14106 7656
rect 16113 7712 16179 7717
rect 16113 7656 16118 7712
rect 16174 7656 16179 7712
rect 11697 7651 11763 7654
rect 16113 7651 16179 7656
rect 16481 7714 16547 7717
rect 19200 7714 20000 7744
rect 16481 7712 20000 7714
rect 16481 7656 16486 7712
rect 16542 7656 20000 7712
rect 16481 7654 20000 7656
rect 16481 7651 16547 7654
rect 5394 7648 5710 7649
rect 0 7578 800 7608
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 19200 7624 20000 7654
rect 14290 7583 14606 7584
rect 2405 7578 2471 7581
rect 0 7576 2471 7578
rect 0 7520 2410 7576
rect 2466 7520 2471 7576
rect 0 7518 2471 7520
rect 0 7488 800 7518
rect 2405 7515 2471 7518
rect 3601 7578 3667 7581
rect 5073 7578 5139 7581
rect 3601 7576 5139 7578
rect 3601 7520 3606 7576
rect 3662 7520 5078 7576
rect 5134 7520 5139 7576
rect 3601 7518 5139 7520
rect 3601 7515 3667 7518
rect 5073 7515 5139 7518
rect 7230 7516 7236 7580
rect 7300 7578 7306 7580
rect 7557 7578 7623 7581
rect 7300 7576 7623 7578
rect 7300 7520 7562 7576
rect 7618 7520 7623 7576
rect 7300 7518 7623 7520
rect 7300 7516 7306 7518
rect 7557 7515 7623 7518
rect 15561 7578 15627 7581
rect 16849 7578 16915 7581
rect 15561 7576 16915 7578
rect 15561 7520 15566 7576
rect 15622 7520 16854 7576
rect 16910 7520 16915 7576
rect 15561 7518 16915 7520
rect 15561 7515 15627 7518
rect 16849 7515 16915 7518
rect 2865 7442 2931 7445
rect 3049 7442 3115 7445
rect 10685 7442 10751 7445
rect 2865 7440 10751 7442
rect 2865 7384 2870 7440
rect 2926 7384 3054 7440
rect 3110 7384 10690 7440
rect 10746 7384 10751 7440
rect 2865 7382 10751 7384
rect 2865 7379 2931 7382
rect 3049 7379 3115 7382
rect 10685 7379 10751 7382
rect 14733 7442 14799 7445
rect 17677 7442 17743 7445
rect 14733 7440 17743 7442
rect 14733 7384 14738 7440
rect 14794 7384 17682 7440
rect 17738 7384 17743 7440
rect 14733 7382 17743 7384
rect 14733 7379 14799 7382
rect 17677 7379 17743 7382
rect 18045 7442 18111 7445
rect 19200 7442 20000 7472
rect 18045 7440 20000 7442
rect 18045 7384 18050 7440
rect 18106 7384 20000 7440
rect 18045 7382 20000 7384
rect 18045 7379 18111 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 3233 7306 3299 7309
rect 3877 7306 3943 7309
rect 4153 7306 4219 7309
rect 3233 7304 3664 7306
rect 3233 7248 3238 7304
rect 3294 7248 3664 7304
rect 3233 7246 3664 7248
rect 3233 7243 3299 7246
rect 3604 7173 3664 7246
rect 3877 7304 4219 7306
rect 3877 7248 3882 7304
rect 3938 7248 4158 7304
rect 4214 7248 4219 7304
rect 3877 7246 4219 7248
rect 3877 7243 3943 7246
rect 4153 7243 4219 7246
rect 6545 7306 6611 7309
rect 7005 7306 7071 7309
rect 8845 7306 8911 7309
rect 12566 7306 12572 7308
rect 6545 7304 7071 7306
rect 6545 7248 6550 7304
rect 6606 7248 7010 7304
rect 7066 7248 7071 7304
rect 6545 7246 7071 7248
rect 6545 7243 6611 7246
rect 7005 7243 7071 7246
rect 7422 7246 8770 7306
rect 3601 7168 3667 7173
rect 3601 7112 3606 7168
rect 3662 7112 3667 7168
rect 3601 7107 3667 7112
rect 6177 7170 6243 7173
rect 7230 7170 7236 7172
rect 6177 7168 7236 7170
rect 6177 7112 6182 7168
rect 6238 7112 7236 7168
rect 6177 7110 7236 7112
rect 6177 7107 6243 7110
rect 7230 7108 7236 7110
rect 7300 7108 7306 7172
rect 3170 7104 3486 7105
rect 0 7034 800 7064
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 1301 7034 1367 7037
rect 0 7032 1367 7034
rect 0 6976 1306 7032
rect 1362 6976 1367 7032
rect 0 6974 1367 6976
rect 0 6944 800 6974
rect 1301 6971 1367 6974
rect 3785 7034 3851 7037
rect 7189 7034 7255 7037
rect 7422 7034 7482 7246
rect 8710 7170 8770 7246
rect 8845 7304 12572 7306
rect 8845 7248 8850 7304
rect 8906 7248 12572 7304
rect 8845 7246 12572 7248
rect 8845 7243 8911 7246
rect 12566 7244 12572 7246
rect 12636 7306 12642 7308
rect 17769 7306 17835 7309
rect 12636 7304 17835 7306
rect 12636 7248 17774 7304
rect 17830 7248 17835 7304
rect 12636 7246 17835 7248
rect 12636 7244 12642 7246
rect 17769 7243 17835 7246
rect 11697 7170 11763 7173
rect 8710 7168 11763 7170
rect 8710 7112 11702 7168
rect 11758 7112 11763 7168
rect 8710 7110 11763 7112
rect 11697 7107 11763 7110
rect 18505 7170 18571 7173
rect 19200 7170 20000 7200
rect 18505 7168 20000 7170
rect 18505 7112 18510 7168
rect 18566 7112 20000 7168
rect 18505 7110 20000 7112
rect 18505 7107 18571 7110
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 18689 7034 18755 7037
rect 3785 7032 7482 7034
rect 3785 6976 3790 7032
rect 3846 6976 7194 7032
rect 7250 6976 7482 7032
rect 3785 6974 7482 6976
rect 18462 7032 18755 7034
rect 18462 6976 18694 7032
rect 18750 6976 18755 7032
rect 18462 6974 18755 6976
rect 3785 6971 3851 6974
rect 7189 6971 7255 6974
rect 1577 6898 1643 6901
rect 3141 6898 3207 6901
rect 3877 6898 3943 6901
rect 8937 6898 9003 6901
rect 17861 6898 17927 6901
rect 1577 6896 1962 6898
rect 1577 6840 1582 6896
rect 1638 6840 1962 6896
rect 1577 6838 1962 6840
rect 1577 6835 1643 6838
rect 0 6762 800 6792
rect 1669 6762 1735 6765
rect 0 6760 1735 6762
rect 0 6704 1674 6760
rect 1730 6704 1735 6760
rect 0 6702 1735 6704
rect 1902 6762 1962 6838
rect 3141 6896 9003 6898
rect 3141 6840 3146 6896
rect 3202 6840 3882 6896
rect 3938 6840 8942 6896
rect 8998 6840 9003 6896
rect 3141 6838 9003 6840
rect 3141 6835 3207 6838
rect 3877 6835 3943 6838
rect 8937 6835 9003 6838
rect 10182 6896 17927 6898
rect 10182 6840 17866 6896
rect 17922 6840 17927 6896
rect 10182 6838 17927 6840
rect 10182 6765 10242 6838
rect 17861 6835 17927 6838
rect 8937 6762 9003 6765
rect 10133 6762 10242 6765
rect 16246 6762 16252 6764
rect 1902 6760 10242 6762
rect 1902 6704 8942 6760
rect 8998 6704 10138 6760
rect 10194 6704 10242 6760
rect 1902 6702 10242 6704
rect 10366 6702 16252 6762
rect 0 6672 800 6702
rect 1669 6699 1735 6702
rect 8937 6699 9003 6702
rect 10133 6699 10199 6702
rect 1301 6626 1367 6629
rect 5257 6626 5323 6629
rect 1301 6624 5323 6626
rect 1301 6568 1306 6624
rect 1362 6568 5262 6624
rect 5318 6568 5323 6624
rect 1301 6566 5323 6568
rect 1301 6563 1367 6566
rect 5257 6563 5323 6566
rect 7741 6626 7807 6629
rect 8150 6626 8156 6628
rect 7741 6624 8156 6626
rect 7741 6568 7746 6624
rect 7802 6568 8156 6624
rect 7741 6566 8156 6568
rect 7741 6563 7807 6566
rect 8150 6564 8156 6566
rect 8220 6564 8226 6628
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 5809 6490 5875 6493
rect 8017 6490 8083 6493
rect 9397 6490 9463 6493
rect 0 6430 2790 6490
rect 0 6400 800 6430
rect 1945 6354 2011 6357
rect 2078 6354 2084 6356
rect 1945 6352 2084 6354
rect 1945 6296 1950 6352
rect 2006 6296 2084 6352
rect 1945 6294 2084 6296
rect 1945 6291 2011 6294
rect 2078 6292 2084 6294
rect 2148 6292 2154 6356
rect 2730 6354 2790 6430
rect 5809 6488 9463 6490
rect 5809 6432 5814 6488
rect 5870 6432 8022 6488
rect 8078 6432 9402 6488
rect 9458 6432 9463 6488
rect 5809 6430 9463 6432
rect 5809 6427 5875 6430
rect 8017 6427 8083 6430
rect 9397 6427 9463 6430
rect 2957 6354 3023 6357
rect 2730 6352 3023 6354
rect 2730 6296 2962 6352
rect 3018 6296 3023 6352
rect 2730 6294 3023 6296
rect 2957 6291 3023 6294
rect 6453 6354 6519 6357
rect 8385 6354 8451 6357
rect 6453 6352 8451 6354
rect 6453 6296 6458 6352
rect 6514 6296 8390 6352
rect 8446 6296 8451 6352
rect 6453 6294 8451 6296
rect 6453 6291 6519 6294
rect 8385 6291 8451 6294
rect 8753 6354 8819 6357
rect 10366 6354 10426 6702
rect 16246 6700 16252 6702
rect 16316 6700 16322 6764
rect 16757 6762 16823 6765
rect 18321 6762 18387 6765
rect 18462 6762 18522 6974
rect 18689 6971 18755 6974
rect 18689 6898 18755 6901
rect 19200 6898 20000 6928
rect 18689 6896 20000 6898
rect 18689 6840 18694 6896
rect 18750 6840 20000 6896
rect 18689 6838 20000 6840
rect 18689 6835 18755 6838
rect 19200 6808 20000 6838
rect 16757 6760 18522 6762
rect 16757 6704 16762 6760
rect 16818 6704 18326 6760
rect 18382 6704 18522 6760
rect 16757 6702 18522 6704
rect 16757 6699 16823 6702
rect 18321 6699 18387 6702
rect 11881 6626 11947 6629
rect 13813 6628 13879 6629
rect 13813 6626 13860 6628
rect 11881 6624 13860 6626
rect 11881 6568 11886 6624
rect 11942 6568 13818 6624
rect 11881 6566 13860 6568
rect 11881 6563 11947 6566
rect 13813 6564 13860 6566
rect 13924 6564 13930 6628
rect 15837 6626 15903 6629
rect 17769 6626 17835 6629
rect 15837 6624 17835 6626
rect 15837 6568 15842 6624
rect 15898 6568 17774 6624
rect 17830 6568 17835 6624
rect 15837 6566 17835 6568
rect 13813 6563 13879 6564
rect 15837 6563 15903 6566
rect 17769 6563 17835 6566
rect 18597 6626 18663 6629
rect 19200 6626 20000 6656
rect 18597 6624 20000 6626
rect 18597 6568 18602 6624
rect 18658 6568 20000 6624
rect 18597 6566 20000 6568
rect 18597 6563 18663 6566
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 19200 6536 20000 6566
rect 14290 6495 14606 6496
rect 12617 6492 12683 6493
rect 12566 6428 12572 6492
rect 12636 6490 12683 6492
rect 16481 6490 16547 6493
rect 18781 6490 18847 6493
rect 12636 6488 12728 6490
rect 12678 6432 12728 6488
rect 12636 6430 12728 6432
rect 16481 6488 18847 6490
rect 16481 6432 16486 6488
rect 16542 6432 18786 6488
rect 18842 6432 18847 6488
rect 16481 6430 18847 6432
rect 12636 6428 12683 6430
rect 12617 6427 12683 6428
rect 16481 6427 16547 6430
rect 18781 6427 18847 6430
rect 8753 6352 10426 6354
rect 8753 6296 8758 6352
rect 8814 6296 10426 6352
rect 8753 6294 10426 6296
rect 11145 6354 11211 6357
rect 16757 6354 16823 6357
rect 11145 6352 16823 6354
rect 11145 6296 11150 6352
rect 11206 6296 16762 6352
rect 16818 6296 16823 6352
rect 11145 6294 16823 6296
rect 8753 6291 8819 6294
rect 11145 6291 11211 6294
rect 16757 6291 16823 6294
rect 17677 6354 17743 6357
rect 19200 6354 20000 6384
rect 17677 6352 20000 6354
rect 17677 6296 17682 6352
rect 17738 6296 20000 6352
rect 17677 6294 20000 6296
rect 17677 6291 17743 6294
rect 19200 6264 20000 6294
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 2037 6218 2103 6221
rect 7741 6218 7807 6221
rect 15694 6218 15700 6220
rect 2037 6216 15700 6218
rect 2037 6160 2042 6216
rect 2098 6160 7746 6216
rect 7802 6160 15700 6216
rect 2037 6158 15700 6160
rect 2037 6155 2103 6158
rect 7741 6155 7807 6158
rect 15694 6156 15700 6158
rect 15764 6156 15770 6220
rect 18137 6082 18203 6085
rect 19200 6082 20000 6112
rect 18137 6080 20000 6082
rect 18137 6024 18142 6080
rect 18198 6024 20000 6080
rect 18137 6022 20000 6024
rect 18137 6019 18203 6022
rect 3170 6016 3486 6017
rect 0 5946 800 5976
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 19200 5992 20000 6022
rect 16514 5951 16830 5952
rect 2773 5946 2839 5949
rect 17309 5948 17375 5949
rect 17309 5946 17356 5948
rect 0 5944 2839 5946
rect 0 5888 2778 5944
rect 2834 5888 2839 5944
rect 0 5886 2839 5888
rect 17264 5944 17356 5946
rect 17264 5888 17314 5944
rect 17264 5886 17356 5888
rect 0 5856 800 5886
rect 2773 5883 2839 5886
rect 17309 5884 17356 5886
rect 17420 5884 17426 5948
rect 17309 5883 17375 5884
rect 11881 5810 11947 5813
rect 12566 5810 12572 5812
rect 11881 5808 12572 5810
rect 11881 5752 11886 5808
rect 11942 5752 12572 5808
rect 11881 5750 12572 5752
rect 11881 5747 11947 5750
rect 12566 5748 12572 5750
rect 12636 5810 12642 5812
rect 14181 5810 14247 5813
rect 15653 5812 15719 5813
rect 15653 5810 15700 5812
rect 12636 5808 14247 5810
rect 12636 5752 14186 5808
rect 14242 5752 14247 5808
rect 12636 5750 14247 5752
rect 15608 5808 15700 5810
rect 15608 5752 15658 5808
rect 15608 5750 15700 5752
rect 12636 5748 12642 5750
rect 14181 5747 14247 5750
rect 15653 5748 15700 5750
rect 15764 5748 15770 5812
rect 16246 5748 16252 5812
rect 16316 5810 16322 5812
rect 17033 5810 17099 5813
rect 16316 5808 17099 5810
rect 16316 5752 17038 5808
rect 17094 5752 17099 5808
rect 16316 5750 17099 5752
rect 16316 5748 16322 5750
rect 15653 5747 15719 5748
rect 17033 5747 17099 5750
rect 18229 5810 18295 5813
rect 19200 5810 20000 5840
rect 18229 5808 20000 5810
rect 18229 5752 18234 5808
rect 18290 5752 20000 5808
rect 18229 5750 20000 5752
rect 18229 5747 18295 5750
rect 19200 5720 20000 5750
rect 0 5674 800 5704
rect 1853 5674 1919 5677
rect 0 5672 1919 5674
rect 0 5616 1858 5672
rect 1914 5616 1919 5672
rect 0 5614 1919 5616
rect 0 5584 800 5614
rect 1853 5611 1919 5614
rect 4981 5674 5047 5677
rect 5533 5674 5599 5677
rect 4981 5672 5599 5674
rect 4981 5616 4986 5672
rect 5042 5616 5538 5672
rect 5594 5616 5599 5672
rect 4981 5614 5599 5616
rect 4981 5611 5047 5614
rect 5533 5611 5599 5614
rect 6729 5674 6795 5677
rect 9673 5674 9739 5677
rect 6729 5672 9739 5674
rect 6729 5616 6734 5672
rect 6790 5616 9678 5672
rect 9734 5616 9739 5672
rect 6729 5614 9739 5616
rect 6729 5611 6795 5614
rect 9673 5611 9739 5614
rect 10961 5674 11027 5677
rect 11237 5674 11303 5677
rect 10961 5672 11303 5674
rect 10961 5616 10966 5672
rect 11022 5616 11242 5672
rect 11298 5616 11303 5672
rect 10961 5614 11303 5616
rect 10961 5611 11027 5614
rect 11237 5611 11303 5614
rect 12525 5674 12591 5677
rect 18597 5674 18663 5677
rect 12525 5672 18663 5674
rect 12525 5616 12530 5672
rect 12586 5616 18602 5672
rect 18658 5616 18663 5672
rect 12525 5614 18663 5616
rect 12525 5611 12591 5614
rect 18597 5611 18663 5614
rect 6821 5538 6887 5541
rect 9305 5538 9371 5541
rect 6821 5536 9371 5538
rect 6821 5480 6826 5536
rect 6882 5480 9310 5536
rect 9366 5480 9371 5536
rect 6821 5478 9371 5480
rect 6821 5475 6887 5478
rect 9305 5475 9371 5478
rect 10409 5538 10475 5541
rect 12801 5538 12867 5541
rect 10409 5536 12867 5538
rect 10409 5480 10414 5536
rect 10470 5480 12806 5536
rect 12862 5480 12867 5536
rect 10409 5478 12867 5480
rect 10409 5475 10475 5478
rect 12801 5475 12867 5478
rect 14917 5538 14983 5541
rect 15469 5538 15535 5541
rect 14917 5536 15535 5538
rect 14917 5480 14922 5536
rect 14978 5480 15474 5536
rect 15530 5480 15535 5536
rect 14917 5478 15535 5480
rect 14917 5475 14983 5478
rect 15469 5475 15535 5478
rect 18321 5538 18387 5541
rect 19200 5538 20000 5568
rect 18321 5536 20000 5538
rect 18321 5480 18326 5536
rect 18382 5480 20000 5536
rect 18321 5478 20000 5480
rect 18321 5475 18387 5478
rect 5394 5472 5710 5473
rect 0 5402 800 5432
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 4061 5402 4127 5405
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 800 5342
rect 4061 5339 4127 5342
rect 7281 5402 7347 5405
rect 7557 5402 7623 5405
rect 7281 5400 7623 5402
rect 7281 5344 7286 5400
rect 7342 5344 7562 5400
rect 7618 5344 7623 5400
rect 7281 5342 7623 5344
rect 7281 5339 7347 5342
rect 7557 5339 7623 5342
rect 15193 5402 15259 5405
rect 17350 5402 17356 5404
rect 15193 5400 17356 5402
rect 15193 5344 15198 5400
rect 15254 5344 17356 5400
rect 15193 5342 17356 5344
rect 15193 5339 15259 5342
rect 17350 5340 17356 5342
rect 17420 5340 17426 5404
rect 17769 5402 17835 5405
rect 18873 5402 18939 5405
rect 17769 5400 18939 5402
rect 17769 5344 17774 5400
rect 17830 5344 18878 5400
rect 18934 5344 18939 5400
rect 17769 5342 18939 5344
rect 17769 5339 17835 5342
rect 18873 5339 18939 5342
rect 2773 5268 2839 5269
rect 2773 5264 2820 5268
rect 2884 5266 2890 5268
rect 3325 5266 3391 5269
rect 8845 5266 8911 5269
rect 2773 5208 2778 5264
rect 2773 5204 2820 5208
rect 2884 5206 2930 5266
rect 3325 5264 8911 5266
rect 3325 5208 3330 5264
rect 3386 5208 8850 5264
rect 8906 5208 8911 5264
rect 3325 5206 8911 5208
rect 2884 5204 2890 5206
rect 2773 5203 2839 5204
rect 3325 5203 3391 5206
rect 8845 5203 8911 5206
rect 9765 5266 9831 5269
rect 14089 5266 14155 5269
rect 9765 5264 14155 5266
rect 9765 5208 9770 5264
rect 9826 5208 14094 5264
rect 14150 5208 14155 5264
rect 9765 5206 14155 5208
rect 9765 5203 9831 5206
rect 14089 5203 14155 5206
rect 15285 5266 15351 5269
rect 19200 5266 20000 5296
rect 15285 5264 20000 5266
rect 15285 5208 15290 5264
rect 15346 5208 20000 5264
rect 15285 5206 20000 5208
rect 15285 5203 15351 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 2773 5130 2839 5133
rect 3417 5130 3483 5133
rect 10777 5130 10843 5133
rect 0 5128 2839 5130
rect 0 5072 2778 5128
rect 2834 5072 2839 5128
rect 0 5070 2839 5072
rect 0 5040 800 5070
rect 2773 5067 2839 5070
rect 2960 5128 10843 5130
rect 2960 5072 3422 5128
rect 3478 5072 10782 5128
rect 10838 5072 10843 5128
rect 2960 5070 10843 5072
rect 2037 4994 2103 4997
rect 2960 4994 3020 5070
rect 3417 5067 3483 5070
rect 10777 5067 10843 5070
rect 13629 5132 13695 5133
rect 13629 5128 13676 5132
rect 13740 5130 13746 5132
rect 15193 5130 15259 5133
rect 13629 5072 13634 5128
rect 13629 5068 13676 5072
rect 13740 5070 13786 5130
rect 15193 5128 17234 5130
rect 15193 5072 15198 5128
rect 15254 5072 17234 5128
rect 15193 5070 17234 5072
rect 13740 5068 13746 5070
rect 13629 5067 13695 5068
rect 15193 5067 15259 5070
rect 2037 4992 3020 4994
rect 2037 4936 2042 4992
rect 2098 4936 3020 4992
rect 2037 4934 3020 4936
rect 13261 4994 13327 4997
rect 15561 4994 15627 4997
rect 13261 4992 15627 4994
rect 13261 4936 13266 4992
rect 13322 4936 15566 4992
rect 15622 4936 15627 4992
rect 13261 4934 15627 4936
rect 17174 4994 17234 5070
rect 19200 4994 20000 5024
rect 17174 4934 20000 4994
rect 2037 4931 2103 4934
rect 13261 4931 13327 4934
rect 15561 4931 15627 4934
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 19200 4904 20000 4934
rect 16514 4863 16830 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 17217 4858 17283 4861
rect 17350 4858 17356 4860
rect 17217 4856 17356 4858
rect 17217 4800 17222 4856
rect 17278 4800 17356 4856
rect 17217 4798 17356 4800
rect 17217 4795 17283 4798
rect 17350 4796 17356 4798
rect 17420 4796 17426 4860
rect 7005 4722 7071 4725
rect 8201 4722 8267 4725
rect 10317 4724 10383 4725
rect 10317 4722 10364 4724
rect 7005 4720 8267 4722
rect 7005 4664 7010 4720
rect 7066 4664 8206 4720
rect 8262 4664 8267 4720
rect 7005 4662 8267 4664
rect 10272 4720 10364 4722
rect 10272 4664 10322 4720
rect 10272 4662 10364 4664
rect 7005 4659 7071 4662
rect 8201 4659 8267 4662
rect 10317 4660 10364 4662
rect 10428 4660 10434 4724
rect 13721 4722 13787 4725
rect 17769 4722 17835 4725
rect 13721 4720 17835 4722
rect 13721 4664 13726 4720
rect 13782 4664 17774 4720
rect 17830 4664 17835 4720
rect 13721 4662 17835 4664
rect 10317 4659 10383 4660
rect 13721 4659 13787 4662
rect 17769 4659 17835 4662
rect 18505 4722 18571 4725
rect 19200 4722 20000 4752
rect 18505 4720 20000 4722
rect 18505 4664 18510 4720
rect 18566 4664 20000 4720
rect 18505 4662 20000 4664
rect 18505 4659 18571 4662
rect 19200 4632 20000 4662
rect 0 4586 800 4616
rect 1853 4586 1919 4589
rect 0 4584 1919 4586
rect 0 4528 1858 4584
rect 1914 4528 1919 4584
rect 0 4526 1919 4528
rect 0 4496 800 4526
rect 1853 4523 1919 4526
rect 3141 4586 3207 4589
rect 3969 4586 4035 4589
rect 10685 4586 10751 4589
rect 17861 4586 17927 4589
rect 3141 4584 10426 4586
rect 3141 4528 3146 4584
rect 3202 4528 3974 4584
rect 4030 4528 10426 4584
rect 3141 4526 10426 4528
rect 3141 4523 3207 4526
rect 3969 4523 4035 4526
rect 10366 4450 10426 4526
rect 10685 4584 17927 4586
rect 10685 4528 10690 4584
rect 10746 4528 17866 4584
rect 17922 4528 17927 4584
rect 10685 4526 17927 4528
rect 10685 4523 10751 4526
rect 17861 4523 17927 4526
rect 13169 4450 13235 4453
rect 10366 4448 13235 4450
rect 10366 4392 13174 4448
rect 13230 4392 13235 4448
rect 10366 4390 13235 4392
rect 13169 4387 13235 4390
rect 14917 4450 14983 4453
rect 16757 4450 16823 4453
rect 14917 4448 16823 4450
rect 14917 4392 14922 4448
rect 14978 4392 16762 4448
rect 16818 4392 16823 4448
rect 14917 4390 16823 4392
rect 14917 4387 14983 4390
rect 16757 4387 16823 4390
rect 16941 4450 17007 4453
rect 19200 4450 20000 4480
rect 16941 4448 20000 4450
rect 16941 4392 16946 4448
rect 17002 4392 20000 4448
rect 16941 4390 20000 4392
rect 16941 4387 17007 4390
rect 5394 4384 5710 4385
rect 0 4314 800 4344
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 19200 4360 20000 4390
rect 14290 4319 14606 4320
rect 2221 4314 2287 4317
rect 0 4312 2287 4314
rect 0 4256 2226 4312
rect 2282 4256 2287 4312
rect 0 4254 2287 4256
rect 0 4224 800 4254
rect 2221 4251 2287 4254
rect 15142 4252 15148 4316
rect 15212 4314 15218 4316
rect 17953 4314 18019 4317
rect 15212 4312 18019 4314
rect 15212 4256 17958 4312
rect 18014 4256 18019 4312
rect 15212 4254 18019 4256
rect 15212 4252 15218 4254
rect 17953 4251 18019 4254
rect 3509 4178 3575 4181
rect 13721 4178 13787 4181
rect 3509 4176 13787 4178
rect 3509 4120 3514 4176
rect 3570 4120 13726 4176
rect 13782 4120 13787 4176
rect 3509 4118 13787 4120
rect 3509 4115 3575 4118
rect 13721 4115 13787 4118
rect 17309 4178 17375 4181
rect 19200 4178 20000 4208
rect 17309 4176 20000 4178
rect 17309 4120 17314 4176
rect 17370 4120 20000 4176
rect 17309 4118 20000 4120
rect 17309 4115 17375 4118
rect 19200 4088 20000 4118
rect 0 4042 800 4072
rect 2773 4042 2839 4045
rect 0 4040 2839 4042
rect 0 3984 2778 4040
rect 2834 3984 2839 4040
rect 0 3982 2839 3984
rect 0 3952 800 3982
rect 2773 3979 2839 3982
rect 4286 3980 4292 4044
rect 4356 4042 4362 4044
rect 10777 4042 10843 4045
rect 12801 4042 12867 4045
rect 12934 4042 12940 4044
rect 4356 4040 10843 4042
rect 4356 3984 10782 4040
rect 10838 3984 10843 4040
rect 4356 3982 10843 3984
rect 4356 3980 4362 3982
rect 10777 3979 10843 3982
rect 10918 3982 12634 4042
rect 2037 3906 2103 3909
rect 9029 3906 9095 3909
rect 10918 3906 10978 3982
rect 2037 3904 2790 3906
rect 2037 3848 2042 3904
rect 2098 3848 2790 3904
rect 2037 3846 2790 3848
rect 2037 3843 2103 3846
rect 0 3770 800 3800
rect 2405 3770 2471 3773
rect 0 3768 2471 3770
rect 0 3712 2410 3768
rect 2466 3712 2471 3768
rect 0 3710 2471 3712
rect 0 3680 800 3710
rect 2405 3707 2471 3710
rect 2129 3634 2195 3637
rect 2262 3634 2268 3636
rect 2129 3632 2268 3634
rect 2129 3576 2134 3632
rect 2190 3576 2268 3632
rect 2129 3574 2268 3576
rect 2129 3571 2195 3574
rect 2262 3572 2268 3574
rect 2332 3572 2338 3636
rect 2730 3634 2790 3846
rect 9029 3904 10978 3906
rect 9029 3848 9034 3904
rect 9090 3848 10978 3904
rect 9029 3846 10978 3848
rect 12574 3906 12634 3982
rect 12801 4040 12940 4042
rect 12801 3984 12806 4040
rect 12862 3984 12940 4040
rect 12801 3982 12940 3984
rect 12801 3979 12867 3982
rect 12934 3980 12940 3982
rect 13004 3980 13010 4044
rect 15377 4042 15443 4045
rect 16982 4042 16988 4044
rect 15377 4040 16988 4042
rect 15377 3984 15382 4040
rect 15438 3984 16988 4040
rect 15377 3982 16988 3984
rect 15377 3979 15443 3982
rect 16982 3980 16988 3982
rect 17052 3980 17058 4044
rect 15285 3906 15351 3909
rect 12574 3904 15351 3906
rect 12574 3848 15290 3904
rect 15346 3848 15351 3904
rect 12574 3846 15351 3848
rect 9029 3843 9095 3846
rect 15285 3843 15351 3846
rect 17401 3906 17467 3909
rect 19200 3906 20000 3936
rect 17401 3904 20000 3906
rect 17401 3848 17406 3904
rect 17462 3848 20000 3904
rect 17401 3846 20000 3848
rect 17401 3843 17467 3846
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 10501 3770 10567 3773
rect 8894 3768 10567 3770
rect 8894 3712 10506 3768
rect 10562 3712 10567 3768
rect 8894 3710 10567 3712
rect 8894 3634 8954 3710
rect 10501 3707 10567 3710
rect 2730 3574 8954 3634
rect 9070 3572 9076 3636
rect 9140 3634 9146 3636
rect 15469 3634 15535 3637
rect 9140 3632 15535 3634
rect 9140 3576 15474 3632
rect 15530 3576 15535 3632
rect 9140 3574 15535 3576
rect 9140 3572 9146 3574
rect 15469 3571 15535 3574
rect 15694 3572 15700 3636
rect 15764 3634 15770 3636
rect 16113 3634 16179 3637
rect 15764 3632 16179 3634
rect 15764 3576 16118 3632
rect 16174 3576 16179 3632
rect 15764 3574 16179 3576
rect 15764 3572 15770 3574
rect 16113 3571 16179 3574
rect 16246 3572 16252 3636
rect 16316 3634 16322 3636
rect 16573 3634 16639 3637
rect 16316 3632 16639 3634
rect 16316 3576 16578 3632
rect 16634 3576 16639 3632
rect 16316 3574 16639 3576
rect 16316 3572 16322 3574
rect 16573 3571 16639 3574
rect 18045 3634 18111 3637
rect 19200 3634 20000 3664
rect 18045 3632 20000 3634
rect 18045 3576 18050 3632
rect 18106 3576 20000 3632
rect 18045 3574 20000 3576
rect 18045 3571 18111 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 3049 3498 3115 3501
rect 11094 3498 11100 3500
rect 0 3496 3115 3498
rect 0 3440 3054 3496
rect 3110 3440 3115 3496
rect 0 3438 3115 3440
rect 0 3408 800 3438
rect 3049 3435 3115 3438
rect 6134 3438 11100 3498
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 3877 3226 3943 3229
rect 0 3224 3943 3226
rect 0 3168 3882 3224
rect 3938 3168 3943 3224
rect 0 3166 3943 3168
rect 0 3136 800 3166
rect 3877 3163 3943 3166
rect 1209 3090 1275 3093
rect 6134 3090 6194 3438
rect 11094 3436 11100 3438
rect 11164 3436 11170 3500
rect 17861 3362 17927 3365
rect 19200 3362 20000 3392
rect 17861 3360 20000 3362
rect 17861 3304 17866 3360
rect 17922 3304 20000 3360
rect 17861 3302 20000 3304
rect 17861 3299 17927 3302
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 19200 3272 20000 3302
rect 14290 3231 14606 3232
rect 15193 3226 15259 3229
rect 18137 3226 18203 3229
rect 15193 3224 18203 3226
rect 15193 3168 15198 3224
rect 15254 3168 18142 3224
rect 18198 3168 18203 3224
rect 15193 3166 18203 3168
rect 15193 3163 15259 3166
rect 18137 3163 18203 3166
rect 1209 3088 6194 3090
rect 1209 3032 1214 3088
rect 1270 3032 6194 3088
rect 1209 3030 6194 3032
rect 1209 3027 1275 3030
rect 6310 3028 6316 3092
rect 6380 3090 6386 3092
rect 15377 3090 15443 3093
rect 6380 3088 15443 3090
rect 6380 3032 15382 3088
rect 15438 3032 15443 3088
rect 6380 3030 15443 3032
rect 6380 3028 6386 3030
rect 15377 3027 15443 3030
rect 16297 3090 16363 3093
rect 17769 3090 17835 3093
rect 19200 3090 20000 3120
rect 16297 3088 17234 3090
rect 16297 3032 16302 3088
rect 16358 3032 17234 3088
rect 16297 3030 17234 3032
rect 16297 3027 16363 3030
rect 0 2954 800 2984
rect 2865 2954 2931 2957
rect 0 2952 2931 2954
rect 0 2896 2870 2952
rect 2926 2896 2931 2952
rect 0 2894 2931 2896
rect 0 2864 800 2894
rect 2865 2891 2931 2894
rect 4102 2892 4108 2956
rect 4172 2954 4178 2956
rect 16941 2954 17007 2957
rect 4172 2952 17007 2954
rect 4172 2896 16946 2952
rect 17002 2896 17007 2952
rect 4172 2894 17007 2896
rect 4172 2892 4178 2894
rect 16941 2891 17007 2894
rect 17174 2818 17234 3030
rect 17769 3088 20000 3090
rect 17769 3032 17774 3088
rect 17830 3032 20000 3088
rect 17769 3030 20000 3032
rect 17769 3027 17835 3030
rect 19200 3000 20000 3030
rect 19200 2818 20000 2848
rect 17174 2758 20000 2818
rect 3170 2752 3486 2753
rect 0 2682 800 2712
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 19200 2728 20000 2758
rect 16514 2687 16830 2688
rect 1485 2682 1551 2685
rect 0 2680 1551 2682
rect 0 2624 1490 2680
rect 1546 2624 1551 2680
rect 0 2622 1551 2624
rect 0 2592 800 2622
rect 1485 2619 1551 2622
rect 15142 2620 15148 2684
rect 15212 2682 15218 2684
rect 16205 2682 16271 2685
rect 15212 2680 16271 2682
rect 15212 2624 16210 2680
rect 16266 2624 16271 2680
rect 15212 2622 16271 2624
rect 15212 2620 15218 2622
rect 16205 2619 16271 2622
rect 17033 2682 17099 2685
rect 17350 2682 17356 2684
rect 17033 2680 17356 2682
rect 17033 2624 17038 2680
rect 17094 2624 17356 2680
rect 17033 2622 17356 2624
rect 17033 2619 17099 2622
rect 17350 2620 17356 2622
rect 17420 2620 17426 2684
rect 15193 2546 15259 2549
rect 19200 2546 20000 2576
rect 15193 2544 20000 2546
rect 15193 2488 15198 2544
rect 15254 2488 20000 2544
rect 15193 2486 20000 2488
rect 15193 2483 15259 2486
rect 19200 2456 20000 2486
rect 0 2410 800 2440
rect 2589 2410 2655 2413
rect 0 2408 2655 2410
rect 0 2352 2594 2408
rect 2650 2352 2655 2408
rect 0 2350 2655 2352
rect 0 2320 800 2350
rect 2589 2347 2655 2350
rect 15009 2410 15075 2413
rect 15929 2410 15995 2413
rect 17861 2410 17927 2413
rect 15009 2408 17927 2410
rect 15009 2352 15014 2408
rect 15070 2352 15934 2408
rect 15990 2352 17866 2408
rect 17922 2352 17927 2408
rect 15009 2350 17927 2352
rect 15009 2347 15075 2350
rect 15929 2347 15995 2350
rect 17861 2347 17927 2350
rect 5394 2208 5710 2209
rect 0 2138 800 2168
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 14290 2143 14606 2144
rect 1853 2138 1919 2141
rect 0 2136 1919 2138
rect 0 2080 1858 2136
rect 1914 2080 1919 2136
rect 0 2078 1919 2080
rect 0 2048 800 2078
rect 1853 2075 1919 2078
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
rect 0 1594 800 1624
rect 1669 1594 1735 1597
rect 0 1592 1735 1594
rect 0 1536 1674 1592
rect 1730 1536 1735 1592
rect 0 1534 1735 1536
rect 0 1504 800 1534
rect 1669 1531 1735 1534
<< via3 >>
rect 9076 14860 9140 14924
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 15700 13908 15764 13972
rect 6316 13636 6380 13700
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 4108 13228 4172 13292
rect 16252 13092 16316 13156
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 12572 12276 12636 12340
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 13860 11732 13924 11796
rect 11100 11520 11164 11524
rect 11100 11464 11114 11520
rect 11114 11464 11164 11520
rect 11100 11460 11164 11464
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 13676 9964 13740 10028
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 2084 9556 2148 9620
rect 16988 9556 17052 9620
rect 12940 9284 13004 9348
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 10364 9148 10428 9212
rect 2268 8876 2332 8940
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 4108 8332 4172 8396
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 8156 8120 8220 8124
rect 8156 8064 8170 8120
rect 8170 8064 8220 8120
rect 8156 8060 8220 8064
rect 2820 7924 2884 7988
rect 15148 7924 15212 7988
rect 17356 7924 17420 7988
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 7236 7516 7300 7580
rect 7236 7108 7300 7172
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 12572 7244 12636 7308
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 8156 6564 8220 6628
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 2084 6292 2148 6356
rect 16252 6700 16316 6764
rect 13860 6624 13924 6628
rect 13860 6568 13874 6624
rect 13874 6568 13924 6624
rect 13860 6564 13924 6568
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 12572 6488 12636 6492
rect 12572 6432 12622 6488
rect 12622 6432 12636 6488
rect 12572 6428 12636 6432
rect 15700 6156 15764 6220
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 17356 5944 17420 5948
rect 17356 5888 17370 5944
rect 17370 5888 17420 5944
rect 17356 5884 17420 5888
rect 12572 5748 12636 5812
rect 15700 5808 15764 5812
rect 15700 5752 15714 5808
rect 15714 5752 15764 5808
rect 15700 5748 15764 5752
rect 16252 5748 16316 5812
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 17356 5340 17420 5404
rect 2820 5264 2884 5268
rect 2820 5208 2834 5264
rect 2834 5208 2884 5264
rect 2820 5204 2884 5208
rect 13676 5128 13740 5132
rect 13676 5072 13690 5128
rect 13690 5072 13740 5128
rect 13676 5068 13740 5072
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 17356 4796 17420 4860
rect 10364 4720 10428 4724
rect 10364 4664 10378 4720
rect 10378 4664 10428 4720
rect 10364 4660 10428 4664
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 15148 4252 15212 4316
rect 4292 3980 4356 4044
rect 2268 3572 2332 3636
rect 12940 3980 13004 4044
rect 16988 3980 17052 4044
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 9076 3572 9140 3636
rect 15700 3572 15764 3636
rect 16252 3572 16316 3636
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 11100 3436 11164 3500
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 6316 3028 6380 3092
rect 4108 2892 4172 2956
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 15148 2620 15212 2684
rect 17356 2620 17420 2684
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 9075 14924 9141 14925
rect 9075 14860 9076 14924
rect 9140 14860 9141 14924
rect 9075 14859 9141 14860
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 4107 13292 4173 13293
rect 4107 13228 4108 13292
rect 4172 13290 4173 13292
rect 4172 13230 4354 13290
rect 4172 13228 4173 13230
rect 4107 13227 4173 13228
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 2083 9620 2149 9621
rect 2083 9556 2084 9620
rect 2148 9556 2149 9620
rect 2083 9555 2149 9556
rect 2086 6357 2146 9555
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 2267 8940 2333 8941
rect 2267 8876 2268 8940
rect 2332 8876 2333 8940
rect 2267 8875 2333 8876
rect 2083 6356 2149 6357
rect 2083 6292 2084 6356
rect 2148 6292 2149 6356
rect 2083 6291 2149 6292
rect 2270 3637 2330 8875
rect 3168 8192 3488 9216
rect 4107 8396 4173 8397
rect 4107 8332 4108 8396
rect 4172 8332 4173 8396
rect 4107 8331 4173 8332
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 2819 7988 2885 7989
rect 2819 7924 2820 7988
rect 2884 7924 2885 7988
rect 2819 7923 2885 7924
rect 2822 5269 2882 7923
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 2819 5268 2885 5269
rect 2819 5204 2820 5268
rect 2884 5204 2885 5268
rect 2819 5203 2885 5204
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 3840 3488 4864
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 2267 3636 2333 3637
rect 2267 3572 2268 3636
rect 2332 3572 2333 3636
rect 2267 3571 2333 3572
rect 3168 2752 3488 3776
rect 4110 2957 4170 8331
rect 4294 4045 4354 13230
rect 5392 13088 5712 14112
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 6315 13700 6381 13701
rect 6315 13636 6316 13700
rect 6380 13636 6381 13700
rect 6315 13635 6381 13636
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 4291 4044 4357 4045
rect 4291 3980 4292 4044
rect 4356 3980 4357 4044
rect 4291 3979 4357 3980
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 4107 2956 4173 2957
rect 4107 2892 4108 2956
rect 4172 2892 4173 2956
rect 4107 2891 4173 2892
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 2208 5712 3232
rect 6318 3093 6378 13635
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7235 7580 7301 7581
rect 7235 7516 7236 7580
rect 7300 7516 7301 7580
rect 7235 7515 7301 7516
rect 7238 7173 7298 7515
rect 7235 7172 7301 7173
rect 7235 7108 7236 7172
rect 7300 7108 7301 7172
rect 7235 7107 7301 7108
rect 7616 7104 7936 8128
rect 8155 8124 8221 8125
rect 8155 8060 8156 8124
rect 8220 8060 8221 8124
rect 8155 8059 8221 8060
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 8158 6629 8218 8059
rect 8155 6628 8221 6629
rect 8155 6564 8156 6628
rect 8220 6564 8221 6628
rect 8155 6563 8221 6564
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 6315 3092 6381 3093
rect 6315 3028 6316 3092
rect 6380 3028 6381 3092
rect 6315 3027 6381 3028
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2752 7936 3776
rect 9078 3637 9138 14859
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 11099 11524 11165 11525
rect 11099 11460 11100 11524
rect 11164 11460 11165 11524
rect 11099 11459 11165 11460
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 10363 9212 10429 9213
rect 10363 9148 10364 9212
rect 10428 9148 10429 9212
rect 10363 9147 10429 9148
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 10366 4725 10426 9147
rect 10363 4724 10429 4725
rect 10363 4660 10364 4724
rect 10428 4660 10429 4724
rect 10363 4659 10429 4660
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9075 3636 9141 3637
rect 9075 3572 9076 3636
rect 9140 3572 9141 3636
rect 9075 3571 9141 3572
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 9840 3296 10160 4320
rect 11102 3501 11162 11459
rect 12064 11456 12384 12480
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 15699 13972 15765 13973
rect 15699 13908 15700 13972
rect 15764 13908 15765 13972
rect 15699 13907 15765 13908
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 12571 12340 12637 12341
rect 12571 12276 12572 12340
rect 12636 12276 12637 12340
rect 12571 12275 12637 12276
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12574 7309 12634 12275
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 13859 11796 13925 11797
rect 13859 11732 13860 11796
rect 13924 11732 13925 11796
rect 13859 11731 13925 11732
rect 13675 10028 13741 10029
rect 13675 9964 13676 10028
rect 13740 9964 13741 10028
rect 13675 9963 13741 9964
rect 12939 9348 13005 9349
rect 12939 9284 12940 9348
rect 13004 9284 13005 9348
rect 12939 9283 13005 9284
rect 12571 7308 12637 7309
rect 12571 7244 12572 7308
rect 12636 7244 12637 7308
rect 12571 7243 12637 7244
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12571 6492 12637 6493
rect 12571 6428 12572 6492
rect 12636 6428 12637 6492
rect 12571 6427 12637 6428
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12574 5813 12634 6427
rect 12571 5812 12637 5813
rect 12571 5748 12572 5812
rect 12636 5748 12637 5812
rect 12571 5747 12637 5748
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12942 4045 13002 9283
rect 13678 5133 13738 9963
rect 13862 6629 13922 11731
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 15147 7988 15213 7989
rect 15147 7924 15148 7988
rect 15212 7924 15213 7988
rect 15147 7923 15213 7924
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 13859 6628 13925 6629
rect 13859 6564 13860 6628
rect 13924 6564 13925 6628
rect 13859 6563 13925 6564
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 13675 5132 13741 5133
rect 13675 5068 13676 5132
rect 13740 5068 13741 5132
rect 13675 5067 13741 5068
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 12939 4044 13005 4045
rect 12939 3980 12940 4044
rect 13004 3980 13005 4044
rect 12939 3979 13005 3980
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 11099 3500 11165 3501
rect 11099 3436 11100 3500
rect 11164 3436 11165 3500
rect 11099 3435 11165 3436
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 3296 14608 4320
rect 15150 4317 15210 7923
rect 15702 6221 15762 13907
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16251 13156 16317 13157
rect 16251 13092 16252 13156
rect 16316 13092 16317 13156
rect 16251 13091 16317 13092
rect 16254 6765 16314 13091
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16987 9620 17053 9621
rect 16987 9556 16988 9620
rect 17052 9556 17053 9620
rect 16987 9555 17053 9556
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16251 6764 16317 6765
rect 16251 6700 16252 6764
rect 16316 6700 16317 6764
rect 16251 6699 16317 6700
rect 15699 6220 15765 6221
rect 15699 6156 15700 6220
rect 15764 6156 15765 6220
rect 15699 6155 15765 6156
rect 15702 5813 15762 6155
rect 16254 5813 16314 6699
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 15699 5812 15765 5813
rect 15699 5748 15700 5812
rect 15764 5748 15765 5812
rect 15699 5747 15765 5748
rect 16251 5812 16317 5813
rect 16251 5748 16252 5812
rect 16316 5748 16317 5812
rect 16251 5747 16317 5748
rect 15147 4316 15213 4317
rect 15147 4252 15148 4316
rect 15212 4252 15213 4316
rect 15147 4251 15213 4252
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 15150 2685 15210 4251
rect 15702 3637 15762 5747
rect 16254 3637 16314 5747
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 3840 16832 4864
rect 16990 4045 17050 9555
rect 17355 7988 17421 7989
rect 17355 7924 17356 7988
rect 17420 7924 17421 7988
rect 17355 7923 17421 7924
rect 17358 5949 17418 7923
rect 17355 5948 17421 5949
rect 17355 5884 17356 5948
rect 17420 5884 17421 5948
rect 17355 5883 17421 5884
rect 17358 5405 17418 5883
rect 17355 5404 17421 5405
rect 17355 5340 17356 5404
rect 17420 5340 17421 5404
rect 17355 5339 17421 5340
rect 17358 4861 17418 5339
rect 17355 4860 17421 4861
rect 17355 4796 17356 4860
rect 17420 4796 17421 4860
rect 17355 4795 17421 4796
rect 16987 4044 17053 4045
rect 16987 3980 16988 4044
rect 17052 3980 17053 4044
rect 16987 3979 17053 3980
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 15699 3636 15765 3637
rect 15699 3572 15700 3636
rect 15764 3572 15765 3636
rect 15699 3571 15765 3572
rect 16251 3636 16317 3637
rect 16251 3572 16252 3636
rect 16316 3572 16317 3636
rect 16251 3571 16317 3572
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 15147 2684 15213 2685
rect 15147 2620 15148 2684
rect 15212 2620 15213 2684
rect 15147 2619 15213 2620
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2128 16832 2688
rect 17358 2685 17418 4795
rect 17355 2684 17421 2685
rect 17355 2620 17356 2684
rect 17420 2620 17421 2684
rect 17355 2619 17421 2620
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform -1 0 2944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1649977179
transform -1 0 13892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 1564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 15824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform -1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 15272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform -1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 17112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 17664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_N_FTB01_A
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_S_FTB01_A
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_E_FTB01_A
timestamp 1649977179
transform -1 0 17296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 2024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_E_FTB01_A
timestamp 1649977179
transform -1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_W_FTB01_A
timestamp 1649977179
transform 1 0 1472 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 18308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1649977179
transform -1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6624 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 4140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 17112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 17112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 16468 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 16192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 18584 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_N_FTB01_A
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_S_FTB01_A
timestamp 1649977179
transform -1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 1472 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1649977179
transform 1 0 1472 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_186
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1649977179
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1649977179
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_88
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_171
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_35
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_47
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_59
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1649977179
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_87
timestamp 1649977179
transform 1 0 9108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_113
timestamp 1649977179
transform 1 0 11500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_164
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_59
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1649977179
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_48
timestamp 1649977179
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_115
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_41
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_147
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_31
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_109
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_18
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_40
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_90
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_91
timestamp 1649977179
transform 1 0 9476 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_45
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_98
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_18
timestamp 1649977179
transform 1 0 2760 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_40
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_52
timestamp 1649977179
transform 1 0 5888 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_64
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1649977179
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_31
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_38
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_187
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_12
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1649977179
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1649977179
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_185
timestamp 1649977179
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _16_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1649977179
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform -1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform -1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform 1 0 3680 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _32_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1649977179
transform -1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform -1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 2760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform -1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform 1 0 16744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_1_S_FTB01
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1649977179
transform -1 0 2760 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1649977179
transform -1 0 2208 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13432 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8648 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13156 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11408 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9568 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11868 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9384 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14444 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14444 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15456 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16192 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16468 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14168 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14444 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15916 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2392 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2300 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1840 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9016 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2944 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2760 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3588 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5980 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6348 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7912 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9476 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4692 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3588 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4876 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7084 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6992 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16284 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9844 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10028 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 15824 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17940 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10948 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11316 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12052 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10672 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_N_FTB01
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_S_FTB01
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1649977179
transform -1 0 2208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1649977179
transform -1 0 2760 0 1 13056
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 REGIN_FEEDTHROUGH
port 0 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 REGOUT_FEEDTHROUGH
port 1 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 2 nsew signal input
flabel metal2 s 2042 16400 2098 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 3 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 4 nsew signal tristate
flabel metal2 s 5998 16400 6054 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 5 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 8 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 9 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 bottom_grid_pin_11_
port 10 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 11 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 bottom_grid_pin_13_
port 12 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 13 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 bottom_grid_pin_15_
port 14 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_1_
port 15 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 16 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 bottom_grid_pin_3_
port 17 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 18 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 bottom_grid_pin_5_
port 19 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 20 nsew signal tristate
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_pin_7_
port 21 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 22 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 bottom_grid_pin_9_
port 23 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 ccff_head
port 24 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 ccff_tail
port 25 nsew signal tristate
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 26 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 27 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 28 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 29 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 30 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 31 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 32 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 33 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 34 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 35 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 36 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 37 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 38 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 39 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 40 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 41 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 42 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 43 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 44 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 45 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 46 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 47 nsew signal tristate
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 48 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 49 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 50 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 51 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 52 nsew signal tristate
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 53 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 54 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 55 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 56 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 57 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 19200 9256 20000 9376 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 66 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 67 nsew signal input
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 68 nsew signal input
flabel metal3 s 19200 12520 20000 12640 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 69 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 70 nsew signal input
flabel metal3 s 19200 13064 20000 13184 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 71 nsew signal input
flabel metal3 s 19200 13336 20000 13456 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 72 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 73 nsew signal input
flabel metal3 s 19200 13880 20000 14000 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 74 nsew signal input
flabel metal3 s 19200 14152 20000 14272 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 75 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 76 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 77 nsew signal input
flabel metal3 s 19200 9800 20000 9920 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 78 nsew signal input
flabel metal3 s 19200 10072 20000 10192 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 79 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 80 nsew signal input
flabel metal3 s 19200 10616 20000 10736 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 81 nsew signal input
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 82 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 83 nsew signal input
flabel metal3 s 19200 11432 20000 11552 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 84 nsew signal input
flabel metal3 s 19200 11704 20000 11824 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 85 nsew signal input
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 86 nsew signal tristate
flabel metal3 s 19200 6536 20000 6656 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 87 nsew signal tristate
flabel metal3 s 19200 6808 20000 6928 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 88 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 89 nsew signal tristate
flabel metal3 s 19200 7352 20000 7472 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 90 nsew signal tristate
flabel metal3 s 19200 7624 20000 7744 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 91 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 92 nsew signal tristate
flabel metal3 s 19200 8168 20000 8288 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 93 nsew signal tristate
flabel metal3 s 19200 8440 20000 8560 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 94 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 95 nsew signal tristate
flabel metal3 s 19200 8984 20000 9104 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 96 nsew signal tristate
flabel metal3 s 19200 4088 20000 4208 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 97 nsew signal tristate
flabel metal3 s 19200 4360 20000 4480 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 98 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 99 nsew signal tristate
flabel metal3 s 19200 4904 20000 5024 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 100 nsew signal tristate
flabel metal3 s 19200 5176 20000 5296 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 101 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 102 nsew signal tristate
flabel metal3 s 19200 5720 20000 5840 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 103 nsew signal tristate
flabel metal3 s 19200 5992 20000 6112 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 104 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 105 nsew signal tristate
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 clk_1_N_out
port 106 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 clk_1_S_out
port 107 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 clk_1_W_in
port 108 nsew signal input
flabel metal3 s 19200 3544 20000 3664 0 FreeSans 480 0 0 0 clk_2_E_out
port 109 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 clk_2_W_in
port 110 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 clk_2_W_out
port 111 nsew signal tristate
flabel metal3 s 19200 3272 20000 3392 0 FreeSans 480 0 0 0 clk_3_E_out
port 112 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 clk_3_W_in
port 113 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 clk_3_W_out
port 114 nsew signal tristate
flabel metal2 s 13910 16400 13966 17200 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 115 nsew signal input
flabel metal2 s 17866 16400 17922 17200 0 FreeSans 224 90 0 0 prog_clk_0_W_out
port 116 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 prog_clk_1_N_out
port 117 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 prog_clk_1_S_out
port 118 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 prog_clk_1_W_in
port 119 nsew signal input
flabel metal3 s 19200 2728 20000 2848 0 FreeSans 480 0 0 0 prog_clk_2_E_out
port 120 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 prog_clk_2_W_in
port 121 nsew signal input
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 prog_clk_2_W_out
port 122 nsew signal tristate
flabel metal3 s 19200 2456 20000 2576 0 FreeSans 480 0 0 0 prog_clk_3_E_out
port 123 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 prog_clk_3_W_in
port 124 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 prog_clk_3_W_out
port 125 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
