magic
tech sky130A
magscale 1 2
timestamp 1656945783
<< viali >>
rect 2881 20553 2915 20587
rect 3341 20553 3375 20587
rect 4445 20553 4479 20587
rect 4813 20553 4847 20587
rect 6377 20553 6411 20587
rect 6653 20553 6687 20587
rect 7389 20553 7423 20587
rect 7849 20553 7883 20587
rect 9229 20553 9263 20587
rect 9689 20553 9723 20587
rect 10149 20553 10183 20587
rect 10609 20553 10643 20587
rect 15761 20553 15795 20587
rect 16313 20553 16347 20587
rect 16865 20553 16899 20587
rect 2973 20485 3007 20519
rect 3249 20485 3283 20519
rect 7481 20485 7515 20519
rect 8217 20485 8251 20519
rect 11069 20485 11103 20519
rect 11805 20485 11839 20519
rect 14473 20485 14507 20519
rect 3525 20417 3559 20451
rect 3985 20417 4019 20451
rect 4997 20417 5031 20451
rect 6193 20417 6227 20451
rect 8309 20417 8343 20451
rect 9321 20417 9355 20451
rect 10977 20417 11011 20451
rect 11897 20417 11931 20451
rect 12357 20417 12391 20451
rect 15577 20417 15611 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 4169 20349 4203 20383
rect 4353 20349 4387 20383
rect 5273 20349 5307 20383
rect 7205 20349 7239 20383
rect 8033 20349 8067 20383
rect 9045 20349 9079 20383
rect 9873 20349 9907 20383
rect 10057 20349 10091 20383
rect 11253 20349 11287 20383
rect 11529 20349 11563 20383
rect 13829 20349 13863 20383
rect 14565 20349 14599 20383
rect 14749 20349 14783 20383
rect 6837 20281 6871 20315
rect 10517 20281 10551 20315
rect 13461 20281 13495 20315
rect 13645 20281 13679 20315
rect 6929 20213 6963 20247
rect 8677 20213 8711 20247
rect 12081 20213 12115 20247
rect 13001 20213 13035 20247
rect 13277 20213 13311 20247
rect 14105 20213 14139 20247
rect 16037 20213 16071 20247
rect 17969 20213 18003 20247
rect 20729 20213 20763 20247
rect 21097 20213 21131 20247
rect 1961 20009 1995 20043
rect 2329 20009 2363 20043
rect 2881 20009 2915 20043
rect 7205 20009 7239 20043
rect 11437 20009 11471 20043
rect 13829 20009 13863 20043
rect 14105 20009 14139 20043
rect 15485 20009 15519 20043
rect 15761 20009 15795 20043
rect 17785 20009 17819 20043
rect 18245 20009 18279 20043
rect 19809 20009 19843 20043
rect 20177 20009 20211 20043
rect 20545 20009 20579 20043
rect 21373 20009 21407 20043
rect 11069 19941 11103 19975
rect 11253 19941 11287 19975
rect 15117 19941 15151 19975
rect 18981 19941 19015 19975
rect 21005 19941 21039 19975
rect 7757 19873 7791 19907
rect 8217 19873 8251 19907
rect 11897 19873 11931 19907
rect 11989 19873 12023 19907
rect 13277 19873 13311 19907
rect 13369 19873 13403 19907
rect 14749 19873 14783 19907
rect 15945 19873 15979 19907
rect 2145 19805 2179 19839
rect 2513 19805 2547 19839
rect 3433 19805 3467 19839
rect 3893 19805 3927 19839
rect 6745 19805 6779 19839
rect 8309 19805 8343 19839
rect 8401 19805 8435 19839
rect 9597 19805 9631 19839
rect 11805 19805 11839 19839
rect 12541 19805 12575 19839
rect 14933 19805 14967 19839
rect 15301 19805 15335 19839
rect 16221 19805 16255 19839
rect 16773 19805 16807 19839
rect 16865 19805 16899 19839
rect 17141 19805 17175 19839
rect 17601 19805 17635 19839
rect 18061 19805 18095 19839
rect 18429 19805 18463 19839
rect 18797 19805 18831 19839
rect 19625 19805 19659 19839
rect 20361 19805 20395 19839
rect 20821 19805 20855 19839
rect 21189 19805 21223 19839
rect 3617 19737 3651 19771
rect 4160 19737 4194 19771
rect 6500 19737 6534 19771
rect 9045 19737 9079 19771
rect 9413 19737 9447 19771
rect 9842 19737 9876 19771
rect 13461 19737 13495 19771
rect 14473 19737 14507 19771
rect 16129 19737 16163 19771
rect 17417 19737 17451 19771
rect 2697 19669 2731 19703
rect 5273 19669 5307 19703
rect 5365 19669 5399 19703
rect 6929 19669 6963 19703
rect 7113 19669 7147 19703
rect 7573 19669 7607 19703
rect 7665 19669 7699 19703
rect 8769 19669 8803 19703
rect 9229 19669 9263 19703
rect 10977 19669 11011 19703
rect 12449 19669 12483 19703
rect 12725 19669 12759 19703
rect 14565 19669 14599 19703
rect 16589 19669 16623 19703
rect 18613 19669 18647 19703
rect 19533 19669 19567 19703
rect 3617 19465 3651 19499
rect 4077 19465 4111 19499
rect 4445 19465 4479 19499
rect 4629 19465 4663 19499
rect 6193 19465 6227 19499
rect 6745 19465 6779 19499
rect 9597 19465 9631 19499
rect 13645 19465 13679 19499
rect 14749 19465 14783 19499
rect 14933 19465 14967 19499
rect 16129 19465 16163 19499
rect 16405 19465 16439 19499
rect 16681 19465 16715 19499
rect 17049 19465 17083 19499
rect 17509 19465 17543 19499
rect 18889 19465 18923 19499
rect 21005 19465 21039 19499
rect 3525 19397 3559 19431
rect 9956 19397 9990 19431
rect 17141 19397 17175 19431
rect 17877 19397 17911 19431
rect 3985 19329 4019 19363
rect 4813 19329 4847 19363
rect 5080 19329 5114 19363
rect 7869 19329 7903 19363
rect 8125 19329 8159 19363
rect 8217 19329 8251 19363
rect 8484 19329 8518 19363
rect 9689 19329 9723 19363
rect 12653 19329 12687 19363
rect 13461 19329 13495 19363
rect 14289 19329 14323 19363
rect 14381 19329 14415 19363
rect 15117 19329 15151 19363
rect 15577 19329 15611 19363
rect 16313 19329 16347 19363
rect 18337 19329 18371 19363
rect 18705 19329 18739 19363
rect 20821 19329 20855 19363
rect 4169 19261 4203 19295
rect 12909 19261 12943 19295
rect 13001 19261 13035 19295
rect 13277 19261 13311 19295
rect 14105 19261 14139 19295
rect 15669 19261 15703 19295
rect 15761 19261 15795 19295
rect 17233 19261 17267 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 11253 19193 11287 19227
rect 18521 19193 18555 19227
rect 6377 19125 6411 19159
rect 6561 19125 6595 19159
rect 11069 19125 11103 19159
rect 11529 19125 11563 19159
rect 13829 19125 13863 19159
rect 15209 19125 15243 19159
rect 20729 19125 20763 19159
rect 4445 18921 4479 18955
rect 4629 18921 4663 18955
rect 7297 18921 7331 18955
rect 10977 18921 11011 18955
rect 13829 18921 13863 18955
rect 17049 18921 17083 18955
rect 21005 18921 21039 18955
rect 7389 18853 7423 18887
rect 9045 18853 9079 18887
rect 11069 18853 11103 18887
rect 15853 18853 15887 18887
rect 4721 18785 4755 18819
rect 6745 18785 6779 18819
rect 12449 18785 12483 18819
rect 13185 18785 13219 18819
rect 15209 18785 15243 18819
rect 16589 18785 16623 18819
rect 17969 18785 18003 18819
rect 18429 18785 18463 18819
rect 6193 18717 6227 18751
rect 6377 18717 6411 18751
rect 6837 18717 6871 18751
rect 8769 18717 8803 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 12182 18717 12216 18751
rect 15485 18717 15519 18751
rect 16865 18717 16899 18751
rect 17233 18717 17267 18751
rect 18245 18717 18279 18751
rect 20821 18717 20855 18751
rect 4077 18649 4111 18683
rect 4988 18649 5022 18683
rect 8524 18649 8558 18683
rect 9864 18649 9898 18683
rect 13001 18649 13035 18683
rect 13553 18649 13587 18683
rect 15393 18649 15427 18683
rect 16405 18649 16439 18683
rect 17509 18649 17543 18683
rect 4261 18581 4295 18615
rect 6101 18581 6135 18615
rect 6929 18581 6963 18615
rect 9137 18581 9171 18615
rect 12633 18581 12667 18615
rect 13093 18581 13127 18615
rect 13645 18581 13679 18615
rect 16037 18581 16071 18615
rect 16497 18581 16531 18615
rect 20729 18581 20763 18615
rect 1961 18377 1995 18411
rect 6009 18377 6043 18411
rect 6193 18377 6227 18411
rect 12541 18377 12575 18411
rect 14289 18377 14323 18411
rect 14749 18377 14783 18411
rect 15577 18377 15611 18411
rect 16865 18377 16899 18411
rect 21005 18377 21039 18411
rect 5558 18309 5592 18343
rect 9413 18309 9447 18343
rect 9781 18309 9815 18343
rect 13645 18309 13679 18343
rect 15117 18309 15151 18343
rect 17417 18309 17451 18343
rect 2145 18241 2179 18275
rect 5825 18241 5859 18275
rect 6377 18241 6411 18275
rect 6644 18241 6678 18275
rect 7941 18241 7975 18275
rect 8208 18241 8242 18275
rect 11089 18241 11123 18275
rect 11345 18241 11379 18275
rect 13921 18241 13955 18275
rect 14381 18241 14415 18275
rect 14841 18241 14875 18275
rect 17141 18241 17175 18275
rect 20821 18241 20855 18275
rect 14105 18173 14139 18207
rect 15853 18173 15887 18207
rect 17693 18173 17727 18207
rect 2329 18105 2363 18139
rect 9321 18105 9355 18139
rect 2421 18037 2455 18071
rect 4445 18037 4479 18071
rect 7757 18037 7791 18071
rect 9965 18037 9999 18071
rect 13277 18037 13311 18071
rect 19165 18037 19199 18071
rect 1961 17833 1995 17867
rect 3341 17833 3375 17867
rect 5917 17833 5951 17867
rect 13921 17833 13955 17867
rect 14933 17833 14967 17867
rect 16037 17833 16071 17867
rect 17233 17833 17267 17867
rect 18245 17833 18279 17867
rect 20269 17833 20303 17867
rect 5825 17765 5859 17799
rect 2421 17697 2455 17731
rect 4445 17697 4479 17731
rect 7297 17697 7331 17731
rect 7389 17697 7423 17731
rect 13369 17697 13403 17731
rect 13553 17697 13587 17731
rect 14657 17697 14691 17731
rect 15393 17697 15427 17731
rect 15485 17697 15519 17731
rect 16221 17697 16255 17731
rect 16497 17697 16531 17731
rect 17785 17697 17819 17731
rect 18797 17697 18831 17731
rect 19809 17697 19843 17731
rect 2145 17629 2179 17663
rect 2605 17629 2639 17663
rect 4712 17629 4746 17663
rect 8953 17629 8987 17663
rect 9873 17629 9907 17663
rect 10057 17629 10091 17663
rect 10324 17629 10358 17663
rect 16681 17629 16715 17663
rect 20085 17629 20119 17663
rect 3065 17561 3099 17595
rect 7030 17561 7064 17595
rect 7656 17561 7690 17595
rect 16773 17561 16807 17595
rect 18613 17561 18647 17595
rect 2513 17493 2547 17527
rect 2973 17493 3007 17527
rect 8769 17493 8803 17527
rect 11437 17493 11471 17527
rect 12909 17493 12943 17527
rect 13277 17493 13311 17527
rect 14105 17493 14139 17527
rect 14473 17493 14507 17527
rect 14565 17493 14599 17527
rect 15301 17493 15335 17527
rect 17141 17493 17175 17527
rect 17601 17493 17635 17527
rect 17693 17493 17727 17527
rect 18705 17493 18739 17527
rect 19257 17493 19291 17527
rect 19625 17493 19659 17527
rect 19717 17493 19751 17527
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 2697 17289 2731 17323
rect 3065 17289 3099 17323
rect 6469 17289 6503 17323
rect 6653 17289 6687 17323
rect 6837 17289 6871 17323
rect 7205 17289 7239 17323
rect 9781 17289 9815 17323
rect 12817 17289 12851 17323
rect 14013 17289 14047 17323
rect 17325 17289 17359 17323
rect 17693 17289 17727 17323
rect 18337 17289 18371 17323
rect 19165 17289 19199 17323
rect 19993 17289 20027 17323
rect 21005 17289 21039 17323
rect 21373 17289 21407 17323
rect 3249 17221 3283 17255
rect 13001 17221 13035 17255
rect 14749 17221 14783 17255
rect 16221 17221 16255 17255
rect 17969 17221 18003 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 5926 17153 5960 17187
rect 6193 17153 6227 17187
rect 7297 17153 7331 17187
rect 7564 17153 7598 17187
rect 9965 17153 9999 17187
rect 10232 17153 10266 17187
rect 13093 17153 13127 17187
rect 13921 17153 13955 17187
rect 14473 17153 14507 17187
rect 16497 17153 16531 17187
rect 16865 17153 16899 17187
rect 18245 17153 18279 17187
rect 18705 17153 18739 17187
rect 19533 17153 19567 17187
rect 20729 17153 20763 17187
rect 20821 17153 20855 17187
rect 21189 17153 21223 17187
rect 13277 17085 13311 17119
rect 13737 17085 13771 17119
rect 17049 17085 17083 17119
rect 17233 17085 17267 17119
rect 18797 17085 18831 17119
rect 18889 17085 18923 17119
rect 19625 17085 19659 17119
rect 19809 17085 19843 17119
rect 11345 17017 11379 17051
rect 4813 16949 4847 16983
rect 8677 16949 8711 16983
rect 12173 16949 12207 16983
rect 14381 16949 14415 16983
rect 20269 16949 20303 16983
rect 6285 16745 6319 16779
rect 6377 16745 6411 16779
rect 6561 16745 6595 16779
rect 7021 16745 7055 16779
rect 16313 16745 16347 16779
rect 18153 16745 18187 16779
rect 19257 16745 19291 16779
rect 18981 16677 19015 16711
rect 2881 16609 2915 16643
rect 4353 16609 4387 16643
rect 4721 16609 4755 16643
rect 8585 16609 8619 16643
rect 16773 16609 16807 16643
rect 16957 16609 16991 16643
rect 1777 16541 1811 16575
rect 2145 16541 2179 16575
rect 2789 16541 2823 16575
rect 12265 16541 12299 16575
rect 12357 16541 12391 16575
rect 14749 16541 14783 16575
rect 15025 16541 15059 16575
rect 15577 16541 15611 16575
rect 15853 16541 15887 16575
rect 17141 16541 17175 16575
rect 2697 16473 2731 16507
rect 4261 16473 4295 16507
rect 4988 16473 5022 16507
rect 8318 16473 8352 16507
rect 12020 16473 12054 16507
rect 12624 16473 12658 16507
rect 17417 16473 17451 16507
rect 1961 16405 1995 16439
rect 2329 16405 2363 16439
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 6101 16405 6135 16439
rect 7205 16405 7239 16439
rect 10701 16405 10735 16439
rect 10885 16405 10919 16439
rect 13737 16405 13771 16439
rect 16681 16405 16715 16439
rect 2605 16201 2639 16235
rect 6377 16201 6411 16235
rect 9781 16201 9815 16235
rect 14473 16201 14507 16235
rect 14841 16201 14875 16235
rect 15669 16201 15703 16235
rect 16037 16201 16071 16235
rect 16497 16201 16531 16235
rect 17785 16201 17819 16235
rect 17969 16201 18003 16235
rect 18429 16133 18463 16167
rect 20729 16133 20763 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2513 16065 2547 16099
rect 3341 16065 3375 16099
rect 4077 16065 4111 16099
rect 5742 16065 5776 16099
rect 6009 16065 6043 16099
rect 7490 16065 7524 16099
rect 7757 16065 7791 16099
rect 7941 16065 7975 16099
rect 8208 16065 8242 16099
rect 9965 16065 9999 16099
rect 10232 16065 10266 16099
rect 12642 16065 12676 16099
rect 12909 16065 12943 16099
rect 16129 16065 16163 16099
rect 17049 16065 17083 16099
rect 18337 16065 18371 16099
rect 18797 16065 18831 16099
rect 20453 16065 20487 16099
rect 2789 15997 2823 16031
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 9505 15997 9539 16031
rect 14933 15997 14967 16031
rect 15025 15997 15059 16031
rect 15945 15997 15979 16031
rect 17141 15997 17175 16031
rect 17325 15997 17359 16031
rect 18521 15997 18555 16031
rect 1869 15929 1903 15963
rect 4261 15929 4295 15963
rect 11345 15929 11379 15963
rect 2145 15861 2179 15895
rect 3709 15861 3743 15895
rect 3893 15861 3927 15895
rect 4629 15861 4663 15895
rect 6193 15861 6227 15895
rect 9321 15861 9355 15895
rect 11529 15861 11563 15895
rect 16681 15861 16715 15895
rect 3985 15657 4019 15691
rect 7021 15657 7055 15691
rect 7205 15657 7239 15691
rect 10425 15657 10459 15691
rect 12081 15657 12115 15691
rect 14289 15657 14323 15691
rect 15301 15657 15335 15691
rect 17233 15657 17267 15691
rect 17417 15657 17451 15691
rect 5549 15589 5583 15623
rect 10333 15589 10367 15623
rect 19993 15589 20027 15623
rect 5457 15521 5491 15555
rect 6929 15521 6963 15555
rect 8769 15521 8803 15555
rect 8953 15521 8987 15555
rect 10609 15521 10643 15555
rect 14105 15521 14139 15555
rect 14565 15521 14599 15555
rect 15853 15521 15887 15555
rect 16497 15521 16531 15555
rect 17969 15521 18003 15555
rect 19349 15521 19383 15555
rect 20545 15521 20579 15555
rect 1961 15453 1995 15487
rect 5201 15453 5235 15487
rect 9220 15453 9254 15487
rect 16405 15453 16439 15487
rect 17877 15453 17911 15487
rect 18245 15453 18279 15487
rect 20269 15453 20303 15487
rect 2237 15385 2271 15419
rect 6684 15385 6718 15419
rect 8524 15385 8558 15419
rect 10854 15385 10888 15419
rect 13829 15385 13863 15419
rect 14749 15385 14783 15419
rect 14841 15385 14875 15419
rect 15669 15385 15703 15419
rect 15761 15385 15795 15419
rect 4077 15317 4111 15351
rect 7389 15317 7423 15351
rect 11989 15317 12023 15351
rect 15209 15317 15243 15351
rect 16865 15317 16899 15351
rect 17785 15317 17819 15351
rect 18521 15317 18555 15351
rect 19533 15317 19567 15351
rect 19625 15317 19659 15351
rect 1961 15113 1995 15147
rect 4445 15113 4479 15147
rect 6469 15113 6503 15147
rect 6653 15113 6687 15147
rect 7021 15113 7055 15147
rect 7665 15113 7699 15147
rect 9229 15113 9263 15147
rect 9413 15113 9447 15147
rect 13185 15113 13219 15147
rect 13461 15113 13495 15147
rect 14013 15113 14047 15147
rect 15761 15113 15795 15147
rect 17233 15113 17267 15147
rect 19165 15113 19199 15147
rect 19625 15113 19659 15147
rect 19717 15113 19751 15147
rect 21005 15113 21039 15147
rect 21373 15113 21407 15147
rect 3801 15045 3835 15079
rect 3893 15045 3927 15079
rect 4629 15045 4663 15079
rect 17601 15045 17635 15079
rect 18429 15045 18463 15079
rect 20177 15045 20211 15079
rect 20637 15045 20671 15079
rect 2145 14977 2179 15011
rect 4813 14977 4847 15011
rect 5069 14977 5103 15011
rect 7849 14977 7883 15011
rect 8116 14977 8150 15011
rect 12653 14977 12687 15011
rect 12909 14977 12943 15011
rect 13921 14977 13955 15011
rect 15209 14977 15243 15011
rect 16129 14977 16163 15011
rect 16681 14977 16715 15011
rect 19257 14977 19291 15011
rect 20085 14977 20119 15011
rect 20821 14977 20855 15011
rect 21189 14977 21223 15011
rect 3709 14909 3743 14943
rect 14105 14909 14139 14943
rect 14473 14909 14507 14943
rect 15301 14909 15335 14943
rect 15393 14909 15427 14943
rect 16221 14909 16255 14943
rect 16405 14909 16439 14943
rect 17141 14909 17175 14943
rect 17693 14909 17727 14943
rect 17785 14909 17819 14943
rect 18153 14909 18187 14943
rect 18337 14909 18371 14943
rect 18981 14909 19015 14943
rect 20269 14909 20303 14943
rect 4261 14841 4295 14875
rect 11529 14841 11563 14875
rect 13553 14841 13587 14875
rect 14565 14841 14599 14875
rect 6193 14773 6227 14807
rect 7297 14773 7331 14807
rect 11253 14773 11287 14807
rect 14841 14773 14875 14807
rect 18797 14773 18831 14807
rect 5641 14569 5675 14603
rect 7205 14569 7239 14603
rect 11161 14569 11195 14603
rect 17785 14569 17819 14603
rect 21005 14569 21039 14603
rect 13645 14501 13679 14535
rect 14105 14501 14139 14535
rect 3341 14433 3375 14467
rect 3525 14433 3559 14467
rect 4261 14433 4295 14467
rect 5733 14433 5767 14467
rect 8769 14433 8803 14467
rect 14565 14433 14599 14467
rect 14657 14433 14691 14467
rect 14933 14433 14967 14467
rect 17141 14433 17175 14467
rect 17325 14433 17359 14467
rect 18521 14433 18555 14467
rect 19625 14433 19659 14467
rect 12725 14365 12759 14399
rect 18705 14365 18739 14399
rect 19349 14365 19383 14399
rect 20821 14365 20855 14399
rect 4169 14297 4203 14331
rect 4528 14297 4562 14331
rect 5978 14297 6012 14331
rect 8524 14297 8558 14331
rect 12480 14297 12514 14331
rect 13829 14297 13863 14331
rect 17417 14297 17451 14331
rect 21189 14297 21223 14331
rect 2881 14229 2915 14263
rect 3249 14229 3283 14263
rect 3985 14229 4019 14263
rect 7113 14229 7147 14263
rect 7389 14229 7423 14263
rect 11345 14229 11379 14263
rect 14473 14229 14507 14263
rect 15577 14229 15611 14263
rect 17877 14229 17911 14263
rect 18245 14229 18279 14263
rect 18337 14229 18371 14263
rect 20729 14229 20763 14263
rect 1593 14025 1627 14059
rect 1961 14025 1995 14059
rect 3525 14025 3559 14059
rect 4537 14025 4571 14059
rect 6193 14025 6227 14059
rect 9413 14025 9447 14059
rect 9781 14025 9815 14059
rect 11345 14025 11379 14059
rect 17509 14025 17543 14059
rect 19349 14025 19383 14059
rect 20269 14025 20303 14059
rect 20637 14025 20671 14059
rect 21281 14025 21315 14059
rect 5661 13957 5695 13991
rect 17693 13957 17727 13991
rect 18061 13957 18095 13991
rect 1777 13889 1811 13923
rect 2145 13889 2179 13923
rect 2697 13889 2731 13923
rect 2973 13889 3007 13923
rect 3433 13889 3467 13923
rect 7490 13889 7524 13923
rect 7757 13889 7791 13923
rect 7849 13889 7883 13923
rect 8116 13889 8150 13923
rect 9965 13889 9999 13923
rect 10232 13889 10266 13923
rect 11529 13889 11563 13923
rect 11785 13889 11819 13923
rect 19165 13889 19199 13923
rect 20085 13889 20119 13923
rect 20729 13889 20763 13923
rect 21097 13889 21131 13923
rect 3709 13821 3743 13855
rect 5917 13821 5951 13855
rect 18981 13821 19015 13855
rect 19625 13821 19659 13855
rect 20821 13821 20855 13855
rect 21465 13821 21499 13855
rect 6377 13753 6411 13787
rect 9229 13753 9263 13787
rect 13001 13753 13035 13787
rect 3065 13685 3099 13719
rect 12909 13685 12943 13719
rect 8585 13481 8619 13515
rect 10977 13481 11011 13515
rect 15301 13481 15335 13515
rect 17233 13481 17267 13515
rect 18981 13481 19015 13515
rect 20085 13481 20119 13515
rect 6193 13413 6227 13447
rect 12541 13413 12575 13447
rect 18153 13413 18187 13447
rect 19257 13413 19291 13447
rect 8309 13345 8343 13379
rect 11161 13345 11195 13379
rect 15485 13345 15519 13379
rect 15669 13345 15703 13379
rect 16589 13345 16623 13379
rect 17509 13345 17543 13379
rect 18337 13345 18371 13379
rect 19809 13345 19843 13379
rect 20637 13345 20671 13379
rect 4813 13277 4847 13311
rect 8053 13277 8087 13311
rect 8493 13277 8527 13311
rect 11428 13277 11462 13311
rect 12633 13277 12667 13311
rect 16773 13277 16807 13311
rect 18613 13277 18647 13311
rect 5080 13209 5114 13243
rect 6285 13209 6319 13243
rect 6469 13209 6503 13243
rect 6745 13209 6779 13243
rect 18521 13209 18555 13243
rect 20453 13209 20487 13243
rect 6929 13141 6963 13175
rect 15761 13141 15795 13175
rect 16129 13141 16163 13175
rect 16313 13141 16347 13175
rect 16865 13141 16899 13175
rect 17693 13141 17727 13175
rect 17785 13141 17819 13175
rect 19625 13141 19659 13175
rect 19717 13141 19751 13175
rect 20545 13141 20579 13175
rect 8033 12937 8067 12971
rect 9597 12937 9631 12971
rect 9781 12937 9815 12971
rect 11345 12937 11379 12971
rect 13369 12937 13403 12971
rect 14013 12937 14047 12971
rect 14473 12937 14507 12971
rect 16957 12937 16991 12971
rect 17417 12937 17451 12971
rect 17509 12937 17543 12971
rect 18613 12937 18647 12971
rect 19441 12937 19475 12971
rect 20269 12937 20303 12971
rect 20637 12937 20671 12971
rect 21189 12937 21223 12971
rect 5304 12869 5338 12903
rect 10232 12869 10266 12903
rect 11796 12869 11830 12903
rect 13553 12869 13587 12903
rect 14105 12869 14139 12903
rect 17969 12869 18003 12903
rect 6828 12801 6862 12835
rect 9157 12801 9191 12835
rect 9413 12801 9447 12835
rect 9965 12801 9999 12835
rect 11529 12801 11563 12835
rect 15853 12801 15887 12835
rect 17049 12801 17083 12835
rect 17877 12801 17911 12835
rect 18337 12801 18371 12835
rect 18981 12801 19015 12835
rect 19809 12801 19843 12835
rect 5549 12733 5583 12767
rect 6561 12733 6595 12767
rect 13829 12733 13863 12767
rect 16129 12733 16163 12767
rect 16865 12733 16899 12767
rect 18061 12733 18095 12767
rect 19073 12733 19107 12767
rect 19257 12733 19291 12767
rect 19901 12733 19935 12767
rect 19993 12733 20027 12767
rect 20729 12733 20763 12767
rect 20821 12733 20855 12767
rect 7941 12665 7975 12699
rect 13001 12665 13035 12699
rect 4169 12597 4203 12631
rect 5641 12597 5675 12631
rect 6101 12597 6135 12631
rect 6377 12597 6411 12631
rect 12909 12597 12943 12631
rect 15025 12597 15059 12631
rect 21281 12597 21315 12631
rect 11161 12393 11195 12427
rect 14105 12393 14139 12427
rect 14933 12393 14967 12427
rect 17877 12393 17911 12427
rect 19533 12393 19567 12427
rect 20177 12393 20211 12427
rect 21189 12393 21223 12427
rect 5917 12325 5951 12359
rect 17969 12325 18003 12359
rect 12725 12257 12759 12291
rect 14657 12257 14691 12291
rect 15669 12257 15703 12291
rect 17233 12257 17267 12291
rect 17417 12257 17451 12291
rect 18521 12257 18555 12291
rect 19257 12257 19291 12291
rect 19809 12257 19843 12291
rect 20729 12257 20763 12291
rect 4169 12189 4203 12223
rect 5825 12189 5859 12223
rect 7297 12189 7331 12223
rect 7389 12189 7423 12223
rect 8953 12189 8987 12223
rect 17049 12189 17083 12223
rect 18429 12189 18463 12223
rect 21005 12189 21039 12223
rect 4414 12121 4448 12155
rect 7030 12121 7064 12155
rect 7634 12121 7668 12155
rect 9198 12121 9232 12155
rect 12480 12121 12514 12155
rect 15485 12121 15519 12155
rect 15945 12121 15979 12155
rect 20545 12121 20579 12155
rect 21373 12121 21407 12155
rect 1777 12053 1811 12087
rect 5549 12053 5583 12087
rect 8769 12053 8803 12087
rect 10333 12053 10367 12087
rect 11345 12053 11379 12087
rect 14473 12053 14507 12087
rect 14565 12053 14599 12087
rect 15117 12053 15151 12087
rect 15577 12053 15611 12087
rect 17509 12053 17543 12087
rect 18337 12053 18371 12087
rect 18797 12053 18831 12087
rect 20637 12053 20671 12087
rect 2329 11849 2363 11883
rect 2789 11849 2823 11883
rect 8677 11849 8711 11883
rect 11253 11849 11287 11883
rect 13553 11849 13587 11883
rect 14749 11849 14783 11883
rect 15025 11849 15059 11883
rect 15393 11849 15427 11883
rect 16681 11849 16715 11883
rect 16957 11849 16991 11883
rect 17417 11849 17451 11883
rect 17969 11849 18003 11883
rect 19717 11849 19751 11883
rect 20821 11849 20855 11883
rect 21097 11849 21131 11883
rect 1961 11781 1995 11815
rect 4620 11781 4654 11815
rect 5917 11781 5951 11815
rect 6101 11781 6135 11815
rect 6469 11781 6503 11815
rect 7297 11781 7331 11815
rect 7481 11781 7515 11815
rect 8401 11781 8435 11815
rect 8585 11781 8619 11815
rect 13001 11781 13035 11815
rect 14381 11781 14415 11815
rect 19901 11781 19935 11815
rect 20361 11781 20395 11815
rect 20453 11781 20487 11815
rect 21281 11781 21315 11815
rect 1685 11713 1719 11747
rect 2237 11713 2271 11747
rect 2697 11713 2731 11747
rect 8217 11713 8251 11747
rect 9801 11713 9835 11747
rect 10057 11713 10091 11747
rect 11529 11713 11563 11747
rect 11796 11713 11830 11747
rect 14289 11713 14323 11747
rect 16497 11713 16531 11747
rect 17325 11713 17359 11747
rect 18613 11713 18647 11747
rect 19625 11713 19659 11747
rect 20913 11713 20947 11747
rect 2973 11645 3007 11679
rect 4353 11645 4387 11679
rect 10241 11645 10275 11679
rect 13645 11645 13679 11679
rect 13737 11645 13771 11679
rect 14105 11645 14139 11679
rect 15485 11645 15519 11679
rect 15577 11645 15611 11679
rect 17509 11645 17543 11679
rect 18705 11645 18739 11679
rect 18889 11645 18923 11679
rect 20177 11645 20211 11679
rect 1501 11577 1535 11611
rect 18245 11577 18279 11611
rect 19165 11577 19199 11611
rect 5733 11509 5767 11543
rect 12909 11509 12943 11543
rect 13185 11509 13219 11543
rect 18061 11509 18095 11543
rect 2329 11305 2363 11339
rect 10701 11305 10735 11339
rect 10885 11305 10919 11339
rect 10977 11305 11011 11339
rect 17049 11305 17083 11339
rect 18981 11305 19015 11339
rect 19349 11305 19383 11339
rect 20177 11305 20211 11339
rect 1961 11237 1995 11271
rect 7205 11237 7239 11271
rect 10333 11237 10367 11271
rect 12541 11237 12575 11271
rect 12909 11237 12943 11271
rect 13093 11237 13127 11271
rect 14657 11237 14691 11271
rect 15761 11237 15795 11271
rect 8953 11169 8987 11203
rect 11161 11169 11195 11203
rect 15209 11169 15243 11203
rect 15301 11169 15335 11203
rect 16313 11169 16347 11203
rect 16405 11169 16439 11203
rect 17601 11169 17635 11203
rect 19901 11169 19935 11203
rect 20729 11169 20763 11203
rect 2145 11101 2179 11135
rect 2513 11101 2547 11135
rect 2697 11101 2731 11135
rect 4353 11101 4387 11135
rect 5825 11101 5859 11135
rect 7297 11101 7331 11135
rect 9220 11101 9254 11135
rect 16865 11101 16899 11135
rect 17509 11101 17543 11135
rect 17969 11101 18003 11135
rect 19717 11101 19751 11135
rect 20637 11101 20671 11135
rect 21281 11101 21315 11135
rect 2881 11033 2915 11067
rect 4620 11033 4654 11067
rect 6070 11033 6104 11067
rect 7542 11033 7576 11067
rect 11428 11033 11462 11067
rect 14841 11033 14875 11067
rect 15393 11033 15427 11067
rect 16221 11033 16255 11067
rect 17417 11033 17451 11067
rect 18337 11033 18371 11067
rect 18429 11033 18463 11067
rect 5733 10965 5767 10999
rect 8677 10965 8711 10999
rect 10425 10965 10459 10999
rect 15853 10965 15887 10999
rect 18061 10965 18095 10999
rect 19809 10965 19843 10999
rect 20545 10965 20579 10999
rect 21005 10965 21039 10999
rect 21465 10965 21499 10999
rect 14565 10761 14599 10795
rect 15485 10761 15519 10795
rect 15669 10761 15703 10795
rect 16957 10761 16991 10795
rect 19901 10761 19935 10795
rect 20545 10761 20579 10795
rect 20913 10761 20947 10795
rect 7266 10693 7300 10727
rect 18153 10693 18187 10727
rect 20361 10693 20395 10727
rect 4454 10625 4488 10659
rect 4721 10625 4755 10659
rect 5937 10625 5971 10659
rect 8493 10625 8527 10659
rect 8760 10625 8794 10659
rect 9965 10625 9999 10659
rect 10232 10625 10266 10659
rect 12642 10625 12676 10659
rect 12909 10625 12943 10659
rect 14114 10625 14148 10659
rect 14381 10625 14415 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 21005 10625 21039 10659
rect 21373 10625 21407 10659
rect 6193 10557 6227 10591
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 7021 10557 7055 10591
rect 16773 10557 16807 10591
rect 19993 10557 20027 10591
rect 20085 10557 20119 10591
rect 21097 10557 21131 10591
rect 4813 10489 4847 10523
rect 19441 10489 19475 10523
rect 3341 10421 3375 10455
rect 6929 10421 6963 10455
rect 8401 10421 8435 10455
rect 9873 10421 9907 10455
rect 11345 10421 11379 10455
rect 11529 10421 11563 10455
rect 13001 10421 13035 10455
rect 14749 10421 14783 10455
rect 17417 10421 17451 10455
rect 19533 10421 19567 10455
rect 2697 10217 2731 10251
rect 6929 10217 6963 10251
rect 7297 10217 7331 10251
rect 9045 10217 9079 10251
rect 9689 10217 9723 10251
rect 12817 10217 12851 10251
rect 15945 10217 15979 10251
rect 16865 10217 16899 10251
rect 16957 10217 16991 10251
rect 17969 10217 18003 10251
rect 20269 10217 20303 10251
rect 21281 10217 21315 10251
rect 7021 10149 7055 10183
rect 8769 10149 8803 10183
rect 14841 10149 14875 10183
rect 21465 10149 21499 10183
rect 3341 10081 3375 10115
rect 7389 10081 7423 10115
rect 11161 10081 11195 10115
rect 12633 10081 12667 10115
rect 13277 10081 13311 10115
rect 14197 10081 14231 10115
rect 14381 10081 14415 10115
rect 15485 10081 15519 10115
rect 16221 10081 16255 10115
rect 16405 10081 16439 10115
rect 17509 10081 17543 10115
rect 18521 10081 18555 10115
rect 20821 10081 20855 10115
rect 5006 10013 5040 10047
rect 5273 10013 5307 10047
rect 5365 10013 5399 10047
rect 5632 10013 5666 10047
rect 10905 10013 10939 10047
rect 17325 10013 17359 10047
rect 18337 10013 18371 10047
rect 19349 10013 19383 10047
rect 20085 10013 20119 10047
rect 20729 10013 20763 10047
rect 21097 10013 21131 10047
rect 7656 9945 7690 9979
rect 12388 9945 12422 9979
rect 13553 9945 13587 9979
rect 14473 9945 14507 9979
rect 15393 9945 15427 9979
rect 16497 9945 16531 9979
rect 19625 9945 19659 9979
rect 2421 9877 2455 9911
rect 3065 9877 3099 9911
rect 3157 9877 3191 9911
rect 3893 9877 3927 9911
rect 6745 9877 6779 9911
rect 9781 9877 9815 9911
rect 11253 9877 11287 9911
rect 13001 9877 13035 9911
rect 13461 9877 13495 9911
rect 13921 9877 13955 9911
rect 14933 9877 14967 9911
rect 15301 9877 15335 9911
rect 15853 9877 15887 9911
rect 17417 9877 17451 9911
rect 17877 9877 17911 9911
rect 18429 9877 18463 9911
rect 18889 9877 18923 9911
rect 19901 9877 19935 9911
rect 20637 9877 20671 9911
rect 3341 9673 3375 9707
rect 4261 9673 4295 9707
rect 4353 9673 4387 9707
rect 4905 9673 4939 9707
rect 5825 9673 5859 9707
rect 9505 9673 9539 9707
rect 11069 9673 11103 9707
rect 11253 9673 11287 9707
rect 14197 9673 14231 9707
rect 18705 9673 18739 9707
rect 20729 9673 20763 9707
rect 2973 9605 3007 9639
rect 3709 9605 3743 9639
rect 9864 9605 9898 9639
rect 15025 9605 15059 9639
rect 16129 9605 16163 9639
rect 17141 9605 17175 9639
rect 18245 9605 18279 9639
rect 19349 9605 19383 9639
rect 20269 9605 20303 9639
rect 2053 9537 2087 9571
rect 2881 9537 2915 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 7196 9537 7230 9571
rect 9597 9537 9631 9571
rect 12642 9537 12676 9571
rect 12909 9537 12943 9571
rect 14749 9537 14783 9571
rect 16221 9537 16255 9571
rect 17049 9537 17083 9571
rect 18337 9537 18371 9571
rect 20177 9537 20211 9571
rect 20821 9537 20855 9571
rect 21189 9537 21223 9571
rect 1777 9469 1811 9503
rect 1961 9469 1995 9503
rect 3157 9469 3191 9503
rect 4077 9469 4111 9503
rect 5181 9469 5215 9503
rect 13921 9469 13955 9503
rect 14105 9469 14139 9503
rect 16405 9469 16439 9503
rect 17233 9469 17267 9503
rect 18153 9469 18187 9503
rect 19441 9469 19475 9503
rect 19625 9469 19659 9503
rect 20361 9469 20395 9503
rect 2421 9401 2455 9435
rect 2513 9401 2547 9435
rect 11529 9401 11563 9435
rect 14565 9401 14599 9435
rect 19809 9401 19843 9435
rect 21005 9401 21039 9435
rect 21373 9401 21407 9435
rect 4721 9333 4755 9367
rect 8309 9333 8343 9367
rect 10977 9333 11011 9367
rect 13645 9333 13679 9367
rect 15761 9333 15795 9367
rect 16681 9333 16715 9367
rect 17877 9333 17911 9367
rect 18797 9333 18831 9367
rect 18981 9333 19015 9367
rect 1961 9129 1995 9163
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 5089 9129 5123 9163
rect 5273 9129 5307 9163
rect 14381 9129 14415 9163
rect 16865 9129 16899 9163
rect 21281 9129 21315 9163
rect 21465 9061 21499 9095
rect 5825 8993 5859 9027
rect 6561 8993 6595 9027
rect 6745 8993 6779 9027
rect 7481 8993 7515 9027
rect 12817 8993 12851 9027
rect 16221 8993 16255 9027
rect 16405 8993 16439 9027
rect 18337 8993 18371 9027
rect 19073 8993 19107 9027
rect 19441 8993 19475 9027
rect 20085 8993 20119 9027
rect 20637 8993 20671 9027
rect 2145 8925 2179 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 6469 8925 6503 8959
rect 7389 8925 7423 8959
rect 18153 8925 18187 8959
rect 19901 8925 19935 8959
rect 20361 8925 20395 8959
rect 7297 8857 7331 8891
rect 7757 8857 7791 8891
rect 13093 8857 13127 8891
rect 13553 8857 13587 8891
rect 14565 8857 14599 8891
rect 16497 8857 16531 8891
rect 18245 8857 18279 8891
rect 21097 8857 21131 8891
rect 3985 8789 4019 8823
rect 4905 8789 4939 8823
rect 5641 8789 5675 8823
rect 5733 8789 5767 8823
rect 6101 8789 6135 8823
rect 6929 8789 6963 8823
rect 13001 8789 13035 8823
rect 13461 8789 13495 8823
rect 14105 8789 14139 8823
rect 14749 8789 14783 8823
rect 17785 8789 17819 8823
rect 19533 8789 19567 8823
rect 19993 8789 20027 8823
rect 20913 8789 20947 8823
rect 1961 8585 1995 8619
rect 3249 8585 3283 8619
rect 3709 8585 3743 8619
rect 4997 8585 5031 8619
rect 6101 8585 6135 8619
rect 13737 8585 13771 8619
rect 14105 8585 14139 8619
rect 14473 8585 14507 8619
rect 14933 8585 14967 8619
rect 18889 8585 18923 8619
rect 21005 8585 21039 8619
rect 21373 8585 21407 8619
rect 2329 8517 2363 8551
rect 3617 8517 3651 8551
rect 4445 8517 4479 8551
rect 13369 8517 13403 8551
rect 15393 8517 15427 8551
rect 18797 8517 18831 8551
rect 2145 8449 2179 8483
rect 5365 8449 5399 8483
rect 5457 8449 5491 8483
rect 5917 8449 5951 8483
rect 15301 8449 15335 8483
rect 15761 8449 15795 8483
rect 19257 8449 19291 8483
rect 20269 8449 20303 8483
rect 20821 8449 20855 8483
rect 21189 8449 21223 8483
rect 3893 8381 3927 8415
rect 4537 8381 4571 8415
rect 4721 8381 4755 8415
rect 5641 8381 5675 8415
rect 6469 8381 6503 8415
rect 12909 8381 12943 8415
rect 13185 8381 13219 8415
rect 13277 8381 13311 8415
rect 13829 8381 13863 8415
rect 14565 8381 14599 8415
rect 14657 8381 14691 8415
rect 15485 8381 15519 8415
rect 19349 8381 19383 8415
rect 19441 8381 19475 8415
rect 20545 8381 20579 8415
rect 4077 8313 4111 8347
rect 19717 8313 19751 8347
rect 20085 8313 20119 8347
rect 19993 8245 20027 8279
rect 2237 8041 2271 8075
rect 13829 8041 13863 8075
rect 14841 8041 14875 8075
rect 15209 8041 15243 8075
rect 18613 8041 18647 8075
rect 19533 8041 19567 8075
rect 21373 8041 21407 8075
rect 17509 7973 17543 8007
rect 21005 7973 21039 8007
rect 1961 7905 1995 7939
rect 2881 7905 2915 7939
rect 4353 7905 4387 7939
rect 4537 7905 4571 7939
rect 5181 7905 5215 7939
rect 6469 7905 6503 7939
rect 9597 7905 9631 7939
rect 14197 7905 14231 7939
rect 16865 7905 16899 7939
rect 18061 7905 18095 7939
rect 18153 7905 18187 7939
rect 20177 7905 20211 7939
rect 20269 7905 20303 7939
rect 2145 7837 2179 7871
rect 5273 7837 5307 7871
rect 14381 7837 14415 7871
rect 15025 7837 15059 7871
rect 18797 7837 18831 7871
rect 19349 7837 19383 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 21189 7837 21223 7871
rect 2605 7769 2639 7803
rect 3065 7769 3099 7803
rect 3617 7769 3651 7803
rect 5365 7769 5399 7803
rect 14473 7769 14507 7803
rect 17049 7769 17083 7803
rect 18429 7769 18463 7803
rect 20085 7769 20119 7803
rect 1593 7701 1627 7735
rect 2697 7701 2731 7735
rect 3893 7701 3927 7735
rect 4261 7701 4295 7735
rect 4905 7701 4939 7735
rect 5733 7701 5767 7735
rect 5825 7701 5859 7735
rect 6193 7701 6227 7735
rect 6285 7701 6319 7735
rect 6745 7701 6779 7735
rect 9689 7701 9723 7735
rect 9781 7701 9815 7735
rect 10149 7701 10183 7735
rect 17141 7701 17175 7735
rect 17601 7701 17635 7735
rect 17969 7701 18003 7735
rect 18981 7701 19015 7735
rect 19717 7701 19751 7735
rect 2053 7497 2087 7531
rect 4353 7497 4387 7531
rect 5273 7497 5307 7531
rect 10333 7497 10367 7531
rect 10701 7497 10735 7531
rect 15945 7497 15979 7531
rect 16405 7497 16439 7531
rect 16957 7497 16991 7531
rect 17049 7497 17083 7531
rect 17509 7497 17543 7531
rect 17969 7497 18003 7531
rect 19165 7497 19199 7531
rect 20361 7497 20395 7531
rect 20453 7497 20487 7531
rect 3985 7429 4019 7463
rect 7113 7429 7147 7463
rect 16037 7429 16071 7463
rect 18797 7429 18831 7463
rect 21189 7429 21223 7463
rect 2237 7361 2271 7395
rect 4261 7361 4295 7395
rect 4721 7361 4755 7395
rect 9965 7361 9999 7395
rect 17877 7361 17911 7395
rect 18705 7361 18739 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 21005 7361 21039 7395
rect 3709 7293 3743 7327
rect 4813 7293 4847 7327
rect 4997 7293 5031 7327
rect 7205 7293 7239 7327
rect 7389 7293 7423 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 15761 7293 15795 7327
rect 16773 7293 16807 7327
rect 18061 7293 18095 7327
rect 18889 7293 18923 7327
rect 19717 7293 19751 7327
rect 20545 7293 20579 7327
rect 5641 7225 5675 7259
rect 17417 7225 17451 7259
rect 21373 7225 21407 7259
rect 6745 7157 6779 7191
rect 10149 7157 10183 7191
rect 18337 7157 18371 7191
rect 19993 7157 20027 7191
rect 20821 7157 20855 7191
rect 2605 6953 2639 6987
rect 17601 6953 17635 6987
rect 19257 6953 19291 6987
rect 20085 6953 20119 6987
rect 21005 6885 21039 6919
rect 3157 6817 3191 6851
rect 4169 6817 4203 6851
rect 4721 6817 4755 6851
rect 5549 6817 5583 6851
rect 5733 6817 5767 6851
rect 10701 6817 10735 6851
rect 18245 6817 18279 6851
rect 19073 6817 19107 6851
rect 19717 6817 19751 6851
rect 19901 6817 19935 6851
rect 20913 6817 20947 6851
rect 4445 6749 4479 6783
rect 19625 6749 19659 6783
rect 17417 6681 17451 6715
rect 17969 6681 18003 6715
rect 18429 6681 18463 6715
rect 2973 6613 3007 6647
rect 3065 6613 3099 6647
rect 5089 6613 5123 6647
rect 5457 6613 5491 6647
rect 18061 6613 18095 6647
rect 18705 6613 18739 6647
rect 21189 6613 21223 6647
rect 3341 6409 3375 6443
rect 3617 6409 3651 6443
rect 3985 6409 4019 6443
rect 4077 6409 4111 6443
rect 4445 6409 4479 6443
rect 4905 6409 4939 6443
rect 5733 6409 5767 6443
rect 6377 6409 6411 6443
rect 6837 6409 6871 6443
rect 8217 6409 8251 6443
rect 9229 6409 9263 6443
rect 9965 6409 9999 6443
rect 12081 6409 12115 6443
rect 12541 6409 12575 6443
rect 13921 6409 13955 6443
rect 16957 6409 16991 6443
rect 17325 6409 17359 6443
rect 17785 6409 17819 6443
rect 18153 6409 18187 6443
rect 18245 6409 18279 6443
rect 18613 6409 18647 6443
rect 19073 6409 19107 6443
rect 19717 6409 19751 6443
rect 4813 6341 4847 6375
rect 10793 6341 10827 6375
rect 11989 6341 12023 6375
rect 13093 6341 13127 6375
rect 19993 6341 20027 6375
rect 2973 6273 3007 6307
rect 5641 6273 5675 6307
rect 6745 6273 6779 6307
rect 8861 6273 8895 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 12449 6273 12483 6307
rect 13001 6273 13035 6307
rect 14289 6273 14323 6307
rect 18981 6273 19015 6307
rect 2697 6205 2731 6239
rect 2881 6205 2915 6239
rect 4169 6205 4203 6239
rect 4997 6205 5031 6239
rect 5825 6205 5859 6239
rect 6929 6205 6963 6239
rect 8585 6205 8619 6239
rect 8769 6205 8803 6239
rect 10517 6205 10551 6239
rect 11069 6205 11103 6239
rect 12633 6205 12667 6239
rect 14381 6205 14415 6239
rect 14473 6205 14507 6239
rect 17417 6205 17451 6239
rect 17509 6205 17543 6239
rect 18337 6205 18371 6239
rect 19165 6205 19199 6239
rect 5273 6137 5307 6171
rect 9321 6137 9355 6171
rect 8309 6069 8343 6103
rect 13829 6069 13863 6103
rect 14841 6069 14875 6103
rect 19533 6069 19567 6103
rect 2697 5865 2731 5899
rect 19257 5865 19291 5899
rect 6377 5797 6411 5831
rect 3341 5729 3375 5763
rect 6193 5729 6227 5763
rect 6929 5729 6963 5763
rect 19809 5729 19843 5763
rect 20637 5729 20671 5763
rect 5825 5661 5859 5695
rect 6745 5661 6779 5695
rect 2605 5593 2639 5627
rect 3065 5593 3099 5627
rect 6101 5593 6135 5627
rect 19625 5593 19659 5627
rect 20453 5593 20487 5627
rect 2237 5525 2271 5559
rect 3157 5525 3191 5559
rect 6837 5525 6871 5559
rect 7297 5525 7331 5559
rect 19717 5525 19751 5559
rect 20085 5525 20119 5559
rect 20545 5525 20579 5559
rect 20913 5525 20947 5559
rect 21189 5525 21223 5559
rect 3249 5321 3283 5355
rect 6193 5321 6227 5355
rect 7113 5321 7147 5355
rect 7205 5321 7239 5355
rect 19441 5321 19475 5355
rect 2789 5253 2823 5287
rect 5825 5253 5859 5287
rect 19349 5253 19383 5287
rect 2881 5185 2915 5219
rect 3801 5185 3835 5219
rect 4445 5185 4479 5219
rect 6745 5185 6779 5219
rect 7573 5185 7607 5219
rect 8033 5185 8067 5219
rect 19809 5185 19843 5219
rect 2697 5117 2731 5151
rect 4537 5117 4571 5151
rect 4721 5117 4755 5151
rect 5549 5117 5583 5151
rect 5733 5117 5767 5151
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 7665 5117 7699 5151
rect 7757 5117 7791 5151
rect 19901 5117 19935 5151
rect 19993 5117 20027 5151
rect 2237 5049 2271 5083
rect 3893 5049 3927 5083
rect 2329 4981 2363 5015
rect 4077 4981 4111 5015
rect 4997 4981 5031 5015
rect 20361 4981 20395 5015
rect 20545 4981 20579 5015
rect 3985 4777 4019 4811
rect 5273 4777 5307 4811
rect 6377 4777 6411 4811
rect 7297 4777 7331 4811
rect 4629 4641 4663 4675
rect 5917 4641 5951 4675
rect 7021 4641 7055 4675
rect 7481 4641 7515 4675
rect 3249 4573 3283 4607
rect 4813 4573 4847 4607
rect 6745 4573 6779 4607
rect 3157 4505 3191 4539
rect 4721 4505 4755 4539
rect 5733 4505 5767 4539
rect 6837 4505 6871 4539
rect 7665 4505 7699 4539
rect 3893 4437 3927 4471
rect 4353 4437 4387 4471
rect 5181 4437 5215 4471
rect 5641 4437 5675 4471
rect 6101 4437 6135 4471
rect 3801 4233 3835 4267
rect 5273 4233 5307 4267
rect 5825 4233 5859 4267
rect 6469 4233 6503 4267
rect 4721 4165 4755 4199
rect 2973 4097 3007 4131
rect 4353 4097 4387 4131
rect 4813 4097 4847 4131
rect 5917 4097 5951 4131
rect 2697 4029 2731 4063
rect 2881 4029 2915 4063
rect 3893 4029 3927 4063
rect 4077 4029 4111 4063
rect 4537 4029 4571 4063
rect 6009 4029 6043 4063
rect 3341 3961 3375 3995
rect 5181 3961 5215 3995
rect 5457 3961 5491 3995
rect 3433 3893 3467 3927
rect 2145 3689 2179 3723
rect 2329 3689 2363 3723
rect 3249 3689 3283 3723
rect 4721 3689 4755 3723
rect 5733 3689 5767 3723
rect 5917 3689 5951 3723
rect 2697 3553 2731 3587
rect 4077 3553 4111 3587
rect 4261 3553 4295 3587
rect 5181 3553 5215 3587
rect 2881 3485 2915 3519
rect 4353 3485 4387 3519
rect 5365 3485 5399 3519
rect 2789 3417 2823 3451
rect 3433 3417 3467 3451
rect 4813 3349 4847 3383
rect 5273 3349 5307 3383
rect 3617 3145 3651 3179
rect 3249 3077 3283 3111
rect 3985 3077 4019 3111
rect 4537 3077 4571 3111
rect 5273 3077 5307 3111
rect 18889 3077 18923 3111
rect 5549 3009 5583 3043
rect 12265 3009 12299 3043
rect 12541 3009 12575 3043
rect 19165 3009 19199 3043
rect 3433 2941 3467 2975
rect 4077 2941 4111 2975
rect 4261 2941 4295 2975
rect 4629 2805 4663 2839
rect 5733 2805 5767 2839
rect 12725 2805 12759 2839
rect 19349 2805 19383 2839
<< metal1 >>
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 7374 21060 7380 21072
rect 5224 21032 7380 21060
rect 5224 21020 5230 21032
rect 7374 21020 7380 21032
rect 7432 21020 7438 21072
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 11054 20992 11060 21004
rect 3936 20964 11060 20992
rect 3936 20952 3942 20964
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 2958 20884 2964 20936
rect 3016 20924 3022 20936
rect 16206 20924 16212 20936
rect 3016 20896 16212 20924
rect 3016 20884 3022 20896
rect 16206 20884 16212 20896
rect 16264 20884 16270 20936
rect 1670 20816 1676 20868
rect 1728 20856 1734 20868
rect 1728 20828 2774 20856
rect 1728 20816 1734 20828
rect 2746 20788 2774 20828
rect 5810 20816 5816 20868
rect 5868 20856 5874 20868
rect 6822 20856 6828 20868
rect 5868 20828 6828 20856
rect 5868 20816 5874 20828
rect 6822 20816 6828 20828
rect 6880 20816 6886 20868
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 15102 20856 15108 20868
rect 13872 20828 15108 20856
rect 13872 20816 13878 20828
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 20162 20788 20168 20800
rect 2746 20760 20168 20788
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 2866 20584 2872 20596
rect 2827 20556 2872 20584
rect 2866 20544 2872 20556
rect 2924 20584 2930 20596
rect 3329 20587 3387 20593
rect 3329 20584 3341 20587
rect 2924 20556 3341 20584
rect 2924 20544 2930 20556
rect 3329 20553 3341 20556
rect 3375 20584 3387 20587
rect 4430 20584 4436 20596
rect 3375 20556 4436 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4801 20587 4859 20593
rect 4801 20553 4813 20587
rect 4847 20584 4859 20587
rect 4847 20556 6132 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 2038 20476 2044 20528
rect 2096 20516 2102 20528
rect 2961 20519 3019 20525
rect 2961 20516 2973 20519
rect 2096 20488 2973 20516
rect 2096 20476 2102 20488
rect 2961 20485 2973 20488
rect 3007 20485 3019 20519
rect 2961 20479 3019 20485
rect 3237 20519 3295 20525
rect 3237 20485 3249 20519
rect 3283 20516 3295 20519
rect 6104 20516 6132 20556
rect 6178 20544 6184 20596
rect 6236 20584 6242 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 6236 20556 6377 20584
rect 6236 20544 6242 20556
rect 6365 20553 6377 20556
rect 6411 20553 6423 20587
rect 6365 20547 6423 20553
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 7190 20584 7196 20596
rect 6687 20556 7196 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 7374 20544 7380 20596
rect 7432 20584 7438 20596
rect 7837 20587 7895 20593
rect 7432 20556 7477 20584
rect 7432 20544 7438 20556
rect 7837 20553 7849 20587
rect 7883 20584 7895 20587
rect 9217 20587 9275 20593
rect 9217 20584 9229 20587
rect 7883 20556 9229 20584
rect 7883 20553 7895 20556
rect 7837 20547 7895 20553
rect 9217 20553 9229 20556
rect 9263 20553 9275 20587
rect 9217 20547 9275 20553
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 9582 20584 9588 20596
rect 9364 20556 9588 20584
rect 9364 20544 9370 20556
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 9677 20587 9735 20593
rect 9677 20553 9689 20587
rect 9723 20584 9735 20587
rect 10042 20584 10048 20596
rect 9723 20556 10048 20584
rect 9723 20553 9735 20556
rect 9677 20547 9735 20553
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10183 20556 10609 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 15562 20584 15568 20596
rect 10597 20547 10655 20553
rect 10704 20556 15568 20584
rect 6730 20516 6736 20528
rect 3283 20488 5028 20516
rect 6104 20488 6736 20516
rect 3283 20485 3295 20488
rect 3237 20479 3295 20485
rect 2976 20448 3004 20479
rect 5000 20460 5028 20488
rect 6730 20476 6736 20488
rect 6788 20476 6794 20528
rect 7006 20516 7012 20528
rect 6919 20488 7012 20516
rect 3513 20451 3571 20457
rect 3513 20448 3525 20451
rect 2976 20420 3525 20448
rect 3513 20417 3525 20420
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20448 4031 20451
rect 4246 20448 4252 20460
rect 4019 20420 4252 20448
rect 4019 20417 4031 20420
rect 3973 20411 4031 20417
rect 3528 20312 3556 20411
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 4982 20448 4988 20460
rect 4943 20420 4988 20448
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 6181 20451 6239 20457
rect 6181 20417 6193 20451
rect 6227 20448 6239 20451
rect 6932 20448 6960 20488
rect 7006 20476 7012 20488
rect 7064 20516 7070 20528
rect 7466 20516 7472 20528
rect 7064 20488 7144 20516
rect 7427 20488 7472 20516
rect 7064 20476 7070 20488
rect 6227 20420 6960 20448
rect 7116 20448 7144 20488
rect 7466 20476 7472 20488
rect 7524 20516 7530 20528
rect 7742 20516 7748 20528
rect 7524 20488 7748 20516
rect 7524 20476 7530 20488
rect 7742 20476 7748 20488
rect 7800 20476 7806 20528
rect 8202 20516 8208 20528
rect 8163 20488 8208 20516
rect 8202 20476 8208 20488
rect 8260 20476 8266 20528
rect 10704 20516 10732 20556
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 15749 20587 15807 20593
rect 15749 20553 15761 20587
rect 15795 20584 15807 20587
rect 16022 20584 16028 20596
rect 15795 20556 16028 20584
rect 15795 20553 15807 20556
rect 15749 20547 15807 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 16301 20587 16359 20593
rect 16301 20553 16313 20587
rect 16347 20584 16359 20587
rect 16390 20584 16396 20596
rect 16347 20556 16396 20584
rect 16347 20553 16359 20556
rect 16301 20547 16359 20553
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 19334 20584 19340 20596
rect 16899 20556 19340 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 11054 20516 11060 20528
rect 8404 20488 10732 20516
rect 10967 20488 11060 20516
rect 7116 20420 7236 20448
rect 6227 20417 6239 20420
rect 6181 20411 6239 20417
rect 4154 20380 4160 20392
rect 4115 20352 4160 20380
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20380 4399 20383
rect 5166 20380 5172 20392
rect 4387 20352 5172 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 4356 20312 4384 20343
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 7208 20389 7236 20420
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 8297 20451 8355 20457
rect 8297 20448 8309 20451
rect 7708 20420 8309 20448
rect 7708 20408 7714 20420
rect 8297 20417 8309 20420
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 5261 20383 5319 20389
rect 5261 20349 5273 20383
rect 5307 20349 5319 20383
rect 5261 20343 5319 20349
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20349 7251 20383
rect 8018 20380 8024 20392
rect 7979 20352 8024 20380
rect 7193 20343 7251 20349
rect 3528 20284 4384 20312
rect 4430 20272 4436 20324
rect 4488 20312 4494 20324
rect 5276 20312 5304 20343
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 8110 20340 8116 20392
rect 8168 20380 8174 20392
rect 8404 20380 8432 20488
rect 11054 20476 11060 20488
rect 11112 20516 11118 20528
rect 11793 20519 11851 20525
rect 11793 20516 11805 20519
rect 11112 20488 11805 20516
rect 11112 20476 11118 20488
rect 11793 20485 11805 20488
rect 11839 20516 11851 20519
rect 12894 20516 12900 20528
rect 11839 20488 12900 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 12894 20476 12900 20488
rect 12952 20476 12958 20528
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 13446 20516 13452 20528
rect 13044 20488 13452 20516
rect 13044 20476 13050 20488
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 14461 20519 14519 20525
rect 14461 20516 14473 20519
rect 13596 20488 14473 20516
rect 13596 20476 13602 20488
rect 14461 20485 14473 20488
rect 14507 20516 14519 20519
rect 14734 20516 14740 20528
rect 14507 20488 14740 20516
rect 14507 20485 14519 20488
rect 14461 20479 14519 20485
rect 14734 20476 14740 20488
rect 14792 20476 14798 20528
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 9122 20448 9128 20460
rect 8720 20420 9128 20448
rect 8720 20408 8726 20420
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 9306 20448 9312 20460
rect 9267 20420 9312 20448
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 10962 20448 10968 20460
rect 10923 20420 10968 20448
rect 10962 20408 10968 20420
rect 11020 20448 11026 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11020 20420 11897 20448
rect 11020 20408 11026 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20448 12403 20451
rect 12434 20448 12440 20460
rect 12391 20420 12440 20448
rect 12391 20417 12403 20420
rect 12345 20411 12403 20417
rect 8168 20352 8432 20380
rect 9033 20383 9091 20389
rect 8168 20340 8174 20352
rect 9033 20349 9045 20383
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 4488 20284 5304 20312
rect 6825 20315 6883 20321
rect 4488 20272 4494 20284
rect 6825 20281 6837 20315
rect 6871 20312 6883 20315
rect 7466 20312 7472 20324
rect 6871 20284 7472 20312
rect 6871 20281 6883 20284
rect 6825 20275 6883 20281
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 8202 20272 8208 20324
rect 8260 20312 8266 20324
rect 9048 20312 9076 20343
rect 9858 20340 9864 20392
rect 9916 20380 9922 20392
rect 10045 20383 10103 20389
rect 9916 20352 9961 20380
rect 9916 20340 9922 20352
rect 10045 20349 10057 20383
rect 10091 20380 10103 20383
rect 10870 20380 10876 20392
rect 10091 20352 10876 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 11241 20383 11299 20389
rect 11241 20349 11253 20383
rect 11287 20380 11299 20383
rect 11514 20380 11520 20392
rect 11287 20352 11520 20380
rect 11287 20349 11299 20352
rect 11241 20343 11299 20349
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 11900 20380 11928 20411
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 15010 20408 15016 20460
rect 15068 20448 15074 20460
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15068 20420 15577 20448
rect 15068 20408 15074 20420
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15896 20420 16129 20448
rect 15896 20408 15902 20420
rect 16117 20417 16129 20420
rect 16163 20417 16175 20451
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16117 20411 16175 20417
rect 16666 20408 16672 20420
rect 16724 20448 16730 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16724 20420 17049 20448
rect 16724 20408 16730 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 11900 20352 13829 20380
rect 13817 20349 13829 20352
rect 13863 20380 13875 20383
rect 14366 20380 14372 20392
rect 13863 20352 14372 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20380 14611 20383
rect 14642 20380 14648 20392
rect 14599 20352 14648 20380
rect 14599 20349 14611 20352
rect 14553 20343 14611 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20349 14795 20383
rect 14737 20343 14795 20349
rect 9490 20312 9496 20324
rect 8260 20284 9076 20312
rect 9324 20284 9496 20312
rect 8260 20272 8266 20284
rect 6546 20204 6552 20256
rect 6604 20244 6610 20256
rect 6914 20244 6920 20256
rect 6604 20216 6920 20244
rect 6604 20204 6610 20216
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7834 20244 7840 20256
rect 7432 20216 7840 20244
rect 7432 20204 7438 20216
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8665 20247 8723 20253
rect 8665 20213 8677 20247
rect 8711 20244 8723 20247
rect 9324 20244 9352 20284
rect 9490 20272 9496 20284
rect 9548 20272 9554 20324
rect 10505 20315 10563 20321
rect 10505 20281 10517 20315
rect 10551 20312 10563 20315
rect 13078 20312 13084 20324
rect 10551 20284 13084 20312
rect 10551 20281 10563 20284
rect 10505 20275 10563 20281
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 13446 20312 13452 20324
rect 13407 20284 13452 20312
rect 13446 20272 13452 20284
rect 13504 20312 13510 20324
rect 13633 20315 13691 20321
rect 13633 20312 13645 20315
rect 13504 20284 13645 20312
rect 13504 20272 13510 20284
rect 13633 20281 13645 20284
rect 13679 20312 13691 20315
rect 14752 20312 14780 20343
rect 14826 20312 14832 20324
rect 13679 20284 14832 20312
rect 13679 20281 13691 20284
rect 13633 20275 13691 20281
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 16390 20272 16396 20324
rect 16448 20312 16454 20324
rect 16448 20284 20760 20312
rect 16448 20272 16454 20284
rect 20732 20256 20760 20284
rect 8711 20216 9352 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 11514 20244 11520 20256
rect 9456 20216 11520 20244
rect 9456 20204 9462 20216
rect 11514 20204 11520 20216
rect 11572 20204 11578 20256
rect 11974 20204 11980 20256
rect 12032 20244 12038 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 12032 20216 12081 20244
rect 12032 20204 12038 20216
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 12069 20207 12127 20213
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 12989 20247 13047 20253
rect 12989 20244 13001 20247
rect 12492 20216 13001 20244
rect 12492 20204 12498 20216
rect 12989 20213 13001 20216
rect 13035 20244 13047 20247
rect 13170 20244 13176 20256
rect 13035 20216 13176 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13538 20244 13544 20256
rect 13320 20216 13544 20244
rect 13320 20204 13326 20216
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14093 20247 14151 20253
rect 14093 20244 14105 20247
rect 13872 20216 14105 20244
rect 13872 20204 13878 20216
rect 14093 20213 14105 20216
rect 14139 20213 14151 20247
rect 16022 20244 16028 20256
rect 15983 20216 16028 20244
rect 14093 20207 14151 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17954 20244 17960 20256
rect 16632 20216 17960 20244
rect 16632 20204 16638 20216
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 20714 20244 20720 20256
rect 20675 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21085 20247 21143 20253
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 21266 20244 21272 20256
rect 21131 20216 21272 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2317 20043 2375 20049
rect 2317 20009 2329 20043
rect 2363 20040 2375 20043
rect 2774 20040 2780 20052
rect 2363 20012 2780 20040
rect 2363 20009 2375 20012
rect 2317 20003 2375 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 2869 20043 2927 20049
rect 2869 20009 2881 20043
rect 2915 20040 2927 20043
rect 2958 20040 2964 20052
rect 2915 20012 2964 20040
rect 2915 20009 2927 20012
rect 2869 20003 2927 20009
rect 2884 19904 2912 20003
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 4246 20000 4252 20052
rect 4304 20040 4310 20052
rect 5534 20040 5540 20052
rect 4304 20012 5540 20040
rect 4304 20000 4310 20012
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 5684 20012 7205 20040
rect 5684 20000 5690 20012
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 7466 20000 7472 20052
rect 7524 20040 7530 20052
rect 10226 20040 10232 20052
rect 7524 20012 10232 20040
rect 7524 20000 7530 20012
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 11425 20043 11483 20049
rect 11425 20040 11437 20043
rect 10928 20012 11437 20040
rect 10928 20000 10934 20012
rect 11425 20009 11437 20012
rect 11471 20009 11483 20043
rect 11425 20003 11483 20009
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 13817 20043 13875 20049
rect 11572 20012 12020 20040
rect 11572 20000 11578 20012
rect 6822 19932 6828 19984
rect 6880 19972 6886 19984
rect 11054 19972 11060 19984
rect 6880 19944 9628 19972
rect 11015 19944 11060 19972
rect 6880 19932 6886 19944
rect 2148 19876 2912 19904
rect 6656 19876 7236 19904
rect 2148 19845 2176 19876
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 3421 19839 3479 19845
rect 2547 19808 2728 19836
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 2700 19712 2728 19808
rect 3421 19805 3433 19839
rect 3467 19836 3479 19839
rect 3881 19839 3939 19845
rect 3881 19836 3893 19839
rect 3467 19808 3893 19836
rect 3467 19805 3479 19808
rect 3421 19799 3479 19805
rect 3881 19805 3893 19808
rect 3927 19836 3939 19839
rect 4430 19836 4436 19848
rect 3927 19808 4436 19836
rect 3927 19805 3939 19808
rect 3881 19799 3939 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 6656 19836 6684 19876
rect 7208 19848 7236 19876
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 7745 19907 7803 19913
rect 7745 19904 7757 19907
rect 7432 19876 7757 19904
rect 7432 19864 7438 19876
rect 7745 19873 7757 19876
rect 7791 19873 7803 19907
rect 7745 19867 7803 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 9490 19904 9496 19916
rect 8251 19876 9496 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 9600 19904 9628 19944
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 11146 19932 11152 19984
rect 11204 19972 11210 19984
rect 11241 19975 11299 19981
rect 11241 19972 11253 19975
rect 11204 19944 11253 19972
rect 11204 19932 11210 19944
rect 11241 19941 11253 19944
rect 11287 19972 11299 19975
rect 11287 19944 11928 19972
rect 11287 19941 11299 19944
rect 11241 19935 11299 19941
rect 9600 19876 9720 19904
rect 4540 19808 6684 19836
rect 6733 19839 6791 19845
rect 3605 19771 3663 19777
rect 3605 19737 3617 19771
rect 3651 19768 3663 19771
rect 4148 19771 4206 19777
rect 4148 19768 4160 19771
rect 3651 19740 4160 19768
rect 3651 19737 3663 19740
rect 3605 19731 3663 19737
rect 4148 19737 4160 19740
rect 4194 19768 4206 19771
rect 4246 19768 4252 19780
rect 4194 19740 4252 19768
rect 4194 19737 4206 19740
rect 4148 19731 4206 19737
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 2682 19700 2688 19712
rect 2643 19672 2688 19700
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 3970 19660 3976 19712
rect 4028 19700 4034 19712
rect 4540 19700 4568 19808
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6914 19836 6920 19848
rect 6779 19808 6920 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 8297 19839 8355 19845
rect 8297 19836 8309 19839
rect 7248 19808 8309 19836
rect 7248 19796 7254 19808
rect 8297 19805 8309 19808
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 9214 19836 9220 19848
rect 8444 19808 9220 19836
rect 8444 19796 8450 19808
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19805 9643 19839
rect 9692 19836 9720 19876
rect 11072 19836 11100 19932
rect 11900 19913 11928 19944
rect 11992 19913 12020 20012
rect 13817 20009 13829 20043
rect 13863 20009 13875 20043
rect 14090 20040 14096 20052
rect 14051 20012 14096 20040
rect 13817 20003 13875 20009
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 12342 19972 12348 19984
rect 12216 19944 12348 19972
rect 12216 19932 12222 19944
rect 12342 19932 12348 19944
rect 12400 19932 12406 19984
rect 13446 19972 13452 19984
rect 12728 19944 13452 19972
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 9692 19808 11008 19836
rect 11072 19808 11805 19836
rect 9585 19799 9643 19805
rect 6488 19771 6546 19777
rect 5276 19740 6408 19768
rect 5276 19709 5304 19740
rect 4028 19672 4568 19700
rect 5261 19703 5319 19709
rect 4028 19660 4034 19672
rect 5261 19669 5273 19703
rect 5307 19669 5319 19703
rect 5261 19663 5319 19669
rect 5353 19703 5411 19709
rect 5353 19669 5365 19703
rect 5399 19700 5411 19703
rect 5534 19700 5540 19712
rect 5399 19672 5540 19700
rect 5399 19669 5411 19672
rect 5353 19663 5411 19669
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 6380 19700 6408 19740
rect 6488 19737 6500 19771
rect 6534 19768 6546 19771
rect 6534 19740 6776 19768
rect 6534 19737 6546 19740
rect 6488 19731 6546 19737
rect 6748 19712 6776 19740
rect 6932 19740 7696 19768
rect 6638 19700 6644 19712
rect 6380 19672 6644 19700
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 6730 19660 6736 19712
rect 6788 19660 6794 19712
rect 6932 19709 6960 19740
rect 7668 19712 7696 19740
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 9033 19771 9091 19777
rect 9033 19768 9045 19771
rect 8260 19740 9045 19768
rect 8260 19728 8266 19740
rect 9033 19737 9045 19740
rect 9079 19768 9091 19771
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 9079 19740 9413 19768
rect 9079 19737 9091 19740
rect 9033 19731 9091 19737
rect 9401 19737 9413 19740
rect 9447 19768 9459 19771
rect 9600 19768 9628 19799
rect 9830 19771 9888 19777
rect 9830 19768 9842 19771
rect 9447 19740 9628 19768
rect 9692 19740 9842 19768
rect 9447 19737 9459 19740
rect 9401 19731 9459 19737
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19669 6975 19703
rect 6917 19663 6975 19669
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 7374 19700 7380 19712
rect 7147 19672 7380 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 7466 19660 7472 19712
rect 7524 19700 7530 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 7524 19672 7573 19700
rect 7524 19660 7530 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7561 19663 7619 19669
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8754 19700 8760 19712
rect 7708 19672 7753 19700
rect 8715 19672 8760 19700
rect 7708 19660 7714 19672
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 8996 19672 9229 19700
rect 8996 19660 9002 19672
rect 9217 19669 9229 19672
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 9490 19660 9496 19712
rect 9548 19700 9554 19712
rect 9692 19700 9720 19740
rect 9830 19737 9842 19740
rect 9876 19737 9888 19771
rect 10980 19768 11008 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 11900 19836 11928 19867
rect 12342 19836 12348 19848
rect 11900 19808 12348 19836
rect 11793 19799 11851 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12526 19836 12532 19848
rect 12487 19808 12532 19836
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12728 19768 12756 19944
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 13832 19972 13860 20003
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 14608 20012 15485 20040
rect 14608 20000 14614 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15746 20040 15752 20052
rect 15659 20012 15752 20040
rect 15473 20003 15531 20009
rect 15746 20000 15752 20012
rect 15804 20040 15810 20052
rect 17773 20043 17831 20049
rect 15804 20012 17540 20040
rect 15804 20000 15810 20012
rect 15102 19972 15108 19984
rect 13832 19944 14964 19972
rect 15063 19944 15108 19972
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19904 13415 19907
rect 13814 19904 13820 19916
rect 13403 19876 13820 19904
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14608 19876 14749 19904
rect 14608 19864 14614 19876
rect 14737 19873 14749 19876
rect 14783 19904 14795 19907
rect 14826 19904 14832 19916
rect 14783 19876 14832 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 14936 19904 14964 19944
rect 15102 19932 15108 19944
rect 15160 19932 15166 19984
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 17402 19972 17408 19984
rect 15252 19944 17408 19972
rect 15252 19932 15258 19944
rect 17402 19932 17408 19944
rect 17460 19932 17466 19984
rect 17512 19972 17540 20012
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 17862 20040 17868 20052
rect 17819 20012 17868 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 18598 20040 18604 20052
rect 18279 20012 18604 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 19702 20000 19708 20052
rect 19760 20040 19766 20052
rect 19797 20043 19855 20049
rect 19797 20040 19809 20043
rect 19760 20012 19809 20040
rect 19760 20000 19766 20012
rect 19797 20009 19809 20012
rect 19843 20009 19855 20043
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 19797 20003 19855 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20533 20043 20591 20049
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 21174 20040 21180 20052
rect 20579 20012 21180 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 18138 19972 18144 19984
rect 17512 19944 18144 19972
rect 18138 19932 18144 19944
rect 18196 19932 18202 19984
rect 18969 19975 19027 19981
rect 18969 19941 18981 19975
rect 19015 19941 19027 19975
rect 20990 19972 20996 19984
rect 20951 19944 20996 19972
rect 18969 19935 19027 19941
rect 15470 19904 15476 19916
rect 14936 19876 15476 19904
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15620 19876 15945 19904
rect 15620 19864 15626 19876
rect 15933 19873 15945 19876
rect 15979 19904 15991 19907
rect 15979 19876 17908 19904
rect 15979 19873 15991 19876
rect 15933 19867 15991 19873
rect 13630 19796 13636 19848
rect 13688 19836 13694 19848
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 13688 19808 14933 19836
rect 13688 19796 13694 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 14921 19799 14979 19805
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 16206 19836 16212 19848
rect 16119 19808 16212 19836
rect 16206 19796 16212 19808
rect 16264 19836 16270 19848
rect 16758 19836 16764 19848
rect 16264 19808 16764 19836
rect 16264 19796 16270 19808
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 16853 19839 16911 19845
rect 16853 19805 16865 19839
rect 16899 19836 16911 19839
rect 16942 19836 16948 19848
rect 16899 19808 16948 19836
rect 16899 19805 16911 19808
rect 16853 19799 16911 19805
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17589 19839 17647 19845
rect 17589 19836 17601 19839
rect 17175 19808 17601 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 17589 19805 17601 19808
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 10980 19740 12756 19768
rect 9830 19731 9888 19737
rect 12894 19728 12900 19780
rect 12952 19768 12958 19780
rect 13449 19771 13507 19777
rect 12952 19740 13308 19768
rect 12952 19728 12958 19740
rect 9548 19672 9720 19700
rect 9548 19660 9554 19672
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 10965 19703 11023 19709
rect 10965 19700 10977 19703
rect 10928 19672 10977 19700
rect 10928 19660 10934 19672
rect 10965 19669 10977 19672
rect 11011 19669 11023 19703
rect 10965 19663 11023 19669
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12713 19703 12771 19709
rect 12492 19672 12537 19700
rect 12492 19660 12498 19672
rect 12713 19669 12725 19703
rect 12759 19700 12771 19703
rect 13170 19700 13176 19712
rect 12759 19672 13176 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13280 19700 13308 19740
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 14090 19768 14096 19780
rect 13495 19740 14096 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 14090 19728 14096 19740
rect 14148 19728 14154 19780
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 14461 19771 14519 19777
rect 14461 19768 14473 19771
rect 14424 19740 14473 19768
rect 14424 19728 14430 19740
rect 14461 19737 14473 19740
rect 14507 19768 14519 19771
rect 16022 19768 16028 19780
rect 14507 19740 16028 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 16022 19728 16028 19740
rect 16080 19768 16086 19780
rect 16117 19771 16175 19777
rect 16117 19768 16129 19771
rect 16080 19740 16129 19768
rect 16080 19728 16086 19740
rect 16117 19737 16129 19740
rect 16163 19737 16175 19771
rect 16117 19731 16175 19737
rect 17405 19771 17463 19777
rect 17405 19737 17417 19771
rect 17451 19768 17463 19771
rect 17678 19768 17684 19780
rect 17451 19740 17684 19768
rect 17451 19737 17463 19740
rect 17405 19731 17463 19737
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 17880 19768 17908 19876
rect 18230 19864 18236 19916
rect 18288 19904 18294 19916
rect 18984 19904 19012 19935
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 18288 19876 19012 19904
rect 18288 19864 18294 19876
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 18049 19839 18107 19845
rect 18049 19836 18061 19839
rect 18012 19808 18061 19836
rect 18012 19796 18018 19808
rect 18049 19805 18061 19808
rect 18095 19805 18107 19839
rect 18414 19836 18420 19848
rect 18375 19808 18420 19836
rect 18049 19799 18107 19805
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18782 19836 18788 19848
rect 18743 19808 18788 19836
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19536 19808 19625 19836
rect 18230 19768 18236 19780
rect 17880 19740 18236 19768
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 19536 19712 19564 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 20162 19796 20168 19848
rect 20220 19836 20226 19848
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 20220 19808 20361 19836
rect 20220 19796 20226 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 20809 19839 20867 19845
rect 20809 19836 20821 19839
rect 20772 19808 20821 19836
rect 20772 19796 20778 19808
rect 20809 19805 20821 19808
rect 20855 19836 20867 19839
rect 20990 19836 20996 19848
rect 20855 19808 20996 19836
rect 20855 19805 20867 19808
rect 20809 19799 20867 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21174 19836 21180 19848
rect 21135 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 14553 19703 14611 19709
rect 14553 19700 14565 19703
rect 13280 19672 14565 19700
rect 14553 19669 14565 19672
rect 14599 19700 14611 19703
rect 15746 19700 15752 19712
rect 14599 19672 15752 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 17218 19700 17224 19712
rect 16623 19672 17224 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 17494 19660 17500 19712
rect 17552 19700 17558 19712
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 17552 19672 18613 19700
rect 17552 19660 17558 19672
rect 18601 19669 18613 19672
rect 18647 19669 18659 19703
rect 19518 19700 19524 19712
rect 19479 19672 19524 19700
rect 18601 19663 18659 19669
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3605 19499 3663 19505
rect 3605 19496 3617 19499
rect 3108 19468 3617 19496
rect 3108 19456 3114 19468
rect 3605 19465 3617 19468
rect 3651 19465 3663 19499
rect 3605 19459 3663 19465
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4065 19499 4123 19505
rect 4065 19496 4077 19499
rect 4028 19468 4077 19496
rect 4028 19456 4034 19468
rect 4065 19465 4077 19468
rect 4111 19465 4123 19499
rect 4430 19496 4436 19508
rect 4391 19468 4436 19496
rect 4065 19459 4123 19465
rect 4430 19456 4436 19468
rect 4488 19496 4494 19508
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 4488 19468 4629 19496
rect 4488 19456 4494 19468
rect 4617 19465 4629 19468
rect 4663 19465 4675 19499
rect 6178 19496 6184 19508
rect 6139 19468 6184 19496
rect 4617 19459 4675 19465
rect 3513 19431 3571 19437
rect 3513 19397 3525 19431
rect 3559 19428 3571 19431
rect 3988 19428 4016 19456
rect 3559 19400 4016 19428
rect 3559 19397 3571 19400
rect 3513 19391 3571 19397
rect 3970 19360 3976 19372
rect 3931 19332 3976 19360
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 4632 19360 4660 19459
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 6730 19496 6736 19508
rect 6691 19468 6736 19496
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 7006 19456 7012 19508
rect 7064 19496 7070 19508
rect 7190 19496 7196 19508
rect 7064 19468 7196 19496
rect 7064 19456 7070 19468
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 9398 19496 9404 19508
rect 8996 19468 9404 19496
rect 8996 19456 9002 19468
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 9631 19468 9904 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 9876 19428 9904 19468
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 12618 19496 12624 19508
rect 10284 19468 12624 19496
rect 10284 19456 10290 19468
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 13262 19496 13268 19508
rect 12952 19468 13268 19496
rect 12952 19456 12958 19468
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13633 19499 13691 19505
rect 13633 19465 13645 19499
rect 13679 19496 13691 19499
rect 13722 19496 13728 19508
rect 13679 19468 13728 19496
rect 13679 19465 13691 19468
rect 13633 19459 13691 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19465 14795 19499
rect 14918 19496 14924 19508
rect 14879 19468 14924 19496
rect 14737 19459 14795 19465
rect 9950 19437 9956 19440
rect 9944 19428 9956 19437
rect 6972 19400 9720 19428
rect 9876 19400 9956 19428
rect 6972 19388 6978 19400
rect 4801 19363 4859 19369
rect 4801 19360 4813 19363
rect 4632 19332 4813 19360
rect 4801 19329 4813 19332
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 5068 19363 5126 19369
rect 5068 19329 5080 19363
rect 5114 19360 5126 19363
rect 5534 19360 5540 19372
rect 5114 19332 5540 19360
rect 5114 19329 5126 19332
rect 5068 19323 5126 19329
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 7374 19320 7380 19372
rect 7432 19360 7438 19372
rect 7857 19363 7915 19369
rect 7857 19360 7869 19363
rect 7432 19332 7869 19360
rect 7432 19320 7438 19332
rect 7857 19329 7869 19332
rect 7903 19360 7915 19363
rect 8018 19360 8024 19372
rect 7903 19332 8024 19360
rect 7903 19329 7915 19332
rect 7857 19323 7915 19329
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 8128 19369 8156 19400
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8202 19360 8208 19372
rect 8159 19332 8208 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8202 19320 8208 19332
rect 8260 19360 8266 19372
rect 8472 19363 8530 19369
rect 8260 19332 8353 19360
rect 8260 19320 8266 19332
rect 8472 19329 8484 19363
rect 8518 19360 8530 19363
rect 9582 19360 9588 19372
rect 8518 19332 9588 19360
rect 8518 19329 8530 19332
rect 8472 19323 8530 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 9692 19369 9720 19400
rect 9944 19391 9956 19400
rect 9950 19388 9956 19391
rect 10008 19388 10014 19440
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 14752 19428 14780 19459
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 15194 19456 15200 19508
rect 15252 19456 15258 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 16117 19499 16175 19505
rect 16117 19496 16129 19499
rect 15436 19468 16129 19496
rect 15436 19456 15442 19468
rect 16117 19465 16129 19468
rect 16163 19465 16175 19499
rect 16390 19496 16396 19508
rect 16351 19468 16396 19496
rect 16117 19459 16175 19465
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16942 19496 16948 19508
rect 16715 19468 16948 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17037 19499 17095 19505
rect 17037 19465 17049 19499
rect 17083 19496 17095 19499
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 17083 19468 17509 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 17497 19465 17509 19468
rect 17543 19465 17555 19499
rect 18877 19499 18935 19505
rect 18877 19496 18889 19499
rect 17497 19459 17555 19465
rect 17788 19468 18889 19496
rect 15212 19428 15240 19456
rect 12400 19400 13124 19428
rect 14752 19400 15240 19428
rect 12400 19388 12406 19400
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 12066 19360 12072 19372
rect 11296 19332 12072 19360
rect 11296 19320 11302 19332
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12641 19363 12699 19369
rect 12641 19329 12653 19363
rect 12687 19360 12699 19363
rect 12802 19360 12808 19372
rect 12687 19332 12808 19360
rect 12687 19329 12699 19332
rect 12641 19323 12699 19329
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4120 19264 4169 19292
rect 4120 19252 4126 19264
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 4157 19255 4215 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12943 19264 13001 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 13096 19292 13124 19400
rect 15654 19388 15660 19440
rect 15712 19428 15718 19440
rect 17129 19431 17187 19437
rect 15712 19400 17080 19428
rect 15712 19388 15718 19400
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13412 19332 13461 19360
rect 13412 19320 13418 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 13449 19323 13507 19329
rect 13740 19332 14289 19360
rect 13265 19295 13323 19301
rect 13265 19292 13277 19295
rect 13096 19264 13277 19292
rect 12989 19255 13047 19261
rect 13265 19261 13277 19264
rect 13311 19292 13323 19295
rect 13740 19292 13768 19332
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14366 19320 14372 19372
rect 14424 19360 14430 19372
rect 15102 19360 15108 19372
rect 14424 19332 14469 19360
rect 15063 19332 15108 19360
rect 14424 19320 14430 19332
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 15562 19360 15568 19372
rect 15523 19332 15568 19360
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 16301 19363 16359 19369
rect 15672 19332 16252 19360
rect 13311 19264 13768 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 11241 19227 11299 19233
rect 6104 19196 7236 19224
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 6104 19156 6132 19196
rect 6362 19156 6368 19168
rect 4672 19128 6132 19156
rect 6323 19128 6368 19156
rect 4672 19116 4678 19128
rect 6362 19116 6368 19128
rect 6420 19156 6426 19168
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6420 19128 6561 19156
rect 6420 19116 6426 19128
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 6914 19156 6920 19168
rect 6595 19128 6920 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7208 19156 7236 19196
rect 11241 19193 11253 19227
rect 11287 19224 11299 19227
rect 11287 19196 11836 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 10962 19156 10968 19168
rect 7208 19128 10968 19156
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11057 19159 11115 19165
rect 11057 19125 11069 19159
rect 11103 19156 11115 19159
rect 11146 19156 11152 19168
rect 11103 19128 11152 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11517 19159 11575 19165
rect 11517 19125 11529 19159
rect 11563 19156 11575 19159
rect 11698 19156 11704 19168
rect 11563 19128 11704 19156
rect 11563 19125 11575 19128
rect 11517 19119 11575 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11808 19156 11836 19196
rect 12526 19156 12532 19168
rect 11808 19128 12532 19156
rect 12526 19116 12532 19128
rect 12584 19156 12590 19168
rect 12912 19156 12940 19255
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 15672 19301 15700 19332
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13872 19264 14105 19292
rect 13872 19252 13878 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 16224 19292 16252 19332
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 16942 19360 16948 19372
rect 16347 19332 16948 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17052 19360 17080 19400
rect 17129 19397 17141 19431
rect 17175 19428 17187 19431
rect 17218 19428 17224 19440
rect 17175 19400 17224 19428
rect 17175 19397 17187 19400
rect 17129 19391 17187 19397
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 17788 19360 17816 19468
rect 18877 19465 18889 19468
rect 18923 19465 18935 19499
rect 18877 19459 18935 19465
rect 20993 19499 21051 19505
rect 20993 19465 21005 19499
rect 21039 19496 21051 19499
rect 21082 19496 21088 19508
rect 21039 19468 21088 19496
rect 21039 19465 21051 19468
rect 20993 19459 21051 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 17865 19431 17923 19437
rect 17865 19397 17877 19431
rect 17911 19428 17923 19431
rect 17954 19428 17960 19440
rect 17911 19400 17960 19428
rect 17911 19397 17923 19400
rect 17865 19391 17923 19397
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18230 19428 18236 19440
rect 18064 19400 18236 19428
rect 17052 19332 17816 19360
rect 16390 19292 16396 19304
rect 15804 19264 15849 19292
rect 16224 19264 16396 19292
rect 15804 19252 15810 19264
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 17218 19292 17224 19304
rect 17179 19264 17224 19292
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 18064 19301 18092 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 18322 19360 18328 19372
rect 18283 19332 18328 19360
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18656 19332 18705 19360
rect 18656 19320 18662 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17736 19264 17969 19292
rect 17736 19252 17742 19264
rect 17957 19261 17969 19264
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 13170 19184 13176 19236
rect 13228 19224 13234 19236
rect 13228 19196 15608 19224
rect 13228 19184 13234 19196
rect 13814 19156 13820 19168
rect 12584 19128 12940 19156
rect 13775 19128 13820 19156
rect 12584 19116 12590 19128
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 15197 19159 15255 19165
rect 15197 19125 15209 19159
rect 15243 19156 15255 19159
rect 15470 19156 15476 19168
rect 15243 19128 15476 19156
rect 15243 19125 15255 19128
rect 15197 19119 15255 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15580 19156 15608 19196
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 18509 19227 18567 19233
rect 18509 19224 18521 19227
rect 17368 19196 18521 19224
rect 17368 19184 17374 19196
rect 18509 19193 18521 19196
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 18966 19156 18972 19168
rect 15580 19128 18972 19156
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 20714 19156 20720 19168
rect 20627 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19156 20778 19168
rect 20824 19156 20852 19323
rect 22370 19156 22376 19168
rect 20772 19128 22376 19156
rect 20772 19116 20778 19128
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 4430 18952 4436 18964
rect 4391 18924 4436 18952
rect 4430 18912 4436 18924
rect 4488 18912 4494 18964
rect 4617 18955 4675 18961
rect 4617 18921 4629 18955
rect 4663 18952 4675 18955
rect 4982 18952 4988 18964
rect 4663 18924 4988 18952
rect 4663 18921 4675 18924
rect 4617 18915 4675 18921
rect 4982 18912 4988 18924
rect 5040 18952 5046 18964
rect 6546 18952 6552 18964
rect 5040 18924 6552 18952
rect 5040 18912 5046 18924
rect 6546 18912 6552 18924
rect 6604 18952 6610 18964
rect 7006 18952 7012 18964
rect 6604 18924 7012 18952
rect 6604 18912 6610 18924
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7285 18955 7343 18961
rect 7285 18921 7297 18955
rect 7331 18952 7343 18955
rect 9306 18952 9312 18964
rect 7331 18924 9312 18952
rect 7331 18921 7343 18924
rect 7285 18915 7343 18921
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 9582 18912 9588 18964
rect 9640 18952 9646 18964
rect 10965 18955 11023 18961
rect 9640 18924 10640 18952
rect 9640 18912 9646 18924
rect 4448 18816 4476 18912
rect 7374 18884 7380 18896
rect 7335 18856 7380 18884
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 9033 18887 9091 18893
rect 9033 18853 9045 18887
rect 9079 18884 9091 18887
rect 9214 18884 9220 18896
rect 9079 18856 9220 18884
rect 9079 18853 9091 18856
rect 9033 18847 9091 18853
rect 9214 18844 9220 18856
rect 9272 18844 9278 18896
rect 10612 18884 10640 18924
rect 10965 18921 10977 18955
rect 11011 18952 11023 18955
rect 12434 18952 12440 18964
rect 11011 18924 12440 18952
rect 11011 18921 11023 18924
rect 10965 18915 11023 18921
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 12676 18924 13829 18952
rect 12676 18912 12682 18924
rect 13817 18921 13829 18924
rect 13863 18952 13875 18955
rect 14366 18952 14372 18964
rect 13863 18924 14372 18952
rect 13863 18921 13875 18924
rect 13817 18915 13875 18921
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 17034 18952 17040 18964
rect 16995 18924 17040 18952
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 20622 18912 20628 18964
rect 20680 18952 20686 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 20680 18924 21005 18952
rect 20680 18912 20686 18924
rect 20993 18921 21005 18924
rect 21039 18921 21051 18955
rect 20993 18915 21051 18921
rect 11054 18884 11060 18896
rect 10612 18856 11060 18884
rect 11054 18844 11060 18856
rect 11112 18844 11118 18896
rect 12452 18884 12480 18912
rect 12802 18884 12808 18896
rect 12452 18856 12808 18884
rect 12802 18844 12808 18856
rect 12860 18844 12866 18896
rect 15841 18887 15899 18893
rect 15841 18853 15853 18887
rect 15887 18884 15899 18887
rect 15887 18856 17264 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4448 18788 4721 18816
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7190 18816 7196 18828
rect 6779 18788 7196 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 4724 18748 4752 18779
rect 7190 18776 7196 18788
rect 7248 18816 7254 18828
rect 7558 18816 7564 18828
rect 7248 18788 7564 18816
rect 7248 18776 7254 18788
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 8938 18776 8944 18828
rect 8996 18816 9002 18828
rect 12437 18819 12495 18825
rect 8996 18788 9720 18816
rect 8996 18776 9002 18788
rect 5994 18748 6000 18760
rect 4724 18720 6000 18748
rect 5994 18708 6000 18720
rect 6052 18748 6058 18760
rect 6181 18751 6239 18757
rect 6181 18748 6193 18751
rect 6052 18720 6193 18748
rect 6052 18708 6058 18720
rect 6181 18717 6193 18720
rect 6227 18748 6239 18751
rect 6362 18748 6368 18760
rect 6227 18720 6368 18748
rect 6227 18717 6239 18720
rect 6181 18711 6239 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 7098 18748 7104 18760
rect 6871 18720 7104 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8757 18751 8815 18757
rect 8757 18748 8769 18751
rect 8260 18720 8769 18748
rect 8260 18708 8266 18720
rect 8757 18717 8769 18720
rect 8803 18748 8815 18751
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 8803 18720 9413 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9401 18717 9413 18720
rect 9447 18748 9459 18751
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9447 18720 9597 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9692 18748 9720 18788
rect 12437 18785 12449 18819
rect 12483 18816 12495 18819
rect 12526 18816 12532 18828
rect 12483 18788 12532 18816
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 15194 18816 15200 18828
rect 15155 18788 15200 18816
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 15804 18788 16589 18816
rect 15804 18776 15810 18788
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 9692 18720 10180 18748
rect 9585 18711 9643 18717
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 4982 18689 4988 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 4028 18652 4077 18680
rect 4028 18640 4034 18652
rect 4065 18649 4077 18652
rect 4111 18680 4123 18683
rect 4111 18652 4936 18680
rect 4111 18649 4123 18652
rect 4065 18643 4123 18649
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 4908 18612 4936 18652
rect 4976 18643 4988 18689
rect 5040 18680 5046 18692
rect 8386 18680 8392 18692
rect 5040 18652 5076 18680
rect 5460 18652 8392 18680
rect 4982 18640 4988 18643
rect 5040 18640 5046 18652
rect 5460 18612 5488 18652
rect 8386 18640 8392 18652
rect 8444 18640 8450 18692
rect 9858 18689 9864 18692
rect 8512 18683 8570 18689
rect 8512 18649 8524 18683
rect 8558 18680 8570 18683
rect 8558 18652 9812 18680
rect 8558 18649 8570 18652
rect 8512 18643 8570 18649
rect 4908 18584 5488 18612
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 6089 18615 6147 18621
rect 6089 18612 6101 18615
rect 5592 18584 6101 18612
rect 5592 18572 5598 18584
rect 6089 18581 6101 18584
rect 6135 18612 6147 18615
rect 6546 18612 6552 18624
rect 6135 18584 6552 18612
rect 6135 18581 6147 18584
rect 6089 18575 6147 18581
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7374 18612 7380 18624
rect 6963 18584 7380 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 7926 18572 7932 18624
rect 7984 18612 7990 18624
rect 8938 18612 8944 18624
rect 7984 18584 8944 18612
rect 7984 18572 7990 18584
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 9088 18584 9137 18612
rect 9088 18572 9094 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9674 18612 9680 18624
rect 9364 18584 9680 18612
rect 9364 18572 9370 18584
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 9784 18612 9812 18652
rect 9852 18643 9864 18689
rect 9916 18680 9922 18692
rect 9916 18652 9952 18680
rect 9858 18640 9864 18643
rect 9916 18640 9922 18652
rect 9950 18612 9956 18624
rect 9784 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10152 18612 10180 18720
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 10928 18720 11652 18748
rect 10928 18708 10934 18720
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11146 18680 11152 18692
rect 10560 18652 11152 18680
rect 10560 18640 10566 18652
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 11624 18680 11652 18720
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12158 18748 12164 18760
rect 12216 18757 12222 18760
rect 11756 18720 12164 18748
rect 11756 18708 11762 18720
rect 12158 18708 12164 18720
rect 12216 18711 12228 18757
rect 15470 18748 15476 18760
rect 12912 18720 15240 18748
rect 15431 18720 15476 18748
rect 12216 18708 12222 18711
rect 12912 18680 12940 18720
rect 15212 18692 15240 18720
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 17236 18757 17264 18856
rect 17678 18844 17684 18896
rect 17736 18884 17742 18896
rect 20714 18884 20720 18896
rect 17736 18856 20720 18884
rect 17736 18844 17742 18856
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 17954 18816 17960 18828
rect 17915 18788 17960 18816
rect 17954 18776 17960 18788
rect 18012 18776 18018 18828
rect 18414 18816 18420 18828
rect 18375 18788 18420 18816
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16264 18720 16865 18748
rect 16264 18708 16270 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 17221 18711 17279 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 20809 18751 20867 18757
rect 20809 18717 20821 18751
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 11624 18652 12940 18680
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 13035 18652 13553 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 13541 18649 13553 18652
rect 13587 18680 13599 18683
rect 13722 18680 13728 18692
rect 13587 18652 13728 18680
rect 13587 18649 13599 18652
rect 13541 18643 13599 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 15194 18640 15200 18692
rect 15252 18640 15258 18692
rect 15381 18683 15439 18689
rect 15381 18649 15393 18683
rect 15427 18680 15439 18683
rect 16390 18680 16396 18692
rect 15427 18652 16068 18680
rect 16351 18652 16396 18680
rect 15427 18649 15439 18652
rect 15381 18643 15439 18649
rect 11882 18612 11888 18624
rect 10152 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 12710 18612 12716 18624
rect 12667 18584 12716 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12860 18584 13093 18612
rect 12860 18572 12866 18584
rect 13081 18581 13093 18584
rect 13127 18612 13139 18615
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13127 18584 13645 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13633 18581 13645 18584
rect 13679 18612 13691 18615
rect 15654 18612 15660 18624
rect 13679 18584 15660 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 16040 18621 16068 18652
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 17497 18683 17555 18689
rect 17497 18649 17509 18683
rect 17543 18680 17555 18683
rect 18782 18680 18788 18692
rect 17543 18652 18788 18680
rect 17543 18649 17555 18652
rect 17497 18643 17555 18649
rect 18782 18640 18788 18652
rect 18840 18640 18846 18692
rect 16025 18615 16083 18621
rect 16025 18581 16037 18615
rect 16071 18581 16083 18615
rect 16025 18575 16083 18581
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 16485 18615 16543 18621
rect 16485 18612 16497 18615
rect 16356 18584 16497 18612
rect 16356 18572 16362 18584
rect 16485 18581 16497 18584
rect 16531 18581 16543 18615
rect 16485 18575 16543 18581
rect 20717 18615 20775 18621
rect 20717 18581 20729 18615
rect 20763 18612 20775 18615
rect 20824 18612 20852 18711
rect 21082 18612 21088 18624
rect 20763 18584 21088 18612
rect 20763 18581 20775 18584
rect 20717 18575 20775 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 2774 18408 2780 18420
rect 1995 18380 2780 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6822 18408 6828 18420
rect 6236 18380 6828 18408
rect 6236 18368 6242 18380
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 12342 18408 12348 18420
rect 7708 18380 12348 18408
rect 7708 18368 7714 18380
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12618 18408 12624 18420
rect 12575 18380 12624 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12618 18368 12624 18380
rect 12676 18408 12682 18420
rect 13170 18408 13176 18420
rect 12676 18380 13176 18408
rect 12676 18368 12682 18380
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 14056 18380 14289 18408
rect 14056 18368 14062 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14737 18411 14795 18417
rect 14737 18377 14749 18411
rect 14783 18408 14795 18411
rect 15562 18408 15568 18420
rect 14783 18380 15424 18408
rect 15523 18380 15568 18408
rect 14783 18377 14795 18380
rect 14737 18371 14795 18377
rect 5534 18300 5540 18352
rect 5592 18349 5598 18352
rect 5592 18340 5604 18349
rect 5592 18312 5637 18340
rect 5592 18303 5604 18312
rect 5592 18300 5598 18303
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2406 18272 2412 18284
rect 2179 18244 2412 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 5813 18275 5871 18281
rect 4304 18244 5764 18272
rect 4304 18232 4310 18244
rect 5736 18204 5764 18244
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6012 18272 6040 18368
rect 7282 18340 7288 18352
rect 6380 18312 7288 18340
rect 6380 18281 6408 18312
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 9401 18343 9459 18349
rect 9401 18340 9413 18343
rect 7944 18312 9413 18340
rect 6638 18281 6644 18284
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5859 18244 6377 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6632 18272 6644 18281
rect 6599 18244 6644 18272
rect 6365 18235 6423 18241
rect 6632 18235 6644 18244
rect 6638 18232 6644 18235
rect 6696 18232 6702 18284
rect 7300 18272 7328 18300
rect 7944 18281 7972 18312
rect 9401 18309 9413 18312
rect 9447 18340 9459 18343
rect 9769 18343 9827 18349
rect 9769 18340 9781 18343
rect 9447 18312 9781 18340
rect 9447 18309 9459 18312
rect 9401 18303 9459 18309
rect 9769 18309 9781 18312
rect 9815 18340 9827 18343
rect 9815 18312 11376 18340
rect 9815 18309 9827 18312
rect 9769 18303 9827 18309
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 7300 18244 7941 18272
rect 7929 18241 7941 18244
rect 7975 18241 7987 18275
rect 7929 18235 7987 18241
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8196 18275 8254 18281
rect 8196 18272 8208 18275
rect 8076 18244 8208 18272
rect 8076 18232 8082 18244
rect 8196 18241 8208 18244
rect 8242 18241 8254 18275
rect 8196 18235 8254 18241
rect 11077 18275 11135 18281
rect 11077 18241 11089 18275
rect 11123 18272 11135 18275
rect 11238 18272 11244 18284
rect 11123 18244 11244 18272
rect 11123 18241 11135 18244
rect 11077 18235 11135 18241
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 11348 18281 11376 18312
rect 12158 18300 12164 18352
rect 12216 18340 12222 18352
rect 12216 18312 12664 18340
rect 12216 18300 12222 18312
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 12526 18272 12532 18284
rect 11379 18244 12532 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 12636 18272 12664 18312
rect 12802 18300 12808 18352
rect 12860 18340 12866 18352
rect 13354 18340 13360 18352
rect 12860 18312 13360 18340
rect 12860 18300 12866 18312
rect 13354 18300 13360 18312
rect 13412 18300 13418 18352
rect 13630 18340 13636 18352
rect 13591 18312 13636 18340
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 15102 18340 15108 18352
rect 13740 18312 14504 18340
rect 15063 18312 15108 18340
rect 13740 18272 13768 18312
rect 12636 18244 13768 18272
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14182 18272 14188 18284
rect 13955 18244 14188 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 10226 18204 10232 18216
rect 5736 18176 6316 18204
rect 2317 18139 2375 18145
rect 2317 18105 2329 18139
rect 2363 18136 2375 18139
rect 2498 18136 2504 18148
rect 2363 18108 2504 18136
rect 2363 18105 2375 18108
rect 2317 18099 2375 18105
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 2406 18068 2412 18080
rect 2367 18040 2412 18068
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 4706 18068 4712 18080
rect 4479 18040 4712 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4706 18028 4712 18040
rect 4764 18068 4770 18080
rect 6178 18068 6184 18080
rect 4764 18040 6184 18068
rect 4764 18028 4770 18040
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6288 18068 6316 18176
rect 8956 18176 10232 18204
rect 7374 18068 7380 18080
rect 6288 18040 7380 18068
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 7745 18071 7803 18077
rect 7745 18068 7757 18071
rect 7708 18040 7757 18068
rect 7708 18028 7714 18040
rect 7745 18037 7757 18040
rect 7791 18037 7803 18071
rect 7745 18031 7803 18037
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8956 18068 8984 18176
rect 10226 18164 10232 18176
rect 10284 18164 10290 18216
rect 13722 18204 13728 18216
rect 11348 18176 13728 18204
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 9858 18136 9864 18148
rect 9355 18108 9864 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 9858 18096 9864 18108
rect 9916 18136 9922 18148
rect 10318 18136 10324 18148
rect 9916 18108 10324 18136
rect 9916 18096 9922 18108
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 9950 18068 9956 18080
rect 7892 18040 8984 18068
rect 9911 18040 9956 18068
rect 7892 18028 7898 18040
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 11348 18068 11376 18176
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 11698 18096 11704 18148
rect 11756 18136 11762 18148
rect 14108 18136 14136 18167
rect 11756 18108 14136 18136
rect 14476 18136 14504 18312
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 15396 18340 15424 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16448 18380 16865 18408
rect 16448 18368 16454 18380
rect 16853 18377 16865 18380
rect 16899 18377 16911 18411
rect 16853 18371 16911 18377
rect 20530 18368 20536 18420
rect 20588 18408 20594 18420
rect 20993 18411 21051 18417
rect 20993 18408 21005 18411
rect 20588 18380 21005 18408
rect 20588 18368 20594 18380
rect 20993 18377 21005 18380
rect 21039 18377 21051 18411
rect 20993 18371 21051 18377
rect 17405 18343 17463 18349
rect 15396 18312 17356 18340
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 17126 18272 17132 18284
rect 17087 18244 17132 18272
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17328 18272 17356 18312
rect 17405 18309 17417 18343
rect 17451 18340 17463 18343
rect 18322 18340 18328 18352
rect 17451 18312 18328 18340
rect 17451 18309 17463 18312
rect 17405 18303 17463 18309
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 19058 18272 19064 18284
rect 17328 18244 19064 18272
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20772 18244 20821 18272
rect 20772 18232 20778 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 15102 18204 15108 18216
rect 14700 18176 15108 18204
rect 14700 18164 14706 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15804 18176 15853 18204
rect 15804 18164 15810 18176
rect 15841 18173 15853 18176
rect 15887 18204 15899 18207
rect 16298 18204 16304 18216
rect 15887 18176 16304 18204
rect 15887 18173 15899 18176
rect 15841 18167 15899 18173
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 17681 18207 17739 18213
rect 17681 18204 17693 18207
rect 17460 18176 17693 18204
rect 17460 18164 17466 18176
rect 17681 18173 17693 18176
rect 17727 18173 17739 18207
rect 17681 18167 17739 18173
rect 17310 18136 17316 18148
rect 14476 18108 17316 18136
rect 11756 18096 11762 18108
rect 10100 18040 11376 18068
rect 10100 18028 10106 18040
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12986 18068 12992 18080
rect 11940 18040 12992 18068
rect 11940 18028 11946 18040
rect 12986 18028 12992 18040
rect 13044 18068 13050 18080
rect 13265 18071 13323 18077
rect 13265 18068 13277 18071
rect 13044 18040 13277 18068
rect 13044 18028 13050 18040
rect 13265 18037 13277 18040
rect 13311 18068 13323 18071
rect 13998 18068 14004 18080
rect 13311 18040 14004 18068
rect 13311 18037 13323 18040
rect 13265 18031 13323 18037
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 14108 18068 14136 18108
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 17218 18068 17224 18080
rect 14108 18040 17224 18068
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 19153 18071 19211 18077
rect 19153 18037 19165 18071
rect 19199 18068 19211 18071
rect 19702 18068 19708 18080
rect 19199 18040 19708 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1949 17867 2007 17873
rect 1949 17833 1961 17867
rect 1995 17864 2007 17867
rect 2866 17864 2872 17876
rect 1995 17836 2872 17864
rect 1995 17833 2007 17836
rect 1949 17827 2007 17833
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 5905 17867 5963 17873
rect 3375 17836 5764 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 2590 17756 2596 17808
rect 2648 17796 2654 17808
rect 3344 17796 3372 17827
rect 2648 17768 3372 17796
rect 2648 17756 2654 17768
rect 2409 17731 2467 17737
rect 2409 17697 2421 17731
rect 2455 17728 2467 17731
rect 4062 17728 4068 17740
rect 2455 17700 4068 17728
rect 2455 17697 2467 17700
rect 2409 17691 2467 17697
rect 4062 17688 4068 17700
rect 4120 17728 4126 17740
rect 4430 17728 4436 17740
rect 4120 17700 4292 17728
rect 4391 17700 4436 17728
rect 4120 17688 4126 17700
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2498 17660 2504 17672
rect 2179 17632 2504 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17660 2651 17663
rect 2639 17632 2774 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 2746 17592 2774 17632
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 2746 17564 3065 17592
rect 3053 17561 3065 17564
rect 3099 17592 3111 17595
rect 4264 17592 4292 17700
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 5736 17728 5764 17836
rect 5905 17833 5917 17867
rect 5951 17864 5963 17867
rect 6362 17864 6368 17876
rect 5951 17836 6368 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 6638 17824 6644 17876
rect 6696 17864 6702 17876
rect 9858 17864 9864 17876
rect 6696 17836 9864 17864
rect 6696 17824 6702 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 12894 17864 12900 17876
rect 10060 17836 12900 17864
rect 5813 17799 5871 17805
rect 5813 17765 5825 17799
rect 5859 17796 5871 17799
rect 5859 17768 6316 17796
rect 5859 17765 5871 17768
rect 5813 17759 5871 17765
rect 5736 17700 6224 17728
rect 4706 17669 4712 17672
rect 4700 17660 4712 17669
rect 4667 17632 4712 17660
rect 4700 17623 4712 17632
rect 4706 17620 4712 17623
rect 4764 17620 4770 17672
rect 4982 17592 4988 17604
rect 3099 17564 3372 17592
rect 4264 17564 4988 17592
rect 3099 17561 3111 17564
rect 3053 17555 3111 17561
rect 3344 17536 3372 17564
rect 4982 17552 4988 17564
rect 5040 17552 5046 17604
rect 6196 17592 6224 17700
rect 6288 17660 6316 17768
rect 7282 17728 7288 17740
rect 7243 17700 7288 17728
rect 7282 17688 7288 17700
rect 7340 17728 7346 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7340 17700 7389 17728
rect 7340 17688 7346 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 10060 17728 10088 17836
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 13909 17867 13967 17873
rect 13004 17836 13860 17864
rect 11054 17756 11060 17808
rect 11112 17796 11118 17808
rect 13004 17796 13032 17836
rect 11112 17768 13032 17796
rect 13832 17796 13860 17836
rect 13909 17833 13921 17867
rect 13955 17864 13967 17867
rect 13998 17864 14004 17876
rect 13955 17836 14004 17864
rect 13955 17833 13967 17836
rect 13909 17827 13967 17833
rect 13998 17824 14004 17836
rect 14056 17864 14062 17876
rect 14366 17864 14372 17876
rect 14056 17836 14372 17864
rect 14056 17824 14062 17836
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 14921 17867 14979 17873
rect 14921 17864 14933 17867
rect 14884 17836 14933 17864
rect 14884 17824 14890 17836
rect 14921 17833 14933 17836
rect 14967 17833 14979 17867
rect 14921 17827 14979 17833
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 16025 17867 16083 17873
rect 16025 17864 16037 17867
rect 15252 17836 16037 17864
rect 15252 17824 15258 17836
rect 16025 17833 16037 17836
rect 16071 17864 16083 17867
rect 16482 17864 16488 17876
rect 16071 17836 16488 17864
rect 16071 17833 16083 17836
rect 16025 17827 16083 17833
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 17184 17836 17233 17864
rect 17184 17824 17190 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 20257 17867 20315 17873
rect 18288 17836 18333 17864
rect 18288 17824 18294 17836
rect 20257 17833 20269 17867
rect 20303 17864 20315 17867
rect 20622 17864 20628 17876
rect 20303 17836 20628 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 17034 17796 17040 17808
rect 13832 17768 17040 17796
rect 11112 17756 11118 17768
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 19886 17796 19892 17808
rect 17144 17768 19892 17796
rect 10060 17700 10180 17728
rect 7377 17691 7435 17697
rect 7392 17660 7420 17691
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 6288 17632 7328 17660
rect 7392 17632 8953 17660
rect 6730 17592 6736 17604
rect 5092 17564 6040 17592
rect 6196 17564 6736 17592
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 2590 17524 2596 17536
rect 2547 17496 2596 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 2958 17524 2964 17536
rect 2919 17496 2964 17524
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 3326 17484 3332 17536
rect 3384 17524 3390 17536
rect 5092 17524 5120 17564
rect 3384 17496 5120 17524
rect 6012 17524 6040 17564
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 7018 17595 7076 17601
rect 7018 17592 7030 17595
rect 6880 17564 7030 17592
rect 6880 17552 6886 17564
rect 7018 17561 7030 17564
rect 7064 17561 7076 17595
rect 7300 17592 7328 17632
rect 8941 17629 8953 17632
rect 8987 17660 8999 17663
rect 9766 17660 9772 17672
rect 8987 17632 9772 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9766 17620 9772 17632
rect 9824 17660 9830 17672
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9824 17632 9873 17660
rect 9824 17620 9830 17632
rect 9861 17629 9873 17632
rect 9907 17660 9919 17663
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9907 17632 10057 17660
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 10045 17629 10057 17632
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 7644 17595 7702 17601
rect 7644 17592 7656 17595
rect 7300 17564 7656 17592
rect 7018 17555 7076 17561
rect 7644 17561 7656 17564
rect 7690 17592 7702 17595
rect 10152 17592 10180 17700
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13538 17728 13544 17740
rect 13412 17700 13457 17728
rect 13499 17700 13544 17728
rect 13412 17688 13418 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 14642 17728 14648 17740
rect 14603 17700 14648 17728
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 10312 17663 10370 17669
rect 10312 17629 10324 17663
rect 10358 17660 10370 17663
rect 15488 17660 15516 17691
rect 16114 17688 16120 17740
rect 16172 17728 16178 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 16172 17700 16221 17728
rect 16172 17688 16178 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16482 17728 16488 17740
rect 16443 17700 16488 17728
rect 16209 17691 16267 17697
rect 10358 17632 13308 17660
rect 10358 17629 10370 17632
rect 10312 17623 10370 17629
rect 7690 17564 10180 17592
rect 7690 17561 7702 17564
rect 7644 17555 7702 17561
rect 8294 17524 8300 17536
rect 6012 17496 8300 17524
rect 3384 17484 3390 17496
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8757 17527 8815 17533
rect 8757 17493 8769 17527
rect 8803 17524 8815 17527
rect 10327 17524 10355 17623
rect 10686 17552 10692 17604
rect 10744 17592 10750 17604
rect 11974 17592 11980 17604
rect 10744 17564 11980 17592
rect 10744 17552 10750 17564
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 13170 17552 13176 17604
rect 13228 17552 13234 17604
rect 13280 17592 13308 17632
rect 13464 17632 15516 17660
rect 13464 17592 13492 17632
rect 13280 17564 13492 17592
rect 16224 17592 16252 17691
rect 16482 17688 16488 17700
rect 16540 17728 16546 17740
rect 17144 17728 17172 17768
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 17770 17728 17776 17740
rect 16540 17700 17172 17728
rect 17731 17700 17776 17728
rect 16540 17688 16546 17700
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 18782 17728 18788 17740
rect 18743 17700 18788 17728
rect 18782 17688 18788 17700
rect 18840 17688 18846 17740
rect 19794 17728 19800 17740
rect 19755 17700 19800 17728
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 16666 17660 16672 17672
rect 16627 17632 16672 17660
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 20073 17663 20131 17669
rect 20073 17660 20085 17663
rect 16868 17632 20085 17660
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 16224 17564 16773 17592
rect 16761 17561 16773 17564
rect 16807 17561 16819 17595
rect 16761 17555 16819 17561
rect 8803 17496 10355 17524
rect 8803 17493 8815 17496
rect 8757 17487 8815 17493
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11296 17496 11437 17524
rect 11296 17484 11302 17496
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 12897 17527 12955 17533
rect 12897 17493 12909 17527
rect 12943 17524 12955 17527
rect 13188 17524 13216 17552
rect 12943 17496 13216 17524
rect 13265 17527 13323 17533
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13265 17493 13277 17527
rect 13311 17524 13323 17527
rect 13814 17524 13820 17536
rect 13311 17496 13820 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 14090 17524 14096 17536
rect 14051 17496 14096 17524
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14458 17524 14464 17536
rect 14419 17496 14464 17524
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 14826 17524 14832 17536
rect 14599 17496 14832 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 15010 17484 15016 17536
rect 15068 17524 15074 17536
rect 15289 17527 15347 17533
rect 15289 17524 15301 17527
rect 15068 17496 15301 17524
rect 15068 17484 15074 17496
rect 15289 17493 15301 17496
rect 15335 17493 15347 17527
rect 15289 17487 15347 17493
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16868 17524 16896 17632
rect 20073 17629 20085 17632
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 18414 17592 18420 17604
rect 17144 17564 18420 17592
rect 17144 17533 17172 17564
rect 18414 17552 18420 17564
rect 18472 17552 18478 17604
rect 18601 17595 18659 17601
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 18647 17564 19288 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 16172 17496 16896 17524
rect 17129 17527 17187 17533
rect 16172 17484 16178 17496
rect 17129 17493 17141 17527
rect 17175 17493 17187 17527
rect 17586 17524 17592 17536
rect 17547 17496 17592 17524
rect 17129 17487 17187 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 17681 17527 17739 17533
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 18322 17524 18328 17536
rect 17727 17496 18328 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 19150 17524 19156 17536
rect 18739 17496 19156 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 19150 17484 19156 17496
rect 19208 17484 19214 17536
rect 19260 17533 19288 17564
rect 19245 17527 19303 17533
rect 19245 17493 19257 17527
rect 19291 17493 19303 17527
rect 19610 17524 19616 17536
rect 19571 17496 19616 17524
rect 19245 17487 19303 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 21174 17524 21180 17536
rect 19760 17496 21180 17524
rect 19760 17484 19766 17496
rect 21174 17484 21180 17496
rect 21232 17524 21238 17536
rect 22462 17524 22468 17536
rect 21232 17496 22468 17524
rect 21232 17484 21238 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 2774 17320 2780 17332
rect 2731 17292 2780 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3053 17323 3111 17329
rect 3053 17289 3065 17323
rect 3099 17320 3111 17323
rect 3326 17320 3332 17332
rect 3099 17292 3332 17320
rect 3099 17289 3111 17292
rect 3053 17283 3111 17289
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 6457 17323 6515 17329
rect 6457 17289 6469 17323
rect 6503 17320 6515 17323
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6503 17292 6653 17320
rect 6503 17289 6515 17292
rect 6457 17283 6515 17289
rect 6641 17289 6653 17292
rect 6687 17320 6699 17323
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6687 17292 6837 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 6825 17289 6837 17292
rect 6871 17320 6883 17323
rect 7193 17323 7251 17329
rect 7193 17320 7205 17323
rect 6871 17292 7205 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7193 17289 7205 17292
rect 7239 17320 7251 17323
rect 7282 17320 7288 17332
rect 7239 17292 7288 17320
rect 7239 17289 7251 17292
rect 7193 17283 7251 17289
rect 3237 17255 3295 17261
rect 3237 17252 3249 17255
rect 2746 17224 3249 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1811 17156 2145 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2133 17153 2145 17156
rect 2179 17184 2191 17187
rect 2222 17184 2228 17196
rect 2179 17156 2228 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2516 17116 2544 17147
rect 2746 17116 2774 17224
rect 3237 17221 3249 17224
rect 3283 17252 3295 17255
rect 3283 17224 6132 17252
rect 3283 17221 3295 17224
rect 3237 17215 3295 17221
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17184 2927 17187
rect 3326 17184 3332 17196
rect 2915 17156 3332 17184
rect 2915 17153 2927 17156
rect 2869 17147 2927 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 5626 17184 5632 17196
rect 4304 17156 5632 17184
rect 4304 17144 4310 17156
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 5902 17144 5908 17196
rect 5960 17193 5966 17196
rect 5960 17184 5972 17193
rect 5960 17156 6005 17184
rect 5960 17147 5972 17156
rect 5960 17144 5966 17147
rect 2516 17088 2774 17116
rect 6104 17116 6132 17224
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 6270 17184 6276 17196
rect 6227 17156 6276 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6270 17144 6276 17156
rect 6328 17184 6334 17196
rect 6472 17184 6500 17283
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 9214 17320 9220 17332
rect 7432 17292 9220 17320
rect 7432 17280 7438 17292
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9766 17320 9772 17332
rect 9727 17292 9772 17320
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 9916 17292 10180 17320
rect 9916 17280 9922 17292
rect 7300 17193 7328 17280
rect 10042 17252 10048 17264
rect 7392 17224 10048 17252
rect 6328 17156 6500 17184
rect 7285 17187 7343 17193
rect 6328 17144 6334 17156
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7392 17116 7420 17224
rect 10042 17212 10048 17224
rect 10100 17212 10106 17264
rect 10152 17252 10180 17292
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10870 17320 10876 17332
rect 10284 17292 10876 17320
rect 10284 17280 10290 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 12805 17323 12863 17329
rect 12805 17320 12817 17323
rect 11204 17292 12817 17320
rect 11204 17280 11210 17292
rect 12805 17289 12817 17292
rect 12851 17320 12863 17323
rect 13998 17320 14004 17332
rect 12851 17292 14004 17320
rect 12851 17289 12863 17292
rect 12805 17283 12863 17289
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 17313 17323 17371 17329
rect 17313 17289 17325 17323
rect 17359 17320 17371 17323
rect 17402 17320 17408 17332
rect 17359 17292 17408 17320
rect 17359 17289 17371 17292
rect 17313 17283 17371 17289
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17681 17323 17739 17329
rect 17681 17320 17693 17323
rect 17644 17292 17693 17320
rect 17644 17280 17650 17292
rect 17681 17289 17693 17292
rect 17727 17289 17739 17323
rect 18322 17320 18328 17332
rect 18283 17292 18328 17320
rect 17681 17283 17739 17289
rect 18322 17280 18328 17292
rect 18380 17280 18386 17332
rect 19150 17320 19156 17332
rect 19111 17292 19156 17320
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 19981 17323 20039 17329
rect 19981 17320 19993 17323
rect 19668 17292 19993 17320
rect 19668 17280 19674 17292
rect 19981 17289 19993 17292
rect 20027 17289 20039 17323
rect 19981 17283 20039 17289
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20496 17292 21005 17320
rect 20496 17280 20502 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 20993 17283 21051 17289
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 11882 17252 11888 17264
rect 10152 17224 11888 17252
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12986 17252 12992 17264
rect 12947 17224 12992 17252
rect 12986 17212 12992 17224
rect 13044 17212 13050 17264
rect 13262 17252 13268 17264
rect 13096 17224 13268 17252
rect 7552 17187 7610 17193
rect 7552 17153 7564 17187
rect 7598 17184 7610 17187
rect 7834 17184 7840 17196
rect 7598 17156 7840 17184
rect 7598 17153 7610 17156
rect 7552 17147 7610 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8662 17184 8668 17196
rect 8076 17156 8668 17184
rect 8076 17144 8082 17156
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9824 17156 9965 17184
rect 9824 17144 9830 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10220 17187 10278 17193
rect 10220 17153 10232 17187
rect 10266 17184 10278 17187
rect 11698 17184 11704 17196
rect 10266 17156 11704 17184
rect 10266 17153 10278 17156
rect 10220 17147 10278 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13096 17193 13124 17224
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 14737 17255 14795 17261
rect 14737 17221 14749 17255
rect 14783 17252 14795 17255
rect 15286 17252 15292 17264
rect 14783 17224 15292 17252
rect 14783 17221 14795 17224
rect 14737 17215 14795 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 16206 17252 16212 17264
rect 16167 17224 16212 17252
rect 16206 17212 16212 17224
rect 16264 17212 16270 17264
rect 17957 17255 18015 17261
rect 17957 17221 17969 17255
rect 18003 17252 18015 17255
rect 18598 17252 18604 17264
rect 18003 17224 18604 17252
rect 18003 17221 18015 17224
rect 17957 17215 18015 17221
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 13081 17187 13139 17193
rect 12860 17156 13032 17184
rect 12860 17144 12866 17156
rect 13004 17116 13032 17156
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 13906 17184 13912 17196
rect 13867 17156 13912 17184
rect 13081 17147 13139 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14090 17144 14096 17196
rect 14148 17184 14154 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14148 17156 14473 17184
rect 14148 17144 14154 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 16482 17184 16488 17196
rect 16443 17156 16488 17184
rect 14461 17147 14519 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 18233 17187 18291 17193
rect 16899 17156 17264 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17236 17128 17264 17156
rect 18233 17153 18245 17187
rect 18279 17184 18291 17187
rect 18506 17184 18512 17196
rect 18279 17156 18512 17184
rect 18279 17153 18291 17156
rect 18233 17147 18291 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18690 17184 18696 17196
rect 18651 17156 18696 17184
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 20254 17184 20260 17196
rect 19567 17156 20260 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 20806 17184 20812 17196
rect 20763 17156 20812 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 6104 17088 7420 17116
rect 11256 17088 12940 17116
rect 13004 17088 13277 17116
rect 8220 17020 9674 17048
rect 4798 16980 4804 16992
rect 4759 16952 4804 16980
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 8220 16980 8248 17020
rect 8662 16980 8668 16992
rect 6880 16952 8248 16980
rect 8623 16952 8668 16980
rect 6880 16940 6886 16952
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9646 16980 9674 17020
rect 11256 16980 11284 17088
rect 11333 17051 11391 17057
rect 11333 17017 11345 17051
rect 11379 17048 11391 17051
rect 12434 17048 12440 17060
rect 11379 17020 12440 17048
rect 11379 17017 11391 17020
rect 11333 17011 11391 17017
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12912 17048 12940 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 17034 17116 17040 17128
rect 16995 17088 17040 17116
rect 13725 17079 13783 17085
rect 13740 17048 13768 17079
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 17218 17116 17224 17128
rect 17179 17088 17224 17116
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18785 17119 18843 17125
rect 18785 17116 18797 17119
rect 18196 17088 18797 17116
rect 18196 17076 18202 17088
rect 18785 17085 18797 17088
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17085 18935 17119
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 18877 17079 18935 17085
rect 18984 17088 19625 17116
rect 17052 17048 17080 17076
rect 18892 17048 18920 17079
rect 12912 17020 13768 17048
rect 14200 17020 16988 17048
rect 17052 17020 18920 17048
rect 12158 16980 12164 16992
rect 9646 16952 11284 16980
rect 12119 16952 12164 16980
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 14200 16980 14228 17020
rect 14366 16980 14372 16992
rect 13044 16952 14228 16980
rect 14327 16952 14372 16980
rect 13044 16940 13050 16952
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 16960 16980 16988 17020
rect 18984 16992 19012 17088
rect 19613 17085 19625 17088
rect 19659 17085 19671 17119
rect 19794 17116 19800 17128
rect 19755 17088 19800 17116
rect 19613 17079 19671 17085
rect 19794 17076 19800 17088
rect 19852 17076 19858 17128
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 21192 17116 21220 17147
rect 20588 17088 21220 17116
rect 20588 17076 20594 17088
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 21082 17048 21088 17060
rect 19300 17020 21088 17048
rect 19300 17008 19306 17020
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 17862 16980 17868 16992
rect 16960 16952 17868 16980
rect 17862 16940 17868 16952
rect 17920 16980 17926 16992
rect 18966 16980 18972 16992
rect 17920 16952 18972 16980
rect 17920 16940 17926 16952
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 20254 16980 20260 16992
rect 20215 16952 20260 16980
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 6270 16776 6276 16788
rect 4632 16748 6276 16776
rect 2884 16680 3188 16708
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 2884 16649 2912 16680
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 1728 16612 2881 16640
rect 1728 16600 1734 16612
rect 2869 16609 2881 16612
rect 2915 16609 2927 16643
rect 3050 16640 3056 16652
rect 2869 16603 2927 16609
rect 2976 16612 3056 16640
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 2133 16575 2191 16581
rect 2133 16572 2145 16575
rect 1811 16544 2145 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 2133 16541 2145 16544
rect 2179 16572 2191 16575
rect 2590 16572 2596 16584
rect 2179 16544 2596 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 2976 16572 3004 16612
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 2823 16544 3004 16572
rect 3160 16572 3188 16680
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4120 16612 4353 16640
rect 4120 16600 4126 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4632 16640 4660 16748
rect 6270 16736 6276 16748
rect 6328 16776 6334 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6328 16748 6377 16776
rect 6328 16736 6334 16748
rect 6365 16745 6377 16748
rect 6411 16776 6423 16779
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6411 16748 6561 16776
rect 6411 16745 6423 16748
rect 6365 16739 6423 16745
rect 6549 16745 6561 16748
rect 6595 16776 6607 16779
rect 6914 16776 6920 16788
rect 6595 16748 6920 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6914 16736 6920 16748
rect 6972 16776 6978 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6972 16748 7021 16776
rect 6972 16736 6978 16748
rect 7009 16745 7021 16748
rect 7055 16776 7067 16779
rect 7055 16748 8616 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 8588 16649 8616 16748
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 16301 16779 16359 16785
rect 8720 16748 16252 16776
rect 8720 16736 8726 16748
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 11146 16708 11152 16720
rect 9272 16680 11152 16708
rect 9272 16668 9278 16680
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 13722 16668 13728 16720
rect 13780 16708 13786 16720
rect 15930 16708 15936 16720
rect 13780 16680 15936 16708
rect 13780 16668 13786 16680
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4632 16612 4721 16640
rect 4430 16572 4436 16584
rect 3160 16544 4436 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 4632 16572 4660 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 4709 16603 4767 16609
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16609 8631 16643
rect 11054 16640 11060 16652
rect 8573 16603 8631 16609
rect 10612 16612 11060 16640
rect 10612 16572 10640 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14550 16640 14556 16652
rect 13872 16612 14556 16640
rect 13872 16600 13878 16612
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 16224 16640 16252 16748
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 16482 16776 16488 16788
rect 16347 16748 16488 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 18138 16776 18144 16788
rect 18099 16748 18144 16776
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18748 16748 19257 16776
rect 18748 16736 18754 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 19245 16739 19303 16745
rect 17954 16708 17960 16720
rect 16776 16680 17960 16708
rect 16776 16649 16804 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18966 16708 18972 16720
rect 18927 16680 18972 16708
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 16761 16643 16819 16649
rect 16224 16612 16712 16640
rect 12158 16572 12164 16584
rect 4580 16544 4660 16572
rect 4908 16544 10640 16572
rect 10704 16544 12164 16572
rect 4580 16532 4586 16544
rect 2685 16507 2743 16513
rect 1964 16476 2452 16504
rect 1964 16445 1992 16476
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16405 2007 16439
rect 2314 16436 2320 16448
rect 2275 16408 2320 16436
rect 1949 16399 2007 16405
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 2424 16436 2452 16476
rect 2685 16473 2697 16507
rect 2731 16504 2743 16507
rect 2958 16504 2964 16516
rect 2731 16476 2964 16504
rect 2731 16473 2743 16476
rect 2685 16467 2743 16473
rect 2958 16464 2964 16476
rect 3016 16464 3022 16516
rect 4246 16504 4252 16516
rect 4207 16476 4252 16504
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 4908 16504 4936 16544
rect 4982 16513 4988 16516
rect 4356 16476 4936 16504
rect 2866 16436 2872 16448
rect 2424 16408 2872 16436
rect 2866 16396 2872 16408
rect 2924 16396 2930 16448
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3384 16408 3801 16436
rect 3384 16396 3390 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 4356 16436 4384 16476
rect 4976 16467 4988 16513
rect 5040 16504 5046 16516
rect 5040 16476 5076 16504
rect 4982 16464 4988 16467
rect 5040 16464 5046 16476
rect 8018 16464 8024 16516
rect 8076 16504 8082 16516
rect 8306 16507 8364 16513
rect 8306 16504 8318 16507
rect 8076 16476 8318 16504
rect 8076 16464 8082 16476
rect 8306 16473 8318 16476
rect 8352 16473 8364 16507
rect 8306 16467 8364 16473
rect 4203 16408 4384 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 6089 16439 6147 16445
rect 6089 16436 6101 16439
rect 4488 16408 6101 16436
rect 4488 16396 4494 16408
rect 6089 16405 6101 16408
rect 6135 16436 6147 16439
rect 7006 16436 7012 16448
rect 6135 16408 7012 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7193 16439 7251 16445
rect 7193 16405 7205 16439
rect 7239 16436 7251 16439
rect 7834 16436 7840 16448
rect 7239 16408 7840 16436
rect 7239 16405 7251 16408
rect 7193 16399 7251 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 10704 16445 10732 16544
rect 12158 16532 12164 16544
rect 12216 16572 12222 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 12216 16544 12265 16572
rect 12216 16532 12222 16544
rect 12253 16541 12265 16544
rect 12299 16572 12311 16575
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12299 16544 12357 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14516 16544 14749 16572
rect 14516 16532 14522 16544
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15013 16575 15071 16581
rect 15013 16572 15025 16575
rect 14976 16544 15025 16572
rect 14976 16532 14982 16544
rect 15013 16541 15025 16544
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15344 16544 15577 16572
rect 15344 16532 15350 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15565 16535 15623 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 12008 16507 12066 16513
rect 12008 16473 12020 16507
rect 12054 16504 12066 16507
rect 12054 16476 12204 16504
rect 12054 16473 12066 16476
rect 12008 16467 12066 16473
rect 10689 16439 10747 16445
rect 10689 16436 10701 16439
rect 9824 16408 10701 16436
rect 9824 16396 9830 16408
rect 10689 16405 10701 16408
rect 10735 16405 10747 16439
rect 10689 16399 10747 16405
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 10873 16439 10931 16445
rect 10873 16436 10885 16439
rect 10836 16408 10885 16436
rect 10836 16396 10842 16408
rect 10873 16405 10885 16408
rect 10919 16405 10931 16439
rect 12176 16436 12204 16476
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 12612 16507 12670 16513
rect 12612 16504 12624 16507
rect 12492 16476 12624 16504
rect 12492 16464 12498 16476
rect 12612 16473 12624 16476
rect 12658 16504 12670 16507
rect 15194 16504 15200 16516
rect 12658 16476 15200 16504
rect 12658 16473 12670 16476
rect 12612 16467 12670 16473
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 16684 16504 16712 16612
rect 16761 16609 16773 16643
rect 16807 16609 16819 16643
rect 16761 16603 16819 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17310 16640 17316 16652
rect 16991 16612 17316 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 17126 16572 17132 16584
rect 17087 16544 17132 16572
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 16684 16476 16896 16504
rect 13722 16436 13728 16448
rect 12176 16408 13728 16436
rect 10873 16399 10931 16405
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 16298 16436 16304 16448
rect 15160 16408 16304 16436
rect 15160 16396 15166 16408
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 16448 16408 16681 16436
rect 16448 16396 16454 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16868 16436 16896 16476
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17405 16507 17463 16513
rect 17405 16504 17417 16507
rect 17000 16476 17417 16504
rect 17000 16464 17006 16476
rect 17405 16473 17417 16476
rect 17451 16473 17463 16507
rect 17405 16467 17463 16473
rect 17310 16436 17316 16448
rect 16868 16408 17316 16436
rect 16669 16399 16727 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2372 16204 2605 16232
rect 2372 16192 2378 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 5902 16232 5908 16244
rect 2593 16195 2651 16201
rect 2792 16204 5908 16232
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 2038 16096 2044 16108
rect 1719 16068 2044 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 2501 16099 2559 16105
rect 2501 16096 2513 16099
rect 2464 16068 2513 16096
rect 2464 16056 2470 16068
rect 2501 16065 2513 16068
rect 2547 16065 2559 16099
rect 2501 16059 2559 16065
rect 2792 16037 2820 16204
rect 5902 16192 5908 16204
rect 5960 16232 5966 16244
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 5960 16204 6377 16232
rect 5960 16192 5966 16204
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 9582 16232 9588 16244
rect 6365 16195 6423 16201
rect 6840 16204 9588 16232
rect 4246 16164 4252 16176
rect 3068 16136 4252 16164
rect 3068 16037 3096 16136
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 6840 16164 6868 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 9766 16232 9772 16244
rect 9727 16204 9772 16232
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 14458 16232 14464 16244
rect 9876 16204 13768 16232
rect 14419 16204 14464 16232
rect 4356 16136 6868 16164
rect 6932 16136 7788 16164
rect 3142 16056 3148 16108
rect 3200 16056 3206 16108
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 4065 16099 4123 16105
rect 4065 16096 4077 16099
rect 3375 16068 4077 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 4065 16065 4077 16068
rect 4111 16096 4123 16099
rect 4356 16096 4384 16136
rect 6932 16108 6960 16136
rect 4111 16068 4384 16096
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 5718 16056 5724 16108
rect 5776 16105 5782 16108
rect 5776 16096 5788 16105
rect 5997 16099 6055 16105
rect 5776 16068 5821 16096
rect 5776 16059 5788 16068
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6914 16096 6920 16108
rect 6043 16068 6920 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 5776 16056 5782 16059
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7760 16105 7788 16136
rect 7834 16124 7840 16176
rect 7892 16164 7898 16176
rect 9876 16164 9904 16204
rect 7892 16136 9904 16164
rect 7892 16124 7898 16136
rect 10318 16124 10324 16176
rect 10376 16124 10382 16176
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 13740 16164 13768 16204
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15102 16232 15108 16244
rect 14875 16204 15108 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15657 16235 15715 16241
rect 15657 16201 15669 16235
rect 15703 16232 15715 16235
rect 16022 16232 16028 16244
rect 15703 16204 16028 16232
rect 15703 16201 15715 16204
rect 15657 16195 15715 16201
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16448 16204 16497 16232
rect 16448 16192 16454 16204
rect 16485 16201 16497 16204
rect 16531 16201 16543 16235
rect 16485 16195 16543 16201
rect 17678 16192 17684 16244
rect 17736 16232 17742 16244
rect 17773 16235 17831 16241
rect 17773 16232 17785 16235
rect 17736 16204 17785 16232
rect 17736 16192 17742 16204
rect 17773 16201 17785 16204
rect 17819 16201 17831 16235
rect 17954 16232 17960 16244
rect 17915 16204 17960 16232
rect 17773 16195 17831 16201
rect 12216 16136 12940 16164
rect 13740 16136 15056 16164
rect 12216 16124 12222 16136
rect 7478 16099 7536 16105
rect 7478 16096 7490 16099
rect 7064 16068 7490 16096
rect 7064 16056 7070 16068
rect 7478 16065 7490 16068
rect 7524 16065 7536 16099
rect 7478 16059 7536 16065
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7791 16068 7941 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 8196 16099 8254 16105
rect 8196 16065 8208 16099
rect 8242 16096 8254 16099
rect 8242 16068 9536 16096
rect 8242 16065 8254 16068
rect 8196 16059 8254 16065
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 15997 2835 16031
rect 2777 15991 2835 15997
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 15997 3111 16031
rect 3053 15991 3111 15997
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15960 1915 15963
rect 3160 15960 3188 16056
rect 9508 16037 9536 16068
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 9950 16096 9956 16108
rect 9824 16068 9956 16096
rect 9824 16056 9830 16068
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 10226 16105 10232 16108
rect 10220 16096 10232 16105
rect 10187 16068 10232 16096
rect 10220 16059 10232 16068
rect 10226 16056 10232 16059
rect 10284 16056 10290 16108
rect 10336 16096 10364 16124
rect 12342 16096 12348 16108
rect 10336 16068 12348 16096
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 12618 16056 12624 16108
rect 12676 16105 12682 16108
rect 12912 16105 12940 16136
rect 12676 16096 12688 16105
rect 12897 16099 12955 16105
rect 12676 16068 12721 16096
rect 12676 16059 12688 16068
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 12676 16056 12682 16059
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 9493 16031 9551 16037
rect 3283 16000 3924 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 1903 15932 3188 15960
rect 1903 15929 1915 15932
rect 1857 15923 1915 15929
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2133 15895 2191 15901
rect 2133 15892 2145 15895
rect 2004 15864 2145 15892
rect 2004 15852 2010 15864
rect 2133 15861 2145 15864
rect 2179 15861 2191 15895
rect 2133 15855 2191 15861
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 3896 15901 3924 16000
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9674 16028 9680 16040
rect 9539 16000 9680 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 15028 16037 15056 16136
rect 15194 16124 15200 16176
rect 15252 16164 15258 16176
rect 17586 16164 17592 16176
rect 15252 16136 17592 16164
rect 15252 16124 15258 16136
rect 17586 16124 17592 16136
rect 17644 16124 17650 16176
rect 17788 16164 17816 16195
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 18417 16167 18475 16173
rect 18417 16164 18429 16167
rect 17788 16136 18429 16164
rect 18417 16133 18429 16136
rect 18463 16133 18475 16167
rect 20714 16164 20720 16176
rect 20675 16136 20720 16164
rect 18417 16127 18475 16133
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 16022 16096 16028 16108
rect 15712 16068 16028 16096
rect 15712 16056 15718 16068
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16482 16096 16488 16108
rect 16163 16068 16488 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 17034 16096 17040 16108
rect 16995 16068 17040 16096
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18325 16099 18383 16105
rect 18325 16096 18337 16099
rect 18012 16068 18337 16096
rect 18012 16056 18018 16068
rect 18325 16065 18337 16068
rect 18371 16096 18383 16099
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 18371 16068 18797 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18785 16065 18797 16068
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 19610 16056 19616 16108
rect 19668 16096 19674 16108
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19668 16068 20453 16096
rect 19668 16056 19674 16068
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 14921 16031 14979 16037
rect 11256 16000 11928 16028
rect 4246 15960 4252 15972
rect 4159 15932 4252 15960
rect 4246 15920 4252 15932
rect 4304 15960 4310 15972
rect 4798 15960 4804 15972
rect 4304 15932 4804 15960
rect 4304 15920 4310 15932
rect 4798 15920 4804 15932
rect 4856 15960 4862 15972
rect 4856 15932 5120 15960
rect 4856 15920 4862 15932
rect 3697 15895 3755 15901
rect 3697 15892 3709 15895
rect 3476 15864 3709 15892
rect 3476 15852 3482 15864
rect 3697 15861 3709 15864
rect 3743 15861 3755 15895
rect 3697 15855 3755 15861
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 4338 15892 4344 15904
rect 3927 15864 4344 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15892 4678 15904
rect 4982 15892 4988 15904
rect 4672 15864 4988 15892
rect 4672 15852 4678 15864
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5092 15892 5120 15932
rect 9140 15932 9628 15960
rect 5350 15892 5356 15904
rect 5092 15864 5356 15892
rect 5350 15852 5356 15864
rect 5408 15892 5414 15904
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 5408 15864 6193 15892
rect 5408 15852 5414 15864
rect 6181 15861 6193 15864
rect 6227 15892 6239 15895
rect 7926 15892 7932 15904
rect 6227 15864 7932 15892
rect 6227 15861 6239 15864
rect 6181 15855 6239 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 9140 15892 9168 15932
rect 8168 15864 9168 15892
rect 8168 15852 8174 15864
rect 9214 15852 9220 15904
rect 9272 15892 9278 15904
rect 9309 15895 9367 15901
rect 9309 15892 9321 15895
rect 9272 15864 9321 15892
rect 9272 15852 9278 15864
rect 9309 15861 9321 15864
rect 9355 15861 9367 15895
rect 9600 15892 9628 15932
rect 11256 15892 11284 16000
rect 11333 15963 11391 15969
rect 11333 15929 11345 15963
rect 11379 15960 11391 15963
rect 11698 15960 11704 15972
rect 11379 15932 11704 15960
rect 11379 15929 11391 15932
rect 11333 15923 11391 15929
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 11900 15960 11928 16000
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15930 16028 15936 16040
rect 15891 16000 15936 16028
rect 15013 15991 15071 15997
rect 14936 15960 14964 15991
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16850 15988 16856 16040
rect 16908 16028 16914 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 16908 16000 17141 16028
rect 16908 15988 16914 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17310 16028 17316 16040
rect 17271 16000 17316 16028
rect 17129 15991 17187 15997
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 18230 15988 18236 16040
rect 18288 16028 18294 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18288 16000 18521 16028
rect 18288 15988 18294 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 17402 15960 17408 15972
rect 11900 15932 12020 15960
rect 14936 15932 17408 15960
rect 11514 15892 11520 15904
rect 9600 15864 11284 15892
rect 11427 15864 11520 15892
rect 9309 15855 9367 15861
rect 11514 15852 11520 15864
rect 11572 15892 11578 15904
rect 11882 15892 11888 15904
rect 11572 15864 11888 15892
rect 11572 15852 11578 15864
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 11992 15892 12020 15932
rect 17402 15920 17408 15932
rect 17460 15920 17466 15972
rect 15562 15892 15568 15904
rect 11992 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 15712 15864 16681 15892
rect 15712 15852 15718 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4522 15688 4528 15700
rect 4019 15660 4528 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 4522 15648 4528 15660
rect 4580 15688 4586 15700
rect 4580 15660 5488 15688
rect 4580 15648 4586 15660
rect 5460 15561 5488 15660
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6972 15660 7021 15688
rect 6972 15648 6978 15660
rect 7009 15657 7021 15660
rect 7055 15688 7067 15691
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 7055 15660 7205 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 7193 15657 7205 15660
rect 7239 15688 7251 15691
rect 7239 15660 8800 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 5537 15623 5595 15629
rect 5537 15589 5549 15623
rect 5583 15620 5595 15623
rect 5583 15592 5948 15620
rect 5583 15589 5595 15592
rect 5537 15583 5595 15589
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 1946 15484 1952 15496
rect 1907 15456 1952 15484
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 5189 15487 5247 15493
rect 5189 15453 5201 15487
rect 5235 15484 5247 15487
rect 5350 15484 5356 15496
rect 5235 15456 5356 15484
rect 5235 15453 5247 15456
rect 5189 15447 5247 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 5920 15484 5948 15592
rect 6932 15561 6960 15648
rect 8772 15561 8800 15660
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 10008 15660 10425 15688
rect 10008 15648 10014 15660
rect 10413 15657 10425 15660
rect 10459 15688 10471 15691
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 10459 15660 12081 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12618 15688 12624 15700
rect 12069 15651 12127 15657
rect 12268 15660 12624 15688
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 10321 15623 10379 15629
rect 10321 15620 10333 15623
rect 10284 15592 10333 15620
rect 10284 15580 10290 15592
rect 10321 15589 10333 15592
rect 10367 15589 10379 15623
rect 10321 15583 10379 15589
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8803 15524 8953 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 10428 15552 10456 15651
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10428 15524 10609 15552
rect 8941 15515 8999 15521
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 7098 15484 7104 15496
rect 5920 15456 7104 15484
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 9214 15493 9220 15496
rect 9208 15484 9220 15493
rect 9127 15456 9220 15484
rect 9208 15447 9220 15456
rect 9272 15484 9278 15496
rect 11882 15484 11888 15496
rect 9272 15456 11888 15484
rect 9214 15444 9220 15447
rect 9272 15444 9278 15456
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 2130 15376 2136 15428
rect 2188 15416 2194 15428
rect 2225 15419 2283 15425
rect 2225 15416 2237 15419
rect 2188 15388 2237 15416
rect 2188 15376 2194 15388
rect 2225 15385 2237 15388
rect 2271 15385 2283 15419
rect 2225 15379 2283 15385
rect 4338 15376 4344 15428
rect 4396 15416 4402 15428
rect 5626 15416 5632 15428
rect 4396 15388 5632 15416
rect 4396 15376 4402 15388
rect 5626 15376 5632 15388
rect 5684 15416 5690 15428
rect 6454 15416 6460 15428
rect 5684 15388 6460 15416
rect 5684 15376 5690 15388
rect 6454 15376 6460 15388
rect 6512 15376 6518 15428
rect 6672 15419 6730 15425
rect 6672 15385 6684 15419
rect 6718 15416 6730 15419
rect 7650 15416 7656 15428
rect 6718 15388 7656 15416
rect 6718 15385 6730 15388
rect 6672 15379 6730 15385
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 8512 15419 8570 15425
rect 8512 15385 8524 15419
rect 8558 15416 8570 15419
rect 8558 15388 10640 15416
rect 8558 15385 8570 15388
rect 8512 15379 8570 15385
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 4065 15351 4123 15357
rect 4065 15348 4077 15351
rect 4028 15320 4077 15348
rect 4028 15308 4034 15320
rect 4065 15317 4077 15320
rect 4111 15317 4123 15351
rect 4065 15311 4123 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7377 15351 7435 15357
rect 7377 15348 7389 15351
rect 7064 15320 7389 15348
rect 7064 15308 7070 15320
rect 7377 15317 7389 15320
rect 7423 15317 7435 15351
rect 7377 15311 7435 15317
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9582 15348 9588 15360
rect 9364 15320 9588 15348
rect 9364 15308 9370 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 10612 15348 10640 15388
rect 10686 15376 10692 15428
rect 10744 15416 10750 15428
rect 10842 15419 10900 15425
rect 10842 15416 10854 15419
rect 10744 15388 10854 15416
rect 10744 15376 10750 15388
rect 10842 15385 10854 15388
rect 10888 15385 10900 15419
rect 12268 15416 12296 15660
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 13872 15660 14289 15688
rect 13872 15648 13878 15660
rect 14277 15657 14289 15660
rect 14323 15688 14335 15691
rect 14826 15688 14832 15700
rect 14323 15660 14832 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 15286 15688 15292 15700
rect 15247 15660 15292 15688
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 15562 15648 15568 15700
rect 15620 15688 15626 15700
rect 16390 15688 16396 15700
rect 15620 15660 16396 15688
rect 15620 15648 15626 15660
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 17218 15688 17224 15700
rect 17179 15660 17224 15688
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17402 15688 17408 15700
rect 17363 15660 17408 15688
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 19981 15623 20039 15629
rect 13780 15592 19380 15620
rect 13780 15580 13786 15592
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 12676 15524 14105 15552
rect 12676 15512 12682 15524
rect 14093 15521 14105 15524
rect 14139 15552 14151 15555
rect 14553 15555 14611 15561
rect 14553 15552 14565 15555
rect 14139 15524 14565 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14553 15521 14565 15524
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15521 15899 15555
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 15841 15515 15899 15521
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 15856 15484 15884 15515
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 19352 15561 19380 15592
rect 19981 15589 19993 15623
rect 20027 15589 20039 15623
rect 19981 15583 20039 15589
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 16632 15524 17969 15552
rect 16632 15512 16638 15524
rect 17957 15521 17969 15524
rect 18003 15521 18015 15555
rect 17957 15515 18015 15521
rect 19337 15555 19395 15561
rect 19337 15521 19349 15555
rect 19383 15521 19395 15555
rect 19337 15515 19395 15521
rect 12400 15456 15884 15484
rect 16393 15487 16451 15493
rect 12400 15444 12406 15456
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 17034 15484 17040 15496
rect 16439 15456 17040 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 17034 15444 17040 15456
rect 17092 15444 17098 15496
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17276 15456 17877 15484
rect 17276 15444 17282 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 18230 15484 18236 15496
rect 18191 15456 18236 15484
rect 17865 15447 17923 15453
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 19996 15484 20024 15583
rect 20530 15552 20536 15564
rect 20491 15524 20536 15552
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 20257 15487 20315 15493
rect 20257 15484 20269 15487
rect 19996 15456 20269 15484
rect 20257 15453 20269 15456
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 13814 15416 13820 15428
rect 10842 15379 10900 15385
rect 11992 15388 13400 15416
rect 13775 15388 13820 15416
rect 11514 15348 11520 15360
rect 10612 15320 11520 15348
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 11992 15357 12020 15388
rect 11977 15351 12035 15357
rect 11977 15317 11989 15351
rect 12023 15317 12035 15351
rect 11977 15311 12035 15317
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 13262 15348 13268 15360
rect 12308 15320 13268 15348
rect 12308 15308 12314 15320
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13372 15348 13400 15388
rect 13814 15376 13820 15388
rect 13872 15416 13878 15428
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 13872 15388 14749 15416
rect 13872 15376 13878 15388
rect 14737 15385 14749 15388
rect 14783 15385 14795 15419
rect 14737 15379 14795 15385
rect 14826 15376 14832 15428
rect 14884 15416 14890 15428
rect 15470 15416 15476 15428
rect 14884 15388 14929 15416
rect 15028 15388 15476 15416
rect 14884 15376 14890 15388
rect 15028 15348 15056 15388
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 15654 15416 15660 15428
rect 15615 15388 15660 15416
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 15749 15419 15807 15425
rect 15749 15385 15761 15419
rect 15795 15416 15807 15419
rect 16942 15416 16948 15428
rect 15795 15388 16948 15416
rect 15795 15385 15807 15388
rect 15749 15379 15807 15385
rect 16942 15376 16948 15388
rect 17000 15376 17006 15428
rect 20530 15416 20536 15428
rect 17052 15388 20536 15416
rect 17052 15360 17080 15388
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 13372 15320 15056 15348
rect 15197 15351 15255 15357
rect 15197 15317 15209 15351
rect 15243 15348 15255 15351
rect 15930 15348 15936 15360
rect 15243 15320 15936 15348
rect 15243 15317 15255 15320
rect 15197 15311 15255 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 16850 15348 16856 15360
rect 16763 15320 16856 15348
rect 16850 15308 16856 15320
rect 16908 15348 16914 15360
rect 17034 15348 17040 15360
rect 16908 15320 17040 15348
rect 16908 15308 16914 15320
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17770 15348 17776 15360
rect 17683 15320 17776 15348
rect 17770 15308 17776 15320
rect 17828 15348 17834 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 17828 15320 18521 15348
rect 17828 15308 17834 15320
rect 18509 15317 18521 15320
rect 18555 15348 18567 15351
rect 18874 15348 18880 15360
rect 18555 15320 18880 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19518 15348 19524 15360
rect 19479 15320 19524 15348
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 19702 15348 19708 15360
rect 19659 15320 19708 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 3234 15144 3240 15156
rect 1995 15116 3240 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 6457 15147 6515 15153
rect 4479 15116 6408 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 3786 15076 3792 15088
rect 3747 15048 3792 15076
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15076 3939 15079
rect 4448 15076 4476 15107
rect 3927 15048 4476 15076
rect 3927 15045 3939 15048
rect 3881 15039 3939 15045
rect 4522 15036 4528 15088
rect 4580 15076 4586 15088
rect 4617 15079 4675 15085
rect 4617 15076 4629 15079
rect 4580 15048 4629 15076
rect 4580 15036 4586 15048
rect 4617 15045 4629 15048
rect 4663 15045 4675 15079
rect 6380 15076 6408 15116
rect 6457 15113 6469 15147
rect 6503 15144 6515 15147
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6503 15116 6653 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6641 15113 6653 15116
rect 6687 15144 6699 15147
rect 6914 15144 6920 15156
rect 6687 15116 6920 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6914 15104 6920 15116
rect 6972 15144 6978 15156
rect 7009 15147 7067 15153
rect 7009 15144 7021 15147
rect 6972 15116 7021 15144
rect 6972 15104 6978 15116
rect 7009 15113 7021 15116
rect 7055 15144 7067 15147
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 7055 15116 7665 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7653 15113 7665 15116
rect 7699 15144 7711 15147
rect 9217 15147 9275 15153
rect 7699 15116 7880 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 6380 15048 7788 15076
rect 4617 15039 4675 15045
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 4632 15008 4660 15039
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4304 14980 4813 15008
rect 4304 14968 4310 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 5057 15011 5115 15017
rect 5057 15008 5069 15011
rect 4801 14971 4859 14977
rect 4908 14980 5069 15008
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14909 3755 14943
rect 3697 14903 3755 14909
rect 3712 14804 3740 14903
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4908 14940 4936 14980
rect 5057 14977 5069 14980
rect 5103 14977 5115 15011
rect 5057 14971 5115 14977
rect 4120 14912 4936 14940
rect 4120 14900 4126 14912
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14872 4307 14875
rect 4798 14872 4804 14884
rect 4295 14844 4804 14872
rect 4295 14841 4307 14844
rect 4249 14835 4307 14841
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 7006 14872 7012 14884
rect 5736 14844 7012 14872
rect 5736 14804 5764 14844
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 3712 14776 5764 14804
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5868 14776 6193 14804
rect 5868 14764 5874 14776
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6181 14767 6239 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 7650 14804 7656 14816
rect 7331 14776 7656 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 7760 14804 7788 15048
rect 7852 15017 7880 15116
rect 9217 15113 9229 15147
rect 9263 15144 9275 15147
rect 9306 15144 9312 15156
rect 9263 15116 9312 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9950 15144 9956 15156
rect 9447 15116 9956 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 13173 15147 13231 15153
rect 13173 15144 13185 15147
rect 10060 15116 13185 15144
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 10060 15076 10088 15116
rect 13173 15113 13185 15116
rect 13219 15113 13231 15147
rect 13173 15107 13231 15113
rect 13188 15076 13216 15107
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13320 15116 13461 15144
rect 13320 15104 13326 15116
rect 13449 15113 13461 15116
rect 13495 15144 13507 15147
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 13495 15116 14013 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 14001 15113 14013 15116
rect 14047 15144 14059 15147
rect 14047 15116 15056 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 15028 15076 15056 15116
rect 15102 15104 15108 15156
rect 15160 15144 15166 15156
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 15160 15116 15761 15144
rect 15160 15104 15166 15116
rect 15749 15113 15761 15116
rect 15795 15113 15807 15147
rect 15749 15107 15807 15113
rect 16942 15104 16948 15156
rect 17000 15144 17006 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 17000 15116 17233 15144
rect 17000 15104 17006 15116
rect 17221 15113 17233 15116
rect 17267 15113 17279 15147
rect 17221 15107 17279 15113
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19153 15147 19211 15153
rect 19153 15144 19165 15147
rect 19116 15116 19165 15144
rect 19116 15104 19122 15116
rect 19153 15113 19165 15116
rect 19199 15113 19211 15147
rect 19153 15107 19211 15113
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19576 15116 19625 15144
rect 19576 15104 19582 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 19702 15104 19708 15156
rect 19760 15144 19766 15156
rect 19760 15116 19805 15144
rect 19760 15104 19766 15116
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20993 15147 21051 15153
rect 20993 15144 21005 15147
rect 20404 15116 21005 15144
rect 20404 15104 20410 15116
rect 20993 15113 21005 15116
rect 21039 15113 21051 15147
rect 21358 15144 21364 15156
rect 21319 15116 21364 15144
rect 20993 15107 21051 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 15286 15076 15292 15088
rect 7984 15048 10088 15076
rect 12544 15048 13124 15076
rect 13188 15048 14136 15076
rect 15028 15048 15292 15076
rect 7984 15036 7990 15048
rect 8110 15017 8116 15020
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 8104 15008 8116 15017
rect 8071 14980 8116 15008
rect 7837 14971 7895 14977
rect 8104 14971 8116 14980
rect 8110 14968 8116 14971
rect 8168 14968 8174 15020
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 12544 15008 12572 15048
rect 8628 14980 12572 15008
rect 12641 15011 12699 15017
rect 8628 14968 8634 14980
rect 12641 14977 12653 15011
rect 12687 15008 12699 15011
rect 12687 14980 12848 15008
rect 12687 14977 12699 14980
rect 12641 14971 12699 14977
rect 9214 14900 9220 14952
rect 9272 14940 9278 14952
rect 12820 14940 12848 14980
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 12952 14980 12997 15008
rect 12952 14968 12958 14980
rect 12986 14940 12992 14952
rect 9272 14912 11652 14940
rect 12820 14912 12992 14940
rect 9272 14900 9278 14912
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11112 14844 11529 14872
rect 11112 14832 11118 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 8570 14804 8576 14816
rect 7760 14776 8576 14804
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 11020 14776 11253 14804
rect 11020 14764 11026 14776
rect 11241 14773 11253 14776
rect 11287 14773 11299 14807
rect 11624 14804 11652 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13096 14940 13124 15048
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 15008 13967 15011
rect 13998 15008 14004 15020
rect 13955 14980 14004 15008
rect 13955 14977 13967 14980
rect 13909 14971 13967 14977
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 14108 14949 14136 15048
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 16298 15036 16304 15088
rect 16356 15076 16362 15088
rect 17589 15079 17647 15085
rect 16356 15048 17172 15076
rect 16356 15036 16362 15048
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14752 14980 15209 15008
rect 14093 14943 14151 14949
rect 13096 14912 13676 14940
rect 13541 14875 13599 14881
rect 13541 14872 13553 14875
rect 13004 14844 13553 14872
rect 13004 14804 13032 14844
rect 13541 14841 13553 14844
rect 13587 14841 13599 14875
rect 13648 14872 13676 14912
rect 14093 14909 14105 14943
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14182 14900 14188 14952
rect 14240 14940 14246 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14240 14912 14473 14940
rect 14240 14900 14246 14912
rect 14461 14909 14473 14912
rect 14507 14940 14519 14943
rect 14642 14940 14648 14952
rect 14507 14912 14648 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 14553 14875 14611 14881
rect 14553 14872 14565 14875
rect 13648 14844 14565 14872
rect 13541 14835 13599 14841
rect 14553 14841 14565 14844
rect 14599 14872 14611 14875
rect 14752 14872 14780 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16163 14980 16681 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 15160 14912 15301 14940
rect 15160 14900 15166 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 16209 14943 16267 14949
rect 15436 14912 15481 14940
rect 15436 14900 15442 14912
rect 16209 14909 16221 14943
rect 16255 14909 16267 14943
rect 16390 14940 16396 14952
rect 16351 14912 16396 14940
rect 16209 14903 16267 14909
rect 14599 14844 14780 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 11624 14776 13032 14804
rect 11241 14767 11299 14773
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14700 14776 14841 14804
rect 14700 14764 14706 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 16224 14804 16252 14903
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 17144 14949 17172 15048
rect 17589 15045 17601 15079
rect 17635 15076 17647 15079
rect 17678 15076 17684 15088
rect 17635 15048 17684 15076
rect 17635 15045 17647 15048
rect 17589 15039 17647 15045
rect 17678 15036 17684 15048
rect 17736 15076 17742 15088
rect 18230 15076 18236 15088
rect 17736 15048 18236 15076
rect 17736 15036 17742 15048
rect 18230 15036 18236 15048
rect 18288 15036 18294 15088
rect 18417 15079 18475 15085
rect 18417 15045 18429 15079
rect 18463 15076 18475 15079
rect 19978 15076 19984 15088
rect 18463 15048 19984 15076
rect 18463 15045 18475 15048
rect 18417 15039 18475 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 20211 15048 20392 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 20364 15020 20392 15048
rect 20530 15036 20536 15088
rect 20588 15076 20594 15088
rect 20625 15079 20683 15085
rect 20625 15076 20637 15079
rect 20588 15048 20637 15076
rect 20588 15036 20594 15048
rect 20625 15045 20637 15048
rect 20671 15045 20683 15079
rect 20625 15039 20683 15045
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 17368 14980 17816 15008
rect 17368 14968 17374 14980
rect 17788 14949 17816 14980
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 19116 14980 19257 15008
rect 19116 14968 19122 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 20070 15008 20076 15020
rect 20031 14980 20076 15008
rect 19245 14971 19303 14977
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 20640 15008 20668 15039
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20640 14980 20821 15008
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 21174 15008 21180 15020
rect 21135 14980 21180 15008
rect 20809 14971 20867 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17681 14943 17739 14949
rect 17681 14940 17693 14943
rect 17175 14912 17693 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17681 14909 17693 14912
rect 17727 14909 17739 14943
rect 17681 14903 17739 14909
rect 17773 14943 17831 14949
rect 17773 14909 17785 14943
rect 17819 14909 17831 14943
rect 18138 14940 18144 14952
rect 18099 14912 18144 14940
rect 17773 14903 17831 14909
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 18322 14940 18328 14952
rect 18283 14912 18328 14940
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14909 20315 14943
rect 20257 14903 20315 14909
rect 17586 14832 17592 14884
rect 17644 14872 17650 14884
rect 18984 14872 19012 14903
rect 20272 14872 20300 14903
rect 17644 14844 20300 14872
rect 17644 14832 17650 14844
rect 15252 14776 16252 14804
rect 15252 14764 15258 14776
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 17862 14804 17868 14816
rect 17276 14776 17868 14804
rect 17276 14764 17282 14776
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 18782 14804 18788 14816
rect 18743 14776 18788 14804
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 5442 14600 5448 14612
rect 4212 14572 5448 14600
rect 4212 14560 4218 14572
rect 5442 14560 5448 14572
rect 5500 14600 5506 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5500 14572 5641 14600
rect 5500 14560 5506 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 6914 14600 6920 14612
rect 5629 14563 5687 14569
rect 5736 14572 6920 14600
rect 3326 14464 3332 14476
rect 3287 14436 3332 14464
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14433 3571 14467
rect 4246 14464 4252 14476
rect 4207 14436 4252 14464
rect 3513 14427 3571 14433
rect 3528 14396 3556 14427
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 5736 14473 5764 14572
rect 6914 14560 6920 14572
rect 6972 14600 6978 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6972 14572 7205 14600
rect 6972 14560 6978 14572
rect 7193 14569 7205 14572
rect 7239 14600 7251 14603
rect 7239 14572 8800 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 7742 14464 7748 14476
rect 7524 14436 7748 14464
rect 7524 14424 7530 14436
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 8772 14473 8800 14572
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10962 14600 10968 14612
rect 10008 14572 10968 14600
rect 10008 14560 10014 14572
rect 10962 14560 10968 14572
rect 11020 14600 11026 14612
rect 11149 14603 11207 14609
rect 11149 14600 11161 14603
rect 11020 14572 11161 14600
rect 11020 14560 11026 14572
rect 11149 14569 11161 14572
rect 11195 14569 11207 14603
rect 12434 14600 12440 14612
rect 11149 14563 11207 14569
rect 11348 14572 12440 14600
rect 10870 14492 10876 14544
rect 10928 14532 10934 14544
rect 11348 14532 11376 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 15378 14600 15384 14612
rect 12584 14572 15384 14600
rect 12584 14560 12590 14572
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 17773 14603 17831 14609
rect 17773 14569 17785 14603
rect 17819 14600 17831 14603
rect 18322 14600 18328 14612
rect 17819 14572 18328 14600
rect 17819 14569 17831 14572
rect 17773 14563 17831 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 20622 14560 20628 14612
rect 20680 14600 20686 14612
rect 20993 14603 21051 14609
rect 20993 14600 21005 14603
rect 20680 14572 21005 14600
rect 20680 14560 20686 14572
rect 20993 14569 21005 14572
rect 21039 14569 21051 14603
rect 20993 14563 21051 14569
rect 13630 14532 13636 14544
rect 10928 14504 11376 14532
rect 13591 14504 13636 14532
rect 10928 14492 10934 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 14093 14535 14151 14541
rect 14093 14501 14105 14535
rect 14139 14532 14151 14535
rect 15102 14532 15108 14544
rect 14139 14504 15108 14532
rect 14139 14501 14151 14504
rect 14093 14495 14151 14501
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 16390 14532 16396 14544
rect 16080 14504 16396 14532
rect 16080 14492 16086 14504
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 20530 14532 20536 14544
rect 17144 14504 20536 14532
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14433 8815 14467
rect 11422 14464 11428 14476
rect 8757 14427 8815 14433
rect 10888 14436 11428 14464
rect 5810 14396 5816 14408
rect 3528 14368 5816 14396
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 10888 14396 10916 14436
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 14553 14467 14611 14473
rect 14553 14464 14565 14467
rect 14424 14436 14565 14464
rect 14424 14424 14430 14436
rect 14553 14433 14565 14436
rect 14599 14433 14611 14467
rect 14553 14427 14611 14433
rect 14645 14467 14703 14473
rect 14645 14433 14657 14467
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 6604 14368 10916 14396
rect 6604 14356 6610 14368
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 12713 14399 12771 14405
rect 12713 14396 12725 14399
rect 11020 14368 12725 14396
rect 11020 14356 11026 14368
rect 12713 14365 12725 14368
rect 12759 14396 12771 14399
rect 12802 14396 12808 14408
rect 12759 14368 12808 14396
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 14660 14396 14688 14427
rect 14826 14424 14832 14476
rect 14884 14464 14890 14476
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 14884 14436 14933 14464
rect 14884 14424 14890 14436
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 16206 14424 16212 14476
rect 16264 14464 16270 14476
rect 17144 14473 17172 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 16264 14436 17141 14464
rect 16264 14424 16270 14436
rect 17129 14433 17141 14436
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17494 14464 17500 14476
rect 17359 14436 17500 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 18509 14467 18567 14473
rect 18196 14436 18368 14464
rect 18196 14424 18202 14436
rect 18046 14396 18052 14408
rect 13832 14368 14688 14396
rect 17328 14368 18052 14396
rect 4157 14331 4215 14337
rect 4157 14297 4169 14331
rect 4203 14328 4215 14331
rect 4516 14331 4574 14337
rect 4516 14328 4528 14331
rect 4203 14300 4528 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 4516 14297 4528 14300
rect 4562 14328 4574 14331
rect 5350 14328 5356 14340
rect 4562 14300 5356 14328
rect 4562 14297 4574 14300
rect 4516 14291 4574 14297
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 5966 14331 6024 14337
rect 5966 14328 5978 14331
rect 5500 14300 5978 14328
rect 5500 14288 5506 14300
rect 5966 14297 5978 14300
rect 6012 14297 6024 14331
rect 8386 14328 8392 14340
rect 5966 14291 6024 14297
rect 7116 14300 8392 14328
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 2958 14260 2964 14272
rect 2915 14232 2964 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 3234 14260 3240 14272
rect 3195 14232 3240 14260
rect 3234 14220 3240 14232
rect 3292 14220 3298 14272
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14260 4031 14263
rect 4338 14260 4344 14272
rect 4019 14232 4344 14260
rect 4019 14229 4031 14232
rect 3973 14223 4031 14229
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 7116 14269 7144 14300
rect 8386 14288 8392 14300
rect 8444 14288 8450 14340
rect 8512 14331 8570 14337
rect 8512 14297 8524 14331
rect 8558 14328 8570 14331
rect 10318 14328 10324 14340
rect 8558 14300 10324 14328
rect 8558 14297 8570 14300
rect 8512 14291 8570 14297
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 10502 14288 10508 14340
rect 10560 14328 10566 14340
rect 12342 14328 12348 14340
rect 10560 14300 12348 14328
rect 10560 14288 10566 14300
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 12468 14331 12526 14337
rect 12468 14297 12480 14331
rect 12514 14328 12526 14331
rect 12894 14328 12900 14340
rect 12514 14300 12900 14328
rect 12514 14297 12526 14300
rect 12468 14291 12526 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13832 14337 13860 14368
rect 13817 14331 13875 14337
rect 13817 14328 13829 14331
rect 13464 14300 13829 14328
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14229 7159 14263
rect 7101 14223 7159 14229
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 8110 14260 8116 14272
rect 7423 14232 8116 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 8110 14220 8116 14232
rect 8168 14260 8174 14272
rect 10042 14260 10048 14272
rect 8168 14232 10048 14260
rect 8168 14220 8174 14232
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 10928 14232 11345 14260
rect 10928 14220 10934 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 13464 14260 13492 14300
rect 13817 14297 13829 14300
rect 13863 14297 13875 14331
rect 17328 14328 17356 14368
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 18340 14396 18368 14436
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 18598 14464 18604 14476
rect 18555 14436 18604 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 21174 14464 21180 14476
rect 19659 14436 21180 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 18340 14368 18705 14396
rect 18693 14365 18705 14368
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 19337 14399 19395 14405
rect 19337 14396 19349 14399
rect 18840 14368 19349 14396
rect 18840 14356 18846 14368
rect 19337 14365 19349 14368
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 13817 14291 13875 14297
rect 14476 14300 17356 14328
rect 17405 14331 17463 14337
rect 11480 14232 13492 14260
rect 11480 14220 11486 14232
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 14476 14269 14504 14300
rect 17405 14297 17417 14331
rect 17451 14328 17463 14331
rect 18248 14328 18276 14356
rect 20824 14328 20852 14359
rect 21177 14331 21235 14337
rect 21177 14328 21189 14331
rect 17451 14300 17908 14328
rect 18248 14300 21189 14328
rect 17451 14297 17463 14300
rect 17405 14291 17463 14297
rect 14461 14263 14519 14269
rect 14461 14260 14473 14263
rect 13688 14232 14473 14260
rect 13688 14220 13694 14232
rect 14461 14229 14473 14232
rect 14507 14229 14519 14263
rect 14461 14223 14519 14229
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 17880 14269 17908 14300
rect 21177 14297 21189 14300
rect 21223 14297 21235 14331
rect 21177 14291 21235 14297
rect 15565 14263 15623 14269
rect 15565 14260 15577 14263
rect 15252 14232 15577 14260
rect 15252 14220 15258 14232
rect 15565 14229 15577 14232
rect 15611 14229 15623 14263
rect 15565 14223 15623 14229
rect 17865 14263 17923 14269
rect 17865 14229 17877 14263
rect 17911 14229 17923 14263
rect 17865 14223 17923 14229
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 18233 14263 18291 14269
rect 18233 14260 18245 14263
rect 18196 14232 18245 14260
rect 18196 14220 18202 14232
rect 18233 14229 18245 14232
rect 18279 14229 18291 14263
rect 18233 14223 18291 14229
rect 18325 14263 18383 14269
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 18690 14260 18696 14272
rect 18371 14232 18696 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 20622 14220 20628 14272
rect 20680 14260 20686 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 20680 14232 20729 14260
rect 20680 14220 20686 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 1949 14059 2007 14065
rect 1949 14025 1961 14059
rect 1995 14056 2007 14059
rect 2774 14056 2780 14068
rect 1995 14028 2780 14056
rect 1995 14025 2007 14028
rect 1949 14019 2007 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 3476 14028 3525 14056
rect 3476 14016 3482 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 3513 14019 3571 14025
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 4525 14059 4583 14065
rect 4525 14056 4537 14059
rect 4120 14028 4537 14056
rect 4120 14016 4126 14028
rect 4525 14025 4537 14028
rect 4571 14025 4583 14059
rect 6181 14059 6239 14065
rect 6181 14056 6193 14059
rect 4525 14019 4583 14025
rect 5736 14028 6193 14056
rect 5534 13988 5540 14000
rect 3436 13960 5540 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 1946 13920 1952 13932
rect 1811 13892 1952 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2179 13892 2697 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 2685 13889 2697 13892
rect 2731 13889 2743 13923
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2685 13883 2743 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3436 13929 3464 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 5649 13991 5707 13997
rect 5649 13957 5661 13991
rect 5695 13988 5707 13991
rect 5736 13988 5764 14028
rect 6181 14025 6193 14028
rect 6227 14056 6239 14059
rect 7466 14056 7472 14068
rect 6227 14028 7472 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 9214 14056 9220 14068
rect 7760 14028 9220 14056
rect 5695 13960 5764 13988
rect 5695 13957 5707 13960
rect 5649 13951 5707 13957
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 7760 13988 7788 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 9447 14028 9781 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9769 14025 9781 14028
rect 9815 14056 9827 14059
rect 9950 14056 9956 14068
rect 9815 14028 9956 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 8570 13988 8576 14000
rect 5868 13960 7788 13988
rect 7852 13960 8576 13988
rect 5868 13948 5874 13960
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3970 13920 3976 13932
rect 3421 13883 3479 13889
rect 3712 13892 3976 13920
rect 3712 13861 3740 13892
rect 3970 13880 3976 13892
rect 4028 13920 4034 13932
rect 7852 13929 7880 13960
rect 8570 13948 8576 13960
rect 8628 13988 8634 14000
rect 9416 13988 9444 14019
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 11204 14028 11345 14056
rect 11204 14016 11210 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 16574 14056 16580 14068
rect 12492 14028 16580 14056
rect 12492 14016 12498 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 17460 14028 17509 14056
rect 17460 14016 17466 14028
rect 17497 14025 17509 14028
rect 17543 14056 17555 14059
rect 18598 14056 18604 14068
rect 17543 14028 18604 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19337 14059 19395 14065
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19886 14056 19892 14068
rect 19383 14028 19892 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20257 14059 20315 14065
rect 20257 14056 20269 14059
rect 20128 14028 20269 14056
rect 20128 14016 20134 14028
rect 20257 14025 20269 14028
rect 20303 14025 20315 14059
rect 20622 14056 20628 14068
rect 20583 14028 20628 14056
rect 20257 14019 20315 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 8628 13960 9444 13988
rect 8628 13948 8634 13960
rect 7478 13923 7536 13929
rect 7478 13920 7490 13923
rect 4028 13892 7490 13920
rect 4028 13880 4034 13892
rect 7478 13889 7490 13892
rect 7524 13889 7536 13923
rect 7478 13883 7536 13889
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13920 7803 13923
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7791 13892 7849 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 8104 13923 8162 13929
rect 8104 13889 8116 13923
rect 8150 13920 8162 13923
rect 8386 13920 8392 13932
rect 8150 13892 8392 13920
rect 8150 13889 8162 13892
rect 8104 13883 8162 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 9968 13929 9996 14016
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 14366 13988 14372 14000
rect 10100 13960 14372 13988
rect 10100 13948 10106 13960
rect 14366 13948 14372 13960
rect 14424 13948 14430 14000
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 17681 13991 17739 13997
rect 17681 13988 17693 13991
rect 16448 13960 17693 13988
rect 16448 13948 16454 13960
rect 17681 13957 17693 13960
rect 17727 13957 17739 13991
rect 18046 13988 18052 14000
rect 18007 13960 18052 13988
rect 17681 13951 17739 13957
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 10220 13923 10278 13929
rect 10220 13889 10232 13923
rect 10266 13920 10278 13923
rect 10502 13920 10508 13932
rect 10266 13892 10508 13920
rect 10266 13889 10278 13892
rect 10220 13883 10278 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11020 13892 11529 13920
rect 11020 13880 11026 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11773 13923 11831 13929
rect 11773 13920 11785 13923
rect 11517 13883 11575 13889
rect 11624 13892 11785 13920
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13821 5963 13855
rect 9490 13852 9496 13864
rect 5905 13815 5963 13821
rect 9232 13824 9496 13852
rect 3050 13716 3056 13728
rect 3011 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5920 13716 5948 13815
rect 6362 13784 6368 13796
rect 6323 13756 6368 13784
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 9232 13793 9260 13824
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 11624 13852 11652 13892
rect 11773 13889 11785 13892
rect 11819 13920 11831 13923
rect 12158 13920 12164 13932
rect 11819 13892 12164 13920
rect 11819 13889 11831 13892
rect 11773 13883 11831 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 17696 13920 17724 13951
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 18616 13988 18644 14016
rect 19702 13988 19708 14000
rect 18616 13960 19708 13988
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 20806 13988 20812 14000
rect 20732 13960 20812 13988
rect 18690 13920 18696 13932
rect 17696 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 19153 13923 19211 13929
rect 19153 13920 19165 13923
rect 18984 13892 19165 13920
rect 18984 13864 19012 13892
rect 19153 13889 19165 13892
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 20732 13929 20760 13960
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19484 13892 20085 13920
rect 19484 13880 19490 13892
rect 20073 13889 20085 13892
rect 20119 13920 20131 13923
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20119 13892 20729 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 20717 13883 20775 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 11296 13824 11652 13852
rect 11296 13812 11302 13824
rect 12894 13812 12900 13864
rect 12952 13852 12958 13864
rect 17586 13852 17592 13864
rect 12952 13824 17592 13852
rect 12952 13812 12958 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 18966 13852 18972 13864
rect 18927 13824 18972 13852
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 20438 13852 20444 13864
rect 19659 13824 20444 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 21100 13852 21128 13883
rect 21266 13852 21272 13864
rect 21100 13824 21272 13852
rect 20809 13815 20867 13821
rect 9217 13787 9275 13793
rect 9217 13753 9229 13787
rect 9263 13753 9275 13787
rect 9217 13747 9275 13753
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 12989 13787 13047 13793
rect 12989 13784 13001 13787
rect 12860 13756 13001 13784
rect 12860 13744 12866 13756
rect 12989 13753 13001 13756
rect 13035 13753 13047 13787
rect 12989 13747 13047 13753
rect 17770 13744 17776 13796
rect 17828 13784 17834 13796
rect 20622 13784 20628 13796
rect 17828 13756 20628 13784
rect 17828 13744 17834 13756
rect 20622 13744 20628 13756
rect 20680 13784 20686 13796
rect 20824 13784 20852 13815
rect 21266 13812 21272 13824
rect 21324 13852 21330 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 21324 13824 21465 13852
rect 21324 13812 21330 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 20680 13756 20852 13784
rect 20680 13744 20686 13756
rect 12894 13716 12900 13728
rect 5224 13688 5948 13716
rect 12855 13688 12900 13716
rect 5224 13676 5230 13688
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18690 13716 18696 13728
rect 18104 13688 18696 13716
rect 18104 13676 18110 13688
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 7558 13512 7564 13524
rect 5132 13484 7564 13512
rect 5132 13472 5138 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8570 13512 8576 13524
rect 8531 13484 8576 13512
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10965 13515 11023 13521
rect 10965 13512 10977 13515
rect 10008 13484 10977 13512
rect 10008 13472 10014 13484
rect 10965 13481 10977 13484
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15746 13512 15752 13524
rect 15335 13484 15752 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 3142 13444 3148 13456
rect 2832 13416 3148 13444
rect 2832 13404 2838 13416
rect 3142 13404 3148 13416
rect 3200 13404 3206 13456
rect 6181 13447 6239 13453
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 6822 13444 6828 13456
rect 6227 13416 6828 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8588 13376 8616 13472
rect 10980 13388 11008 13475
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 17221 13515 17279 13521
rect 17221 13512 17233 13515
rect 17184 13484 17233 13512
rect 17184 13472 17190 13484
rect 17221 13481 17233 13484
rect 17267 13481 17279 13515
rect 17221 13475 17279 13481
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17770 13512 17776 13524
rect 17368 13484 17776 13512
rect 17368 13472 17374 13484
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19058 13512 19064 13524
rect 19015 13484 19064 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 20036 13484 20085 13512
rect 20036 13472 20042 13484
rect 20073 13481 20085 13484
rect 20119 13481 20131 13515
rect 20073 13475 20131 13481
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 12710 13444 12716 13456
rect 12575 13416 12716 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 12986 13404 12992 13456
rect 13044 13444 13050 13456
rect 18046 13444 18052 13456
rect 13044 13416 18052 13444
rect 13044 13404 13050 13416
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18141 13447 18199 13453
rect 18141 13413 18153 13447
rect 18187 13444 18199 13447
rect 18187 13416 18460 13444
rect 18187 13413 18199 13416
rect 18141 13407 18199 13413
rect 10962 13376 10968 13388
rect 8343 13348 8616 13376
rect 10875 13348 10968 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 10962 13336 10968 13348
rect 11020 13376 11026 13388
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 11020 13348 11161 13376
rect 11020 13336 11026 13348
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 12216 13348 15485 13376
rect 12216 13336 12222 13348
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 15746 13376 15752 13388
rect 15703 13348 15752 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16574 13376 16580 13388
rect 16535 13348 16580 13376
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 3142 13268 3148 13320
rect 3200 13308 3206 13320
rect 3878 13308 3884 13320
rect 3200 13280 3884 13308
rect 3200 13268 3206 13280
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 8041 13311 8099 13317
rect 4847 13280 5212 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5184 13252 5212 13280
rect 8041 13277 8053 13311
rect 8087 13308 8099 13311
rect 8481 13311 8539 13317
rect 8481 13308 8493 13311
rect 8087 13280 8493 13308
rect 8087 13277 8099 13280
rect 8041 13271 8099 13277
rect 8481 13277 8493 13280
rect 8527 13308 8539 13311
rect 9306 13308 9312 13320
rect 8527 13280 9312 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 11416 13311 11474 13317
rect 11416 13277 11428 13311
rect 11462 13308 11474 13311
rect 12250 13308 12256 13320
rect 11462 13280 12256 13308
rect 11462 13277 11474 13280
rect 11416 13271 11474 13277
rect 12250 13268 12256 13280
rect 12308 13308 12314 13320
rect 12618 13308 12624 13320
rect 12308 13280 12624 13308
rect 12308 13268 12314 13280
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16298 13308 16304 13320
rect 15896 13280 16304 13308
rect 15896 13268 15902 13280
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 17402 13308 17408 13320
rect 16807 13280 17408 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 5068 13243 5126 13249
rect 5068 13209 5080 13243
rect 5114 13209 5126 13243
rect 5068 13203 5126 13209
rect 5092 13172 5120 13203
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 6273 13243 6331 13249
rect 6273 13240 6285 13243
rect 5224 13212 6285 13240
rect 5224 13200 5230 13212
rect 6273 13209 6285 13212
rect 6319 13240 6331 13243
rect 6457 13243 6515 13249
rect 6457 13240 6469 13243
rect 6319 13212 6469 13240
rect 6319 13209 6331 13212
rect 6273 13203 6331 13209
rect 6457 13209 6469 13212
rect 6503 13240 6515 13243
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 6503 13212 6745 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 9582 13240 9588 13252
rect 6733 13203 6791 13209
rect 6932 13212 9588 13240
rect 5626 13172 5632 13184
rect 5092 13144 5632 13172
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 6932 13181 6960 13212
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 17512 13240 17540 13339
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 18325 13379 18383 13385
rect 18325 13376 18337 13379
rect 17828 13348 18337 13376
rect 17828 13336 17834 13348
rect 18325 13345 18337 13348
rect 18371 13345 18383 13379
rect 18432 13376 18460 13416
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 19245 13447 19303 13453
rect 19245 13444 19257 13447
rect 18564 13416 19257 13444
rect 18564 13404 18570 13416
rect 19245 13413 19257 13416
rect 19291 13413 19303 13447
rect 19245 13407 19303 13413
rect 19518 13376 19524 13388
rect 18432 13348 19524 13376
rect 18325 13339 18383 13345
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19794 13376 19800 13388
rect 19755 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 20438 13336 20444 13388
rect 20496 13336 20502 13388
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20588 13348 20637 13376
rect 20588 13336 20594 13348
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 20456 13308 20484 13336
rect 18647 13280 20484 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 12032 13212 17540 13240
rect 18509 13243 18567 13249
rect 12032 13200 12038 13212
rect 18509 13209 18521 13243
rect 18555 13240 18567 13243
rect 18690 13240 18696 13252
rect 18555 13212 18696 13240
rect 18555 13209 18567 13212
rect 18509 13203 18567 13209
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 20441 13243 20499 13249
rect 20441 13209 20453 13243
rect 20487 13240 20499 13243
rect 20806 13240 20812 13252
rect 20487 13212 20812 13240
rect 20487 13209 20499 13212
rect 20441 13203 20499 13209
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13141 6975 13175
rect 6917 13135 6975 13141
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 12526 13172 12532 13184
rect 8720 13144 12532 13172
rect 8720 13132 8726 13144
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 15749 13175 15807 13181
rect 15749 13141 15761 13175
rect 15795 13172 15807 13175
rect 15838 13172 15844 13184
rect 15795 13144 15844 13172
rect 15795 13141 15807 13144
rect 15749 13135 15807 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 16114 13172 16120 13184
rect 16075 13144 16120 13172
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16298 13172 16304 13184
rect 16259 13144 16304 13172
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17310 13172 17316 13184
rect 16899 13144 17316 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17460 13144 17693 13172
rect 17460 13132 17466 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 17770 13132 17776 13184
rect 17828 13172 17834 13184
rect 17828 13144 17873 13172
rect 17828 13132 17834 13144
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19484 13144 19625 13172
rect 19484 13132 19490 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 19705 13175 19763 13181
rect 19705 13141 19717 13175
rect 19751 13172 19763 13175
rect 20254 13172 20260 13184
rect 19751 13144 20260 13172
rect 19751 13141 19763 13144
rect 19705 13135 19763 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20530 13132 20536 13184
rect 20588 13172 20594 13184
rect 20588 13144 20633 13172
rect 20588 13132 20594 13144
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 6730 12968 6736 12980
rect 2648 12940 6736 12968
rect 2648 12928 2654 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9585 12971 9643 12977
rect 9585 12937 9597 12971
rect 9631 12968 9643 12971
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9631 12940 9781 12968
rect 9631 12937 9643 12940
rect 9585 12931 9643 12937
rect 9769 12937 9781 12940
rect 9815 12968 9827 12971
rect 9950 12968 9956 12980
rect 9815 12940 9956 12968
rect 9815 12937 9827 12940
rect 9769 12931 9827 12937
rect 5292 12903 5350 12909
rect 5292 12869 5304 12903
rect 5338 12900 5350 12903
rect 7006 12900 7012 12912
rect 5338 12872 7012 12900
rect 5338 12869 5350 12872
rect 5292 12863 5350 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 4982 12832 4988 12844
rect 2096 12804 4988 12832
rect 2096 12792 2102 12804
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 6822 12841 6828 12844
rect 6816 12832 6828 12841
rect 6783 12804 6828 12832
rect 6816 12795 6828 12804
rect 6822 12792 6828 12795
rect 6880 12792 6886 12844
rect 9145 12835 9203 12841
rect 9145 12801 9157 12835
rect 9191 12832 9203 12835
rect 9401 12835 9459 12841
rect 9191 12804 9352 12832
rect 9191 12801 9203 12804
rect 9145 12795 9203 12801
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5537 12727 5595 12733
rect 6380 12736 6561 12764
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5552 12628 5580 12727
rect 6380 12637 6408 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 9324 12764 9352 12804
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9600 12832 9628 12931
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 11054 12968 11060 12980
rect 10060 12940 11060 12968
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9447 12804 9965 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10060 12764 10088 12940
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 10220 12903 10278 12909
rect 10220 12869 10232 12903
rect 10266 12900 10278 12903
rect 10870 12900 10876 12912
rect 10266 12872 10876 12900
rect 10266 12869 10278 12872
rect 10220 12863 10278 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 11348 12900 11376 12931
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 12584 12940 13369 12968
rect 12584 12928 12590 12940
rect 13357 12937 13369 12940
rect 13403 12968 13415 12971
rect 13630 12968 13636 12980
rect 13403 12940 13636 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13630 12928 13636 12940
rect 13688 12968 13694 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13688 12940 14013 12968
rect 13688 12928 13694 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 14001 12931 14059 12937
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 14507 12940 16957 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 16945 12931 17003 12937
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17552 12940 17597 12968
rect 17552 12928 17558 12940
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 17828 12940 18613 12968
rect 17828 12928 17834 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 18601 12931 18659 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20254 12968 20260 12980
rect 20215 12940 20260 12968
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 20625 12971 20683 12977
rect 20625 12937 20637 12971
rect 20671 12968 20683 12971
rect 21174 12968 21180 12980
rect 20671 12940 21180 12968
rect 20671 12937 20683 12940
rect 20625 12931 20683 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 11784 12903 11842 12909
rect 11784 12900 11796 12903
rect 11020 12872 11100 12900
rect 11348 12872 11796 12900
rect 11020 12860 11026 12872
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11072 12832 11100 12872
rect 11784 12869 11796 12872
rect 11830 12900 11842 12903
rect 13538 12900 13544 12912
rect 11830 12872 13400 12900
rect 13499 12872 13544 12900
rect 11830 12869 11842 12872
rect 11784 12863 11842 12869
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10744 12804 11008 12832
rect 11072 12804 11529 12832
rect 10744 12792 10750 12804
rect 9324 12736 10088 12764
rect 10980 12764 11008 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 13372 12832 13400 12872
rect 13538 12860 13544 12872
rect 13596 12900 13602 12912
rect 14093 12903 14151 12909
rect 14093 12900 14105 12903
rect 13596 12872 14105 12900
rect 13596 12860 13602 12872
rect 14093 12869 14105 12872
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 15562 12860 15568 12912
rect 15620 12900 15626 12912
rect 15620 12872 15976 12900
rect 15620 12860 15626 12872
rect 15838 12832 15844 12844
rect 11517 12795 11575 12801
rect 11624 12804 13308 12832
rect 13372 12804 13952 12832
rect 15799 12804 15844 12832
rect 11624 12764 11652 12804
rect 10980 12736 11652 12764
rect 13280 12764 13308 12804
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13280 12736 13829 12764
rect 6549 12727 6607 12733
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13924 12764 13952 12804
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 15948 12832 15976 12872
rect 16114 12860 16120 12912
rect 16172 12900 16178 12912
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 16172 12872 17969 12900
rect 16172 12860 16178 12872
rect 17957 12869 17969 12872
rect 18003 12869 18015 12903
rect 17957 12863 18015 12869
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 18104 12872 19932 12900
rect 18104 12860 18110 12872
rect 17037 12835 17095 12841
rect 15948 12804 16896 12832
rect 15746 12764 15752 12776
rect 13924 12736 15752 12764
rect 13817 12727 13875 12733
rect 7929 12699 7987 12705
rect 7929 12665 7941 12699
rect 7975 12696 7987 12699
rect 7975 12668 8524 12696
rect 7975 12665 7987 12668
rect 7929 12659 7987 12665
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5224 12600 5641 12628
rect 5224 12588 5230 12600
rect 5629 12597 5641 12600
rect 5675 12628 5687 12631
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 5675 12600 6101 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 6089 12597 6101 12600
rect 6135 12628 6147 12631
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 6135 12600 6377 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 8496 12628 8524 12668
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 12989 12699 13047 12705
rect 12989 12696 13001 12699
rect 12860 12668 13001 12696
rect 12860 12656 12866 12668
rect 12989 12665 13001 12668
rect 13035 12665 13047 12699
rect 13832 12696 13860 12727
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16206 12764 16212 12776
rect 16163 12736 16212 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16868 12773 16896 12804
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17770 12832 17776 12844
rect 17083 12804 17776 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 17911 12804 18337 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 18414 12832 18420 12844
rect 18371 12804 18420 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18966 12832 18972 12844
rect 18927 12804 18972 12832
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19794 12832 19800 12844
rect 19168 12804 19380 12832
rect 19755 12804 19800 12832
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 16899 12736 17080 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 16942 12696 16948 12708
rect 13832 12668 16948 12696
rect 12989 12659 13047 12665
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 11238 12628 11244 12640
rect 8496 12600 11244 12628
rect 6365 12591 6423 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 12894 12628 12900 12640
rect 12855 12600 12900 12628
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 15013 12631 15071 12637
rect 15013 12597 15025 12631
rect 15059 12628 15071 12631
rect 15654 12628 15660 12640
rect 15059 12600 15660 12628
rect 15059 12597 15071 12600
rect 15013 12591 15071 12597
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 17052 12628 17080 12736
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 18046 12764 18052 12776
rect 17644 12736 18052 12764
rect 17644 12724 17650 12736
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 19058 12764 19064 12776
rect 19019 12736 19064 12764
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 17862 12656 17868 12708
rect 17920 12696 17926 12708
rect 19168 12696 19196 12804
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 17920 12668 19196 12696
rect 17920 12656 17926 12668
rect 19260 12628 19288 12727
rect 19352 12696 19380 12804
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 19904 12832 19932 12872
rect 19904 12804 20852 12832
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 19996 12773 20024 12804
rect 20824 12773 20852 12804
rect 19889 12767 19947 12773
rect 19889 12764 19901 12767
rect 19576 12736 19901 12764
rect 19576 12724 19582 12736
rect 19889 12733 19901 12736
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12733 20039 12767
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 19981 12727 20039 12733
rect 20088 12736 20729 12764
rect 20088 12696 20116 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 19352 12668 20116 12696
rect 17052 12600 19288 12628
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20404 12600 21281 12628
rect 20404 12588 20410 12600
rect 21269 12597 21281 12600
rect 21315 12597 21327 12631
rect 21269 12591 21327 12597
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3476 12396 9904 12424
rect 3476 12384 3482 12396
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 5905 12359 5963 12365
rect 5905 12356 5917 12359
rect 5776 12328 5917 12356
rect 5776 12316 5782 12328
rect 5905 12325 5917 12328
rect 5951 12325 5963 12359
rect 9876 12356 9904 12396
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 11020 12396 11161 12424
rect 11020 12384 11026 12396
rect 11149 12393 11161 12396
rect 11195 12393 11207 12427
rect 14093 12427 14151 12433
rect 11149 12387 11207 12393
rect 11256 12396 12848 12424
rect 11256 12356 11284 12396
rect 9876 12328 11284 12356
rect 12820 12356 12848 12396
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14274 12424 14280 12436
rect 14139 12396 14280 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14792 12396 14933 12424
rect 14792 12384 14798 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 14921 12387 14979 12393
rect 14458 12356 14464 12368
rect 12820 12328 14464 12356
rect 5905 12319 5963 12325
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 12713 12291 12771 12297
rect 10008 12260 11100 12288
rect 10008 12248 10014 12260
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 5166 12220 5172 12232
rect 4203 12192 5172 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 5166 12180 5172 12192
rect 5224 12220 5230 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5224 12192 5825 12220
rect 5224 12180 5230 12192
rect 5813 12189 5825 12192
rect 5859 12220 5871 12223
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 5859 12192 7297 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 7285 12189 7297 12192
rect 7331 12220 7343 12223
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7331 12192 7389 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7377 12189 7389 12192
rect 7423 12220 7435 12223
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 7423 12192 8953 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 8941 12189 8953 12192
rect 8987 12220 8999 12223
rect 10962 12220 10968 12232
rect 8987 12192 10968 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11072 12220 11100 12260
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 12802 12288 12808 12300
rect 12759 12260 12808 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 14424 12260 14657 12288
rect 14424 12248 14430 12260
rect 14645 12257 14657 12260
rect 14691 12257 14703 12291
rect 14936 12288 14964 12387
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 17862 12424 17868 12436
rect 15252 12396 15516 12424
rect 17823 12396 17868 12424
rect 15252 12384 15258 12396
rect 15488 12368 15516 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19518 12424 19524 12436
rect 19479 12396 19524 12424
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 21450 12424 21456 12436
rect 21223 12396 21456 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 15470 12316 15476 12368
rect 15528 12316 15534 12368
rect 16206 12356 16212 12368
rect 15672 12328 16212 12356
rect 15672 12297 15700 12328
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 17368 12328 17969 12356
rect 17368 12316 17374 12328
rect 17957 12325 17969 12328
rect 18003 12325 18015 12359
rect 17957 12319 18015 12325
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 22370 12356 22376 12368
rect 20312 12328 22376 12356
rect 20312 12316 20318 12328
rect 22370 12316 22376 12328
rect 22428 12316 22434 12368
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14936 12260 15669 12288
rect 14645 12251 14703 12257
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 15804 12260 17233 12288
rect 15804 12248 15810 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 17494 12288 17500 12300
rect 17451 12260 17500 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 16390 12220 16396 12232
rect 11072 12192 16396 12220
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17420 12220 17448 12251
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18509 12291 18567 12297
rect 18509 12288 18521 12291
rect 18104 12260 18521 12288
rect 18104 12248 18110 12260
rect 18509 12257 18521 12260
rect 18555 12257 18567 12291
rect 18509 12251 18567 12257
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19024 12260 19257 12288
rect 19024 12248 19030 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19794 12288 19800 12300
rect 19755 12260 19800 12288
rect 19245 12251 19303 12257
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 20622 12248 20628 12300
rect 20680 12288 20686 12300
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 20680 12260 20729 12288
rect 20680 12248 20686 12260
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 20717 12251 20775 12257
rect 17083 12192 17448 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 17736 12192 18429 12220
rect 17736 12180 17742 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 20993 12223 21051 12229
rect 20993 12220 21005 12223
rect 19576 12192 21005 12220
rect 19576 12180 19582 12192
rect 20993 12189 21005 12192
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4402 12155 4460 12161
rect 4402 12152 4414 12155
rect 4304 12124 4414 12152
rect 4304 12112 4310 12124
rect 4402 12121 4414 12124
rect 4448 12121 4460 12155
rect 4402 12115 4460 12121
rect 7018 12155 7076 12161
rect 7018 12121 7030 12155
rect 7064 12121 7076 12155
rect 7018 12115 7076 12121
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 5626 12084 5632 12096
rect 5583 12056 5632 12084
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 5626 12044 5632 12056
rect 5684 12084 5690 12096
rect 5810 12084 5816 12096
rect 5684 12056 5816 12084
rect 5684 12044 5690 12056
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7033 12084 7061 12115
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 7622 12155 7680 12161
rect 7622 12152 7634 12155
rect 7524 12124 7634 12152
rect 7524 12112 7530 12124
rect 7622 12121 7634 12124
rect 7668 12121 7680 12155
rect 7622 12115 7680 12121
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9186 12155 9244 12161
rect 9186 12152 9198 12155
rect 9088 12124 9198 12152
rect 9088 12112 9094 12124
rect 9186 12121 9198 12124
rect 9232 12121 9244 12155
rect 11054 12152 11060 12164
rect 9186 12115 9244 12121
rect 9324 12124 11060 12152
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 7033 12056 8769 12084
rect 8757 12053 8769 12056
rect 8803 12084 8815 12087
rect 9324 12084 9352 12124
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 12526 12161 12532 12164
rect 12468 12155 12532 12161
rect 12468 12121 12480 12155
rect 12514 12121 12532 12155
rect 12468 12115 12532 12121
rect 12526 12112 12532 12115
rect 12584 12112 12590 12164
rect 15473 12155 15531 12161
rect 15473 12121 15485 12155
rect 15519 12152 15531 12155
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15519 12124 15945 12152
rect 15519 12121 15531 12124
rect 15473 12115 15531 12121
rect 15933 12121 15945 12124
rect 15979 12121 15991 12155
rect 15933 12115 15991 12121
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 18874 12152 18880 12164
rect 17000 12124 18880 12152
rect 17000 12112 17006 12124
rect 18874 12112 18880 12124
rect 18932 12112 18938 12164
rect 19426 12112 19432 12164
rect 19484 12152 19490 12164
rect 20533 12155 20591 12161
rect 20533 12152 20545 12155
rect 19484 12124 20545 12152
rect 19484 12112 19490 12124
rect 20533 12121 20545 12124
rect 20579 12152 20591 12155
rect 21266 12152 21272 12164
rect 20579 12124 21272 12152
rect 20579 12121 20591 12124
rect 20533 12115 20591 12121
rect 21266 12112 21272 12124
rect 21324 12152 21330 12164
rect 21361 12155 21419 12161
rect 21361 12152 21373 12155
rect 21324 12124 21373 12152
rect 21324 12112 21330 12124
rect 21361 12121 21373 12124
rect 21407 12121 21419 12155
rect 21361 12115 21419 12121
rect 8803 12056 9352 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 9950 12084 9956 12096
rect 9548 12056 9956 12084
rect 9548 12044 9554 12056
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10321 12087 10379 12093
rect 10321 12053 10333 12087
rect 10367 12084 10379 12087
rect 10778 12084 10784 12096
rect 10367 12056 10784 12084
rect 10367 12053 10379 12056
rect 10321 12047 10379 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 11790 12084 11796 12096
rect 11379 12056 11796 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 14458 12084 14464 12096
rect 14419 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14553 12087 14611 12093
rect 14553 12053 14565 12087
rect 14599 12084 14611 12087
rect 14734 12084 14740 12096
rect 14599 12056 14740 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15378 12084 15384 12096
rect 15151 12056 15384 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 15654 12084 15660 12096
rect 15611 12056 15660 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 16080 12056 17509 12084
rect 16080 12044 16086 12056
rect 17497 12053 17509 12056
rect 17543 12084 17555 12087
rect 18046 12084 18052 12096
rect 17543 12056 18052 12084
rect 17543 12053 17555 12056
rect 17497 12047 17555 12053
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 18322 12084 18328 12096
rect 18283 12056 18328 12084
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 18785 12087 18843 12093
rect 18785 12084 18797 12087
rect 18748 12056 18797 12084
rect 18748 12044 18754 12056
rect 18785 12053 18797 12056
rect 18831 12053 18843 12087
rect 18785 12047 18843 12053
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 20622 12084 20628 12096
rect 20404 12056 20628 12084
rect 20404 12044 20410 12056
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 3050 11880 3056 11892
rect 2823 11852 3056 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 1946 11812 1952 11824
rect 1907 11784 1952 11812
rect 1946 11772 1952 11784
rect 2004 11772 2010 11824
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1762 11744 1768 11756
rect 1719 11716 1768 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1688 11676 1716 11707
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2332 11744 2360 11843
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 5534 11880 5540 11892
rect 3988 11852 5540 11880
rect 2682 11744 2688 11756
rect 2271 11716 2360 11744
rect 2643 11716 2688 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 2961 11679 3019 11685
rect 1688 11648 2912 11676
rect 1489 11611 1547 11617
rect 1489 11577 1501 11611
rect 1535 11608 1547 11611
rect 2884 11608 2912 11648
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3988 11676 4016 11852
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 8662 11880 8668 11892
rect 5644 11852 8668 11880
rect 4608 11815 4666 11821
rect 4608 11781 4620 11815
rect 4654 11812 4666 11815
rect 5644 11812 5672 11852
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9180 11852 10180 11880
rect 9180 11840 9186 11852
rect 4654 11784 5672 11812
rect 5905 11815 5963 11821
rect 4654 11781 4666 11784
rect 4608 11775 4666 11781
rect 5905 11781 5917 11815
rect 5951 11812 5963 11815
rect 6089 11815 6147 11821
rect 6089 11812 6101 11815
rect 5951 11784 6101 11812
rect 5951 11781 5963 11784
rect 5905 11775 5963 11781
rect 6089 11781 6101 11784
rect 6135 11812 6147 11815
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 6135 11784 6469 11812
rect 6135 11781 6147 11784
rect 6089 11775 6147 11781
rect 6457 11781 6469 11784
rect 6503 11812 6515 11815
rect 7285 11815 7343 11821
rect 7285 11812 7297 11815
rect 6503 11784 7297 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 7285 11781 7297 11784
rect 7331 11812 7343 11815
rect 7469 11815 7527 11821
rect 7469 11812 7481 11815
rect 7331 11784 7481 11812
rect 7331 11781 7343 11784
rect 7285 11775 7343 11781
rect 7469 11781 7481 11784
rect 7515 11812 7527 11815
rect 8389 11815 8447 11821
rect 8389 11812 8401 11815
rect 7515 11784 8401 11812
rect 7515 11781 7527 11784
rect 7469 11775 7527 11781
rect 8389 11781 8401 11784
rect 8435 11812 8447 11815
rect 8573 11815 8631 11821
rect 8573 11812 8585 11815
rect 8435 11784 8585 11812
rect 8435 11781 8447 11784
rect 8389 11775 8447 11781
rect 8573 11781 8585 11784
rect 8619 11812 8631 11815
rect 10152 11812 10180 11852
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 11241 11883 11299 11889
rect 11241 11880 11253 11883
rect 11020 11852 11253 11880
rect 11020 11840 11026 11852
rect 11241 11849 11253 11852
rect 11287 11849 11299 11883
rect 13538 11880 13544 11892
rect 11241 11843 11299 11849
rect 11440 11852 13400 11880
rect 13499 11852 13544 11880
rect 11440 11812 11468 11852
rect 12158 11812 12164 11824
rect 8619 11784 10088 11812
rect 10152 11784 11468 11812
rect 11624 11784 12164 11812
rect 8619 11781 8631 11784
rect 8573 11775 8631 11781
rect 7834 11744 7840 11756
rect 3007 11648 4016 11676
rect 4172 11716 7840 11744
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 4172 11608 4200 11716
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8478 11744 8484 11756
rect 8251 11716 8484 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8478 11704 8484 11716
rect 8536 11744 8542 11756
rect 9490 11744 9496 11756
rect 8536 11716 9496 11744
rect 8536 11704 8542 11716
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9766 11744 9772 11756
rect 9824 11753 9830 11756
rect 10060 11753 10088 11784
rect 9824 11747 9847 11753
rect 9699 11716 9772 11744
rect 9766 11704 9772 11716
rect 9835 11744 9847 11747
rect 10045 11747 10103 11753
rect 9835 11716 9996 11744
rect 9835 11713 9847 11716
rect 9824 11707 9847 11713
rect 9824 11704 9830 11707
rect 4338 11676 4344 11688
rect 4299 11648 4344 11676
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 9968 11676 9996 11716
rect 10045 11713 10057 11747
rect 10091 11744 10103 11747
rect 10962 11744 10968 11756
rect 10091 11716 10968 11744
rect 10091 11713 10103 11716
rect 10045 11707 10103 11713
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11020 11716 11529 11744
rect 11020 11704 11026 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 9968 11648 10241 11676
rect 10229 11645 10241 11648
rect 10275 11676 10287 11679
rect 11624 11676 11652 11784
rect 12158 11772 12164 11784
rect 12216 11812 12222 11824
rect 12989 11815 13047 11821
rect 12989 11812 13001 11815
rect 12216 11784 13001 11812
rect 12216 11772 12222 11784
rect 12989 11781 13001 11784
rect 13035 11781 13047 11815
rect 13372 11812 13400 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 15010 11880 15016 11892
rect 14971 11852 15016 11880
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 16390 11840 16396 11892
rect 16448 11880 16454 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16448 11852 16681 11880
rect 16448 11840 16454 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 16669 11843 16727 11849
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11849 17003 11883
rect 16945 11843 17003 11849
rect 13814 11812 13820 11824
rect 13372 11784 13820 11812
rect 12989 11775 13047 11781
rect 11790 11753 11796 11756
rect 11784 11744 11796 11753
rect 11751 11716 11796 11744
rect 11784 11707 11796 11716
rect 11848 11744 11854 11756
rect 12710 11744 12716 11756
rect 11848 11716 12716 11744
rect 11790 11704 11796 11707
rect 11848 11704 11854 11716
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 13004 11744 13032 11775
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 14369 11815 14427 11821
rect 14369 11781 14381 11815
rect 14415 11812 14427 11815
rect 16960 11812 16988 11843
rect 17218 11840 17224 11892
rect 17276 11880 17282 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17276 11852 17417 11880
rect 17276 11840 17282 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11880 18015 11883
rect 18322 11880 18328 11892
rect 18003 11852 18328 11880
rect 18003 11849 18015 11852
rect 17957 11843 18015 11849
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 19702 11880 19708 11892
rect 19663 11852 19708 11880
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20806 11880 20812 11892
rect 20767 11852 20812 11880
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 21048 11852 21097 11880
rect 21048 11840 21054 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 14415 11784 16988 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 14274 11744 14280 11756
rect 13004 11716 13768 11744
rect 14235 11716 14280 11744
rect 10275 11648 11652 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 13630 11676 13636 11688
rect 12952 11648 13636 11676
rect 12952 11636 12958 11648
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13740 11685 13768 11716
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 17236 11744 17264 11840
rect 18046 11772 18052 11824
rect 18104 11812 18110 11824
rect 18690 11812 18696 11824
rect 18104 11784 18696 11812
rect 18104 11772 18110 11784
rect 18690 11772 18696 11784
rect 18748 11772 18754 11824
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 19889 11815 19947 11821
rect 19889 11812 19901 11815
rect 19852 11784 19901 11812
rect 19852 11772 19858 11784
rect 19889 11781 19901 11784
rect 19935 11812 19947 11815
rect 20254 11812 20260 11824
rect 19935 11784 20260 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 20254 11772 20260 11784
rect 20312 11812 20318 11824
rect 20349 11815 20407 11821
rect 20349 11812 20361 11815
rect 20312 11784 20361 11812
rect 20312 11772 20318 11784
rect 20349 11781 20361 11784
rect 20395 11781 20407 11815
rect 20349 11775 20407 11781
rect 20441 11815 20499 11821
rect 20441 11781 20453 11815
rect 20487 11812 20499 11815
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 20487 11784 21281 11812
rect 20487 11781 20499 11784
rect 20441 11775 20499 11781
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 21269 11775 21327 11781
rect 16531 11716 17264 11744
rect 17313 11747 17371 11753
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17954 11744 17960 11756
rect 17359 11716 17960 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11744 18659 11747
rect 19610 11744 19616 11756
rect 18647 11716 19196 11744
rect 19523 11716 19616 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11645 15531 11679
rect 15473 11639 15531 11645
rect 1535 11580 2774 11608
rect 2884 11580 4200 11608
rect 1535 11577 1547 11580
rect 1489 11571 1547 11577
rect 2746 11552 2774 11580
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 7466 11608 7472 11620
rect 5500 11580 7472 11608
rect 5500 11568 5506 11580
rect 7466 11568 7472 11580
rect 7524 11568 7530 11620
rect 11514 11608 11520 11620
rect 10244 11580 11520 11608
rect 2746 11512 2780 11552
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 5721 11543 5779 11549
rect 5721 11540 5733 11543
rect 4304 11512 5733 11540
rect 4304 11500 4310 11512
rect 5721 11509 5733 11512
rect 5767 11540 5779 11543
rect 6638 11540 6644 11552
rect 5767 11512 6644 11540
rect 5767 11509 5779 11512
rect 5721 11503 5779 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 10244 11540 10272 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 14108 11608 14136 11639
rect 12820 11580 14136 11608
rect 15488 11608 15516 11639
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 15620 11648 15665 11676
rect 15620 11636 15626 11648
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 16448 11648 17509 11676
rect 16448 11636 16454 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18104 11648 18705 11676
rect 18104 11636 18110 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18874 11676 18880 11688
rect 18835 11648 18880 11676
rect 18693 11639 18751 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 17034 11608 17040 11620
rect 15488 11580 17040 11608
rect 9088 11512 10272 11540
rect 9088 11500 9094 11512
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 12820 11540 12848 11580
rect 17034 11568 17040 11580
rect 17092 11568 17098 11620
rect 17770 11568 17776 11620
rect 17828 11608 17834 11620
rect 19168 11617 19196 11716
rect 19610 11704 19616 11716
rect 19668 11744 19674 11756
rect 20806 11744 20812 11756
rect 19668 11716 20812 11744
rect 19668 11704 19674 11716
rect 20806 11704 20812 11716
rect 20864 11744 20870 11756
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 20864 11716 20913 11744
rect 20864 11704 20870 11716
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 19702 11636 19708 11688
rect 19760 11676 19766 11688
rect 20162 11676 20168 11688
rect 19760 11648 20168 11676
rect 19760 11636 19766 11648
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 18233 11611 18291 11617
rect 18233 11608 18245 11611
rect 17828 11580 18245 11608
rect 17828 11568 17834 11580
rect 18233 11577 18245 11580
rect 18279 11577 18291 11611
rect 18233 11571 18291 11577
rect 19153 11611 19211 11617
rect 19153 11577 19165 11611
rect 19199 11608 19211 11611
rect 20254 11608 20260 11620
rect 19199 11580 20260 11608
rect 19199 11577 19211 11580
rect 19153 11571 19211 11577
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 10376 11512 12848 11540
rect 12897 11543 12955 11549
rect 10376 11500 10382 11512
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 12986 11540 12992 11552
rect 12943 11512 12992 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13170 11540 13176 11552
rect 13131 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 17494 11540 17500 11552
rect 15252 11512 17500 11540
rect 15252 11500 15258 11512
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 17678 11500 17684 11552
rect 17736 11540 17742 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17736 11512 18061 11540
rect 17736 11500 17742 11512
rect 18049 11509 18061 11512
rect 18095 11540 18107 11543
rect 19610 11540 19616 11552
rect 18095 11512 19616 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2866 11336 2872 11348
rect 2363 11308 2872 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3786 11296 3792 11348
rect 3844 11336 3850 11348
rect 8846 11336 8852 11348
rect 3844 11308 8852 11336
rect 3844 11296 3850 11308
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 8956 11308 10701 11336
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11268 2007 11271
rect 3142 11268 3148 11280
rect 1995 11240 3148 11268
rect 1995 11237 2007 11240
rect 1949 11231 2007 11237
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 7190 11268 7196 11280
rect 7151 11240 7196 11268
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 8956 11209 8984 11308
rect 10689 11305 10701 11308
rect 10735 11336 10747 11339
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10735 11308 10885 11336
rect 10735 11305 10747 11308
rect 10689 11299 10747 11305
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 10962 11336 10968 11348
rect 10919 11308 10968 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 17034 11336 17040 11348
rect 11112 11308 16436 11336
rect 16995 11308 17040 11336
rect 11112 11296 11118 11308
rect 10318 11268 10324 11280
rect 10279 11240 10324 11268
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 8941 11203 8999 11209
rect 2148 11172 2912 11200
rect 2148 11141 2176 11172
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2133 11095 2191 11101
rect 2498 11092 2504 11104
rect 2556 11132 2562 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2556 11104 2697 11132
rect 2556 11092 2562 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2884 11073 2912 11172
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 10980 11200 11008 11296
rect 12526 11268 12532 11280
rect 12487 11240 12532 11268
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12894 11268 12900 11280
rect 12855 11240 12900 11268
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 13081 11271 13139 11277
rect 13081 11237 13093 11271
rect 13127 11268 13139 11271
rect 13538 11268 13544 11280
rect 13127 11240 13544 11268
rect 13127 11237 13139 11240
rect 13081 11231 13139 11237
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 13872 11240 14657 11268
rect 13872 11228 13878 11240
rect 14645 11237 14657 11240
rect 14691 11268 14703 11271
rect 15749 11271 15807 11277
rect 14691 11240 15332 11268
rect 14691 11237 14703 11240
rect 14645 11231 14703 11237
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 10980 11172 11161 11200
rect 8941 11163 8999 11169
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 15194 11200 15200 11212
rect 12768 11172 15200 11200
rect 12768 11160 12774 11172
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15304 11209 15332 11240
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 16206 11268 16212 11280
rect 15795 11240 16212 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15470 11200 15476 11212
rect 15335 11172 15476 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15470 11160 15476 11172
rect 15528 11200 15534 11212
rect 16408 11209 16436 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 18969 11339 19027 11345
rect 18969 11336 18981 11339
rect 18288 11308 18981 11336
rect 18288 11296 18294 11308
rect 16301 11203 16359 11209
rect 16301 11200 16313 11203
rect 15528 11172 16313 11200
rect 15528 11160 15534 11172
rect 16301 11169 16313 11172
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11169 16451 11203
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 16393 11163 16451 11169
rect 16868 11172 17601 11200
rect 4338 11132 4344 11144
rect 4251 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11132 4402 11144
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 4396 11104 5825 11132
rect 4396 11092 4402 11104
rect 5813 11101 5825 11104
rect 5859 11132 5871 11135
rect 6914 11132 6920 11144
rect 5859 11104 6920 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7285 11135 7343 11141
rect 7285 11132 7297 11135
rect 6972 11104 7297 11132
rect 6972 11092 6978 11104
rect 7285 11101 7297 11104
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 9208 11135 9266 11141
rect 9208 11101 9220 11135
rect 9254 11132 9266 11135
rect 9490 11132 9496 11144
rect 9254 11104 9496 11132
rect 9254 11101 9266 11104
rect 9208 11095 9266 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 11072 11104 12020 11132
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 4246 11064 4252 11076
rect 2915 11036 4252 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4608 11067 4666 11073
rect 4608 11033 4620 11067
rect 4654 11064 4666 11067
rect 5626 11064 5632 11076
rect 4654 11036 5632 11064
rect 4654 11033 4666 11036
rect 4608 11027 4666 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 5902 11064 5908 11076
rect 5736 11036 5908 11064
rect 5736 11005 5764 11036
rect 5902 11024 5908 11036
rect 5960 11064 5966 11076
rect 6058 11067 6116 11073
rect 6058 11064 6070 11067
rect 5960 11036 6070 11064
rect 5960 11024 5966 11036
rect 6058 11033 6070 11036
rect 6104 11033 6116 11067
rect 6058 11027 6116 11033
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7530 11067 7588 11073
rect 7530 11064 7542 11067
rect 7248 11036 7542 11064
rect 7248 11024 7254 11036
rect 7530 11033 7542 11036
rect 7576 11033 7588 11067
rect 7530 11027 7588 11033
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 10686 11064 10692 11076
rect 7892 11036 10692 11064
rect 7892 11024 7898 11036
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 5721 10999 5779 11005
rect 5721 10965 5733 10999
rect 5767 10965 5779 10999
rect 5721 10959 5779 10965
rect 8665 10999 8723 11005
rect 8665 10965 8677 10999
rect 8711 10996 8723 10999
rect 9766 10996 9772 11008
rect 8711 10968 9772 10996
rect 8711 10965 8723 10968
rect 8665 10959 8723 10965
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10134 10996 10140 11008
rect 9916 10968 10140 10996
rect 9916 10956 9922 10968
rect 10134 10956 10140 10968
rect 10192 10996 10198 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10192 10968 10425 10996
rect 10192 10956 10198 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 11072 10996 11100 11104
rect 11238 11024 11244 11076
rect 11296 11064 11302 11076
rect 11416 11067 11474 11073
rect 11416 11064 11428 11067
rect 11296 11036 11428 11064
rect 11296 11024 11302 11036
rect 11416 11033 11428 11036
rect 11462 11064 11474 11067
rect 11698 11064 11704 11076
rect 11462 11036 11704 11064
rect 11462 11033 11474 11036
rect 11416 11027 11474 11033
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 10560 10968 11100 10996
rect 10560 10956 10566 10968
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11882 10996 11888 11008
rect 11204 10968 11888 10996
rect 11204 10956 11210 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 11992 10996 12020 11104
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 16022 11132 16028 11144
rect 12492 11104 16028 11132
rect 12492 11092 12498 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16868 11141 16896 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 17696 11172 18644 11200
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16172 11104 16865 11132
rect 16172 11092 16178 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 17368 11104 17509 11132
rect 17368 11092 17374 11104
rect 17497 11101 17509 11104
rect 17543 11132 17555 11135
rect 17696 11132 17724 11172
rect 17954 11132 17960 11144
rect 17543 11104 17724 11132
rect 17867 11104 17960 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 17954 11092 17960 11104
rect 18012 11132 18018 11144
rect 18506 11132 18512 11144
rect 18012 11104 18512 11132
rect 18012 11092 18018 11104
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 12124 11036 14841 11064
rect 12124 11024 12130 11036
rect 14829 11033 14841 11036
rect 14875 11064 14887 11067
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 14875 11036 15393 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15381 11033 15393 11036
rect 15427 11064 15439 11067
rect 15654 11064 15660 11076
rect 15427 11036 15660 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 15654 11024 15660 11036
rect 15712 11064 15718 11076
rect 16209 11067 16267 11073
rect 16209 11064 16221 11067
rect 15712 11036 16221 11064
rect 15712 11024 15718 11036
rect 16209 11033 16221 11036
rect 16255 11033 16267 11067
rect 16209 11027 16267 11033
rect 17405 11067 17463 11073
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 18322 11064 18328 11076
rect 17451 11036 18328 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18417 11067 18475 11073
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18616 11064 18644 11172
rect 18800 11132 18828 11308
rect 18969 11305 18981 11308
rect 19015 11305 19027 11339
rect 18969 11299 19027 11305
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19116 11308 19349 11336
rect 19116 11296 19122 11308
rect 19337 11305 19349 11308
rect 19383 11305 19395 11339
rect 19337 11299 19395 11305
rect 20165 11339 20223 11345
rect 20165 11305 20177 11339
rect 20211 11336 20223 11339
rect 20530 11336 20536 11348
rect 20211 11308 20536 11336
rect 20211 11305 20223 11308
rect 20165 11299 20223 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 19794 11228 19800 11280
rect 19852 11268 19858 11280
rect 20622 11268 20628 11280
rect 19852 11240 20628 11268
rect 19852 11228 19858 11240
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 18874 11160 18880 11212
rect 18932 11200 18938 11212
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 18932 11172 19901 11200
rect 18932 11160 18938 11172
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 20220 11172 20729 11200
rect 20220 11160 20226 11172
rect 20717 11169 20729 11172
rect 20763 11169 20775 11203
rect 20717 11163 20775 11169
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 18800 11104 19717 11132
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 20588 11104 20637 11132
rect 20588 11092 20594 11104
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 20864 11104 21281 11132
rect 20864 11092 20870 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 19058 11064 19064 11076
rect 18463 11036 19064 11064
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 13078 10996 13084 11008
rect 11992 10968 13084 10996
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 15838 10996 15844 11008
rect 15799 10968 15844 10996
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 18046 10996 18052 11008
rect 16080 10968 18052 10996
rect 16080 10956 16086 10968
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 19797 10999 19855 11005
rect 19797 10965 19809 10999
rect 19843 10996 19855 10999
rect 19978 10996 19984 11008
rect 19843 10968 19984 10996
rect 19843 10965 19855 10968
rect 19797 10959 19855 10965
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 20533 10999 20591 11005
rect 20533 10965 20545 10999
rect 20579 10996 20591 10999
rect 20806 10996 20812 11008
rect 20579 10968 20812 10996
rect 20579 10965 20591 10968
rect 20533 10959 20591 10965
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 20990 10996 20996 11008
rect 20951 10968 20996 10996
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 21450 10996 21456 11008
rect 21411 10968 21456 10996
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 10502 10792 10508 10804
rect 3936 10764 10508 10792
rect 3936 10752 3942 10764
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 13262 10792 13268 10804
rect 10836 10764 11100 10792
rect 10836 10752 10842 10764
rect 5718 10724 5724 10736
rect 4632 10696 5724 10724
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 4442 10659 4500 10665
rect 4442 10656 4454 10659
rect 3476 10628 4454 10656
rect 3476 10616 3482 10628
rect 4442 10625 4454 10628
rect 4488 10625 4500 10659
rect 4442 10619 4500 10625
rect 4632 10588 4660 10696
rect 5718 10684 5724 10696
rect 5776 10724 5782 10736
rect 7254 10727 7312 10733
rect 7254 10724 7266 10727
rect 5776 10696 7266 10724
rect 5776 10684 5782 10696
rect 7254 10693 7266 10696
rect 7300 10693 7312 10727
rect 10962 10724 10968 10736
rect 7254 10687 7312 10693
rect 8496 10696 10968 10724
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5350 10656 5356 10668
rect 4755 10628 5356 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5925 10659 5983 10665
rect 5925 10625 5937 10659
rect 5971 10656 5983 10659
rect 6822 10656 6828 10668
rect 5971 10628 6828 10656
rect 5971 10625 5983 10628
rect 5925 10619 5983 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 8496 10665 8524 10696
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8748 10659 8806 10665
rect 8748 10625 8760 10659
rect 8794 10656 8806 10659
rect 9858 10656 9864 10668
rect 8794 10628 9864 10656
rect 8794 10625 8806 10628
rect 8748 10619 8806 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 9968 10665 9996 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11072 10724 11100 10764
rect 12820 10764 13268 10792
rect 12820 10724 12848 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 13872 10764 14565 10792
rect 13872 10752 13878 10764
rect 14553 10761 14565 10764
rect 14599 10792 14611 10795
rect 14826 10792 14832 10804
rect 14599 10764 14832 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15470 10792 15476 10804
rect 15431 10764 15476 10792
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15654 10792 15660 10804
rect 15615 10764 15660 10792
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 15930 10752 15936 10804
rect 15988 10792 15994 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 15988 10764 16957 10792
rect 15988 10752 15994 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 16945 10755 17003 10761
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 19935 10764 20545 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20533 10755 20591 10761
rect 20901 10795 20959 10801
rect 20901 10761 20913 10795
rect 20947 10792 20959 10795
rect 20990 10792 20996 10804
rect 20947 10764 20996 10792
rect 20947 10761 20959 10764
rect 20901 10755 20959 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 11072 10696 12848 10724
rect 12912 10696 14412 10724
rect 10226 10665 10232 10668
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 10220 10656 10232 10665
rect 10187 10628 10232 10656
rect 9953 10619 10011 10625
rect 10220 10619 10232 10628
rect 10226 10616 10232 10619
rect 10284 10616 10290 10668
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 11146 10656 11152 10668
rect 10744 10628 11152 10656
rect 10744 10616 10750 10628
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12342 10656 12348 10668
rect 11940 10628 12348 10656
rect 11940 10616 11946 10628
rect 12342 10616 12348 10628
rect 12400 10656 12406 10668
rect 12630 10659 12688 10665
rect 12630 10656 12642 10659
rect 12400 10628 12642 10656
rect 12400 10616 12406 10628
rect 12630 10625 12642 10628
rect 12676 10625 12688 10659
rect 12630 10619 12688 10625
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 12912 10665 12940 10696
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12860 10628 12909 10656
rect 12860 10616 12866 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 14384 10665 14412 10696
rect 15562 10684 15568 10736
rect 15620 10724 15626 10736
rect 18141 10727 18199 10733
rect 15620 10696 18092 10724
rect 15620 10684 15626 10696
rect 14102 10659 14160 10665
rect 14102 10656 14114 10659
rect 13044 10628 14114 10656
rect 13044 10616 13050 10628
rect 14102 10625 14114 10628
rect 14148 10656 14160 10659
rect 14369 10659 14427 10665
rect 14148 10628 14320 10656
rect 14148 10625 14160 10628
rect 14102 10619 14160 10625
rect 6181 10591 6239 10597
rect 4632 10560 4844 10588
rect 4816 10529 4844 10560
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6227 10560 6469 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6457 10557 6469 10560
rect 6503 10588 6515 10591
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6503 10560 6653 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 6641 10557 6653 10560
rect 6687 10588 6699 10591
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 6687 10560 7021 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10489 4859 10523
rect 4801 10483 4859 10489
rect 6932 10464 6960 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 14292 10588 14320 10628
rect 14369 10625 14381 10659
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16908 10628 17049 10656
rect 16908 10616 16914 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 17954 10656 17960 10668
rect 17911 10628 17960 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18064 10656 18092 10696
rect 18141 10693 18153 10727
rect 18187 10724 18199 10727
rect 19518 10724 19524 10736
rect 18187 10696 19524 10724
rect 18187 10693 18199 10696
rect 18141 10687 18199 10693
rect 19518 10684 19524 10696
rect 19576 10684 19582 10736
rect 20162 10684 20168 10736
rect 20220 10724 20226 10736
rect 20349 10727 20407 10733
rect 20349 10724 20361 10727
rect 20220 10696 20361 10724
rect 20220 10684 20226 10696
rect 20349 10693 20361 10696
rect 20395 10693 20407 10727
rect 20349 10687 20407 10693
rect 19610 10656 19616 10668
rect 18064 10628 19616 10656
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10656 21054 10668
rect 21361 10659 21419 10665
rect 21361 10656 21373 10659
rect 21048 10628 21373 10656
rect 21048 10616 21054 10628
rect 21361 10625 21373 10628
rect 21407 10656 21419 10659
rect 22462 10656 22468 10668
rect 21407 10628 22468 10656
rect 21407 10625 21419 10628
rect 21361 10619 21419 10625
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 16482 10588 16488 10600
rect 14292 10560 16488 10588
rect 7009 10551 7067 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16632 10560 16773 10588
rect 16632 10548 16638 10560
rect 16761 10557 16773 10560
rect 16807 10588 16819 10591
rect 17770 10588 17776 10600
rect 16807 10560 17776 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 19978 10588 19984 10600
rect 19939 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 21085 10591 21143 10597
rect 20128 10560 20173 10588
rect 20128 10548 20134 10560
rect 21085 10557 21097 10591
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 17218 10520 17224 10532
rect 9548 10492 9996 10520
rect 9548 10480 9554 10492
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3329 10455 3387 10461
rect 3329 10452 3341 10455
rect 2832 10424 3341 10452
rect 2832 10412 2838 10424
rect 3329 10421 3341 10424
rect 3375 10452 3387 10455
rect 5442 10452 5448 10464
rect 3375 10424 5448 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6914 10452 6920 10464
rect 6875 10424 6920 10452
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 7800 10424 8401 10452
rect 7800 10412 7806 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 8389 10415 8447 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 9968 10452 9996 10492
rect 12912 10492 13216 10520
rect 11054 10452 11060 10464
rect 9968 10424 11060 10452
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11330 10452 11336 10464
rect 11291 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 12912 10452 12940 10492
rect 11572 10424 12940 10452
rect 11572 10412 11578 10424
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 13188 10452 13216 10492
rect 14384 10492 17224 10520
rect 14384 10452 14412 10492
rect 17218 10480 17224 10492
rect 17276 10480 17282 10532
rect 19429 10523 19487 10529
rect 19429 10489 19441 10523
rect 19475 10520 19487 10523
rect 19886 10520 19892 10532
rect 19475 10492 19892 10520
rect 19475 10489 19487 10492
rect 19429 10483 19487 10489
rect 19886 10480 19892 10492
rect 19944 10520 19950 10532
rect 21100 10520 21128 10551
rect 19944 10492 21128 10520
rect 19944 10480 19950 10492
rect 13044 10424 13089 10452
rect 13188 10424 14412 10452
rect 13044 10412 13050 10424
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 17405 10455 17463 10461
rect 14792 10424 14837 10452
rect 14792 10412 14798 10424
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 18046 10452 18052 10464
rect 17451 10424 18052 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2682 10248 2688 10260
rect 2643 10220 2688 10248
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 6914 10248 6920 10260
rect 2924 10220 6408 10248
rect 6827 10220 6920 10248
rect 2924 10208 2930 10220
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3970 10112 3976 10124
rect 3375 10084 3976 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4522 10044 4528 10056
rect 4212 10016 4528 10044
rect 4212 10004 4218 10016
rect 4522 10004 4528 10016
rect 4580 10044 4586 10056
rect 4994 10047 5052 10053
rect 4994 10044 5006 10047
rect 4580 10016 5006 10044
rect 4580 10004 4586 10016
rect 4994 10013 5006 10016
rect 5040 10013 5052 10047
rect 4994 10007 5052 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5350 10044 5356 10056
rect 5307 10016 5356 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5620 10047 5678 10053
rect 5620 10044 5632 10047
rect 5552 10016 5632 10044
rect 5552 9988 5580 10016
rect 5620 10013 5632 10016
rect 5666 10044 5678 10047
rect 5994 10044 6000 10056
rect 5666 10016 6000 10044
rect 5666 10013 5678 10016
rect 5620 10007 5678 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6380 10044 6408 10220
rect 6914 10208 6920 10220
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10248 7343 10251
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 7331 10220 9045 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 6546 10140 6552 10192
rect 6604 10180 6610 10192
rect 7009 10183 7067 10189
rect 7009 10180 7021 10183
rect 6604 10152 7021 10180
rect 6604 10140 6610 10152
rect 7009 10149 7021 10152
rect 7055 10149 7067 10183
rect 7009 10143 7067 10149
rect 7392 10121 7420 10220
rect 9033 10217 9045 10220
rect 9079 10248 9091 10251
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 9079 10220 9689 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9677 10217 9689 10220
rect 9723 10248 9735 10251
rect 10962 10248 10968 10260
rect 9723 10220 10968 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10962 10208 10968 10220
rect 11020 10248 11026 10260
rect 12802 10248 12808 10260
rect 11020 10220 11192 10248
rect 12763 10220 12808 10248
rect 11020 10208 11026 10220
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 10134 10180 10140 10192
rect 8803 10152 10140 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 11164 10121 11192 10220
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 14366 10248 14372 10260
rect 13044 10220 14372 10248
rect 13044 10208 13050 10220
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15933 10251 15991 10257
rect 15933 10248 15945 10251
rect 15344 10220 15945 10248
rect 15344 10208 15350 10220
rect 15933 10217 15945 10220
rect 15979 10248 15991 10251
rect 16390 10248 16396 10260
rect 15979 10220 16396 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 16942 10208 16948 10260
rect 17000 10248 17006 10260
rect 17954 10248 17960 10260
rect 17000 10220 17045 10248
rect 17915 10220 17960 10248
rect 17000 10208 17006 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20036 10220 20269 10248
rect 20036 10208 20042 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 21082 10208 21088 10260
rect 21140 10248 21146 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 21140 10220 21281 10248
rect 21140 10208 21146 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 21269 10211 21327 10217
rect 14829 10183 14887 10189
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 17126 10180 17132 10192
rect 14875 10152 17132 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 19702 10180 19708 10192
rect 18064 10152 19708 10180
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 12802 10112 12808 10124
rect 12667 10084 12808 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 14148 10084 14197 10112
rect 14148 10072 14154 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10112 14427 10115
rect 14642 10112 14648 10124
rect 14415 10084 14648 10112
rect 14415 10081 14427 10084
rect 14369 10075 14427 10081
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 16209 10115 16267 10121
rect 16209 10112 16221 10115
rect 16172 10084 16221 10112
rect 16172 10072 16178 10084
rect 16209 10081 16221 10084
rect 16255 10081 16267 10115
rect 16390 10112 16396 10124
rect 16351 10084 16396 10112
rect 16209 10075 16267 10081
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 17494 10112 17500 10124
rect 17455 10084 17500 10112
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 10502 10044 10508 10056
rect 6380 10016 10508 10044
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 10870 10044 10876 10056
rect 10928 10053 10934 10056
rect 10928 10047 10951 10053
rect 10803 10016 10876 10044
rect 10870 10004 10876 10016
rect 10939 10044 10951 10047
rect 15194 10044 15200 10056
rect 10939 10016 15200 10044
rect 10939 10013 10951 10016
rect 10928 10007 10951 10013
rect 10928 10004 10934 10007
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 18064 10044 18092 10152
rect 19702 10140 19708 10152
rect 19760 10180 19766 10192
rect 20438 10180 20444 10192
rect 19760 10152 20444 10180
rect 19760 10140 19766 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 20530 10140 20536 10192
rect 20588 10180 20594 10192
rect 21453 10183 21511 10189
rect 21453 10180 21465 10183
rect 20588 10152 21465 10180
rect 20588 10140 20594 10152
rect 21453 10149 21465 10152
rect 21499 10149 21511 10183
rect 21453 10143 21511 10149
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18196 10084 18521 10112
rect 18196 10072 18202 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 19518 10112 19524 10124
rect 18509 10075 18567 10081
rect 18892 10084 19524 10112
rect 17359 10016 18092 10044
rect 18325 10047 18383 10053
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 18325 10013 18337 10047
rect 18371 10044 18383 10047
rect 18892 10044 18920 10084
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19610 10072 19616 10124
rect 19668 10072 19674 10124
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 20809 10115 20867 10121
rect 20809 10112 20821 10115
rect 19944 10084 20821 10112
rect 19944 10072 19950 10084
rect 20809 10081 20821 10084
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 18371 10016 18920 10044
rect 19337 10047 19395 10053
rect 18371 10013 18383 10016
rect 18325 10007 18383 10013
rect 19337 10013 19349 10047
rect 19383 10013 19395 10047
rect 19628 10044 19656 10072
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 19628 10016 20085 10044
rect 19337 10007 19395 10013
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 5534 9936 5540 9988
rect 5592 9936 5598 9988
rect 7644 9979 7702 9985
rect 5736 9948 7144 9976
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2590 9908 2596 9920
rect 2455 9880 2596 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3050 9908 3056 9920
rect 3011 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3200 9880 3245 9908
rect 3200 9868 3206 9880
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3568 9880 3893 9908
rect 3568 9868 3574 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 5736 9908 5764 9948
rect 4028 9880 5764 9908
rect 6733 9911 6791 9917
rect 4028 9868 4034 9880
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 6822 9908 6828 9920
rect 6779 9880 6828 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7116 9908 7144 9948
rect 7644 9945 7656 9979
rect 7690 9976 7702 9979
rect 10042 9976 10048 9988
rect 7690 9948 10048 9976
rect 7690 9945 7702 9948
rect 7644 9939 7702 9945
rect 10042 9936 10048 9948
rect 10100 9936 10106 9988
rect 12376 9979 12434 9985
rect 12376 9945 12388 9979
rect 12422 9976 12434 9979
rect 13078 9976 13084 9988
rect 12422 9948 13084 9976
rect 12422 9945 12434 9948
rect 12376 9939 12434 9945
rect 13078 9936 13084 9948
rect 13136 9936 13142 9988
rect 13541 9979 13599 9985
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13814 9976 13820 9988
rect 13587 9948 13820 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 13924 9948 14473 9976
rect 9490 9908 9496 9920
rect 7116 9880 9496 9908
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 10410 9908 10416 9920
rect 9815 9880 10416 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 11054 9908 11060 9920
rect 10560 9880 11060 9908
rect 10560 9868 10566 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11241 9911 11299 9917
rect 11241 9877 11253 9911
rect 11287 9908 11299 9911
rect 11790 9908 11796 9920
rect 11287 9880 11796 9908
rect 11287 9877 11299 9880
rect 11241 9871 11299 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12894 9908 12900 9920
rect 12768 9880 12900 9908
rect 12768 9868 12774 9880
rect 12894 9868 12900 9880
rect 12952 9908 12958 9920
rect 13924 9917 13952 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 14734 9936 14740 9988
rect 14792 9976 14798 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14792 9948 15393 9976
rect 14792 9936 14798 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 16485 9979 16543 9985
rect 16485 9945 16497 9979
rect 16531 9976 16543 9979
rect 16531 9948 17448 9976
rect 16531 9945 16543 9948
rect 16485 9939 16543 9945
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12952 9880 13001 9908
rect 12952 9868 12958 9880
rect 12989 9877 13001 9880
rect 13035 9908 13047 9911
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13035 9880 13461 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 13909 9911 13967 9917
rect 13909 9877 13921 9911
rect 13955 9877 13967 9911
rect 13909 9871 13967 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15286 9908 15292 9920
rect 14976 9880 15021 9908
rect 15247 9880 15292 9908
rect 14976 9868 14982 9880
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15841 9911 15899 9917
rect 15841 9877 15853 9911
rect 15887 9908 15899 9911
rect 16114 9908 16120 9920
rect 15887 9880 16120 9908
rect 15887 9877 15899 9880
rect 15841 9871 15899 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 17420 9917 17448 9948
rect 17586 9936 17592 9988
rect 17644 9976 17650 9988
rect 19352 9976 19380 10007
rect 19610 9976 19616 9988
rect 17644 9948 19380 9976
rect 19571 9948 19616 9976
rect 17644 9936 17650 9948
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 17862 9908 17868 9920
rect 17451 9880 17868 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18877 9911 18935 9917
rect 18472 9880 18517 9908
rect 18472 9868 18478 9880
rect 18877 9877 18889 9911
rect 18923 9908 18935 9911
rect 19702 9908 19708 9920
rect 18923 9880 19708 9908
rect 18923 9877 18935 9880
rect 18877 9871 18935 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 19886 9908 19892 9920
rect 19847 9880 19892 9908
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20088 9908 20116 10007
rect 20438 10004 20444 10056
rect 20496 10044 20502 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20496 10016 20729 10044
rect 20496 10004 20502 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10044 21143 10047
rect 21131 10016 21312 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20088 9880 20637 9908
rect 20625 9877 20637 9880
rect 20671 9908 20683 9911
rect 20806 9908 20812 9920
rect 20671 9880 20812 9908
rect 20671 9877 20683 9880
rect 20625 9871 20683 9877
rect 20806 9868 20812 9880
rect 20864 9908 20870 9920
rect 21284 9908 21312 10016
rect 20864 9880 21312 9908
rect 20864 9868 20870 9880
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3329 9707 3387 9713
rect 3329 9704 3341 9707
rect 3108 9676 3341 9704
rect 3108 9664 3114 9676
rect 3329 9673 3341 9676
rect 3375 9673 3387 9707
rect 4246 9704 4252 9716
rect 4207 9676 4252 9704
rect 3329 9667 3387 9673
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4430 9704 4436 9716
rect 4387 9676 4436 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 4430 9664 4436 9676
rect 4488 9704 4494 9716
rect 4706 9704 4712 9716
rect 4488 9676 4712 9704
rect 4488 9664 4494 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4893 9707 4951 9713
rect 4893 9673 4905 9707
rect 4939 9704 4951 9707
rect 5350 9704 5356 9716
rect 4939 9676 5356 9704
rect 4939 9673 4951 9676
rect 4893 9667 4951 9673
rect 5350 9664 5356 9676
rect 5408 9704 5414 9716
rect 5813 9707 5871 9713
rect 5408 9676 5672 9704
rect 5408 9664 5414 9676
rect 2961 9639 3019 9645
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 3694 9636 3700 9648
rect 3007 9608 3700 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 5534 9636 5540 9648
rect 4080 9608 5540 9636
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2740 9540 2881 9568
rect 2740 9528 2746 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1728 9472 1777 9500
rect 1728 9460 1734 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 1995 9472 2544 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2406 9432 2412 9444
rect 2367 9404 2412 9432
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 2516 9441 2544 9472
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3050 9500 3056 9512
rect 2832 9472 3056 9500
rect 2832 9460 2838 9472
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 4080 9509 4108 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 5442 9568 5448 9580
rect 4488 9540 5304 9568
rect 5403 9540 5448 9568
rect 4488 9528 4494 9540
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4614 9500 4620 9512
rect 4065 9463 4123 9469
rect 4264 9472 4620 9500
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9401 2559 9435
rect 3160 9432 3188 9463
rect 4154 9432 4160 9444
rect 3160 9404 4160 9432
rect 2501 9395 2559 9401
rect 4154 9392 4160 9404
rect 4212 9432 4218 9444
rect 4264 9432 4292 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 4982 9500 4988 9512
rect 4764 9472 4988 9500
rect 4764 9460 4770 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5166 9500 5172 9512
rect 5127 9472 5172 9500
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5276 9500 5304 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5644 9577 5672 9676
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 5994 9704 6000 9716
rect 5859 9676 6000 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 5994 9664 6000 9676
rect 6052 9704 6058 9716
rect 6546 9704 6552 9716
rect 6052 9676 6552 9704
rect 6052 9664 6058 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 9493 9707 9551 9713
rect 9493 9673 9505 9707
rect 9539 9704 9551 9707
rect 10962 9704 10968 9716
rect 9539 9676 10968 9704
rect 9539 9673 9551 9676
rect 9493 9667 9551 9673
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 5675 9540 6837 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6825 9537 6837 9540
rect 6871 9568 6883 9571
rect 6914 9568 6920 9580
rect 6871 9540 6920 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7006 9528 7012 9580
rect 7064 9528 7070 9580
rect 9600 9577 9628 9676
rect 10962 9664 10968 9676
rect 11020 9704 11026 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 11020 9676 11069 9704
rect 11020 9664 11026 9676
rect 11057 9673 11069 9676
rect 11103 9704 11115 9707
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 11103 9676 11253 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 11241 9673 11253 9676
rect 11287 9673 11299 9707
rect 11241 9667 11299 9673
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 14090 9704 14096 9716
rect 12400 9676 14096 9704
rect 12400 9664 12406 9676
rect 14090 9664 14096 9676
rect 14148 9664 14154 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14918 9704 14924 9716
rect 14231 9676 14924 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 18138 9704 18144 9716
rect 15252 9676 18144 9704
rect 15252 9664 15258 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 18693 9707 18751 9713
rect 18693 9704 18705 9707
rect 18472 9676 18705 9704
rect 18472 9664 18478 9676
rect 18693 9673 18705 9676
rect 18739 9673 18751 9707
rect 18693 9667 18751 9673
rect 19610 9664 19616 9716
rect 19668 9704 19674 9716
rect 20717 9707 20775 9713
rect 19668 9676 20668 9704
rect 19668 9664 19674 9676
rect 9858 9645 9864 9648
rect 9852 9636 9864 9645
rect 9771 9608 9864 9636
rect 9852 9599 9864 9608
rect 9916 9636 9922 9648
rect 15013 9639 15071 9645
rect 9916 9608 14320 9636
rect 9858 9596 9864 9599
rect 9916 9596 9922 9608
rect 7184 9571 7242 9577
rect 7184 9537 7196 9571
rect 7230 9568 7242 9571
rect 9585 9571 9643 9577
rect 7230 9540 9536 9568
rect 7230 9537 7242 9540
rect 7184 9531 7242 9537
rect 7024 9500 7052 9528
rect 5276 9472 7052 9500
rect 4212 9404 4292 9432
rect 4212 9392 4218 9404
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 6914 9432 6920 9444
rect 5684 9404 6920 9432
rect 5684 9392 5690 9404
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3510 9364 3516 9376
rect 2832 9336 3516 9364
rect 2832 9324 2838 9336
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4706 9364 4712 9376
rect 4667 9336 4712 9364
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8386 9364 8392 9376
rect 8343 9336 8392 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8386 9324 8392 9336
rect 8444 9364 8450 9376
rect 9122 9364 9128 9376
rect 8444 9336 9128 9364
rect 8444 9324 8450 9336
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9508 9364 9536 9540
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 12618 9528 12624 9580
rect 12676 9577 12682 9580
rect 12676 9568 12688 9577
rect 12676 9540 12721 9568
rect 12676 9531 12688 9540
rect 12676 9528 12682 9531
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12860 9540 12909 9568
rect 12860 9528 12866 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13648 9472 13921 9500
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 10520 9404 11529 9432
rect 10520 9364 10548 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 9508 9336 10548 9364
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10928 9336 10977 9364
rect 10928 9324 10934 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 11532 9364 11560 9395
rect 13648 9376 13676 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14292 9500 14320 9608
rect 15013 9605 15025 9639
rect 15059 9636 15071 9639
rect 15286 9636 15292 9648
rect 15059 9608 15292 9636
rect 15059 9605 15071 9608
rect 15013 9599 15071 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 16117 9639 16175 9645
rect 16117 9605 16129 9639
rect 16163 9636 16175 9639
rect 16942 9636 16948 9648
rect 16163 9608 16948 9636
rect 16163 9605 16175 9608
rect 16117 9599 16175 9605
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 17126 9636 17132 9648
rect 17087 9608 17132 9636
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 18233 9639 18291 9645
rect 18233 9605 18245 9639
rect 18279 9636 18291 9639
rect 18598 9636 18604 9648
rect 18279 9608 18604 9636
rect 18279 9605 18291 9608
rect 18233 9599 18291 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 19337 9639 19395 9645
rect 19337 9605 19349 9639
rect 19383 9636 19395 9639
rect 19518 9636 19524 9648
rect 19383 9608 19524 9636
rect 19383 9605 19395 9608
rect 19337 9599 19395 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 20254 9636 20260 9648
rect 20215 9608 20260 9636
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 20640 9636 20668 9676
rect 20717 9673 20729 9707
rect 20763 9704 20775 9707
rect 20806 9704 20812 9716
rect 20763 9676 20812 9704
rect 20763 9673 20775 9676
rect 20717 9667 20775 9673
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 20640 9608 21220 9636
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15194 9568 15200 9580
rect 14783 9540 15200 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15194 9528 15200 9540
rect 15252 9568 15258 9580
rect 15470 9568 15476 9580
rect 15252 9540 15476 9568
rect 15252 9528 15258 9540
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17402 9568 17408 9580
rect 17083 9540 17408 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 18874 9568 18880 9580
rect 18371 9540 18880 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 20070 9568 20076 9580
rect 19352 9540 20076 9568
rect 16390 9500 16396 9512
rect 14292 9472 14964 9500
rect 16351 9472 16396 9500
rect 14093 9463 14151 9469
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14108 9432 14136 9463
rect 13780 9404 14136 9432
rect 14553 9435 14611 9441
rect 13780 9392 13786 9404
rect 14553 9401 14565 9435
rect 14599 9432 14611 9435
rect 14826 9432 14832 9444
rect 14599 9404 14832 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 14936 9432 14964 9472
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 17218 9500 17224 9512
rect 17179 9472 17224 9500
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 17328 9472 18153 9500
rect 17328 9432 17356 9472
rect 18141 9469 18153 9472
rect 18187 9500 18199 9503
rect 19352 9500 19380 9540
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20530 9568 20536 9580
rect 20211 9540 20536 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 21192 9577 21220 9608
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20680 9540 20821 9568
rect 20680 9528 20686 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 18187 9472 19380 9500
rect 18187 9469 18199 9472
rect 18141 9463 18199 9469
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19484 9472 19529 9500
rect 19484 9460 19490 9472
rect 19610 9460 19616 9512
rect 19668 9500 19674 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 19668 9472 20361 9500
rect 19668 9460 19674 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 14936 9404 17356 9432
rect 17402 9392 17408 9444
rect 17460 9432 17466 9444
rect 19797 9435 19855 9441
rect 19797 9432 19809 9435
rect 17460 9404 19809 9432
rect 17460 9392 17466 9404
rect 19797 9401 19809 9404
rect 19843 9401 19855 9435
rect 19797 9395 19855 9401
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 20993 9435 21051 9441
rect 20993 9432 21005 9435
rect 20956 9404 21005 9432
rect 20956 9392 20962 9404
rect 20993 9401 21005 9404
rect 21039 9401 21051 9435
rect 21358 9432 21364 9444
rect 21319 9404 21364 9432
rect 20993 9395 21051 9401
rect 21358 9392 21364 9404
rect 21416 9392 21422 9444
rect 13446 9364 13452 9376
rect 11532 9336 13452 9364
rect 10965 9327 11023 9333
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 13630 9364 13636 9376
rect 13591 9336 13636 9364
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16390 9324 16396 9376
rect 16448 9364 16454 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16448 9336 16681 9364
rect 16448 9324 16454 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16669 9327 16727 9333
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17586 9364 17592 9376
rect 16908 9336 17592 9364
rect 16908 9324 16914 9336
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 17862 9364 17868 9376
rect 17823 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 18785 9367 18843 9373
rect 18785 9364 18797 9367
rect 18656 9336 18797 9364
rect 18656 9324 18662 9336
rect 18785 9333 18797 9336
rect 18831 9333 18843 9367
rect 18966 9364 18972 9376
rect 18927 9336 18972 9364
rect 18785 9327 18843 9333
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1912 9132 1961 9160
rect 1912 9120 1918 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 1949 9123 2007 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3326 9160 3332 9172
rect 2823 9132 3332 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 5074 9160 5080 9172
rect 4304 9132 5080 9160
rect 4304 9120 4310 9132
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5442 9160 5448 9172
rect 5307 9132 5448 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 13630 9160 13636 9172
rect 7432 9132 13636 9160
rect 7432 9120 7438 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 13964 9132 14381 9160
rect 13964 9120 13970 9132
rect 14369 9129 14381 9132
rect 14415 9160 14427 9163
rect 15930 9160 15936 9172
rect 14415 9132 15936 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16850 9160 16856 9172
rect 16811 9132 16856 9160
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 18414 9160 18420 9172
rect 17052 9132 18420 9160
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 9674 9092 9680 9104
rect 4028 9064 9680 9092
rect 4028 9052 4034 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10284 9064 16252 9092
rect 10284 9052 10290 9064
rect 5166 9024 5172 9036
rect 2148 8996 5172 9024
rect 2148 8965 2176 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5776 8996 5825 9024
rect 5776 8984 5782 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 6546 9024 6552 9036
rect 6507 8996 6552 9024
rect 5813 8987 5871 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 9024 6791 9027
rect 6822 9024 6828 9036
rect 6779 8996 6828 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 6972 8996 7481 9024
rect 6972 8984 6978 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12584 8996 12817 9024
rect 12584 8984 12590 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 16224 9033 16252 9064
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 17052 9092 17080 9132
rect 18414 9120 18420 9132
rect 18472 9120 18478 9172
rect 20070 9120 20076 9172
rect 20128 9160 20134 9172
rect 20254 9160 20260 9172
rect 20128 9132 20260 9160
rect 20128 9120 20134 9132
rect 20254 9120 20260 9132
rect 20312 9160 20318 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20312 9132 21281 9160
rect 20312 9120 20318 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 19610 9092 19616 9104
rect 16540 9064 17080 9092
rect 17144 9064 19616 9092
rect 16540 9052 16546 9064
rect 16209 9027 16267 9033
rect 14332 8996 16160 9024
rect 14332 8984 14338 8996
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2516 8888 2544 8919
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 2648 8928 2693 8956
rect 2648 8916 2654 8928
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 4764 8928 6469 8956
rect 4764 8916 4770 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 6457 8919 6515 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 13354 8956 13360 8968
rect 12768 8928 13360 8956
rect 12768 8916 12774 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 15654 8956 15660 8968
rect 13740 8928 15660 8956
rect 3326 8888 3332 8900
rect 2516 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 3510 8848 3516 8900
rect 3568 8888 3574 8900
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 3568 8860 7297 8888
rect 3568 8848 3574 8860
rect 7285 8857 7297 8860
rect 7331 8888 7343 8891
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7331 8860 7757 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 7745 8857 7757 8860
rect 7791 8888 7803 8891
rect 13081 8891 13139 8897
rect 7791 8860 12434 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4430 8820 4436 8832
rect 4019 8792 4436 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 4982 8820 4988 8832
rect 4939 8792 4988 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5626 8820 5632 8832
rect 5587 8792 5632 8820
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8820 5779 8823
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5767 8792 6101 8820
rect 5767 8789 5779 8792
rect 5721 8783 5779 8789
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 6089 8783 6147 8789
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 6604 8792 6929 8820
rect 6604 8780 6610 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 12406 8820 12434 8860
rect 13081 8857 13093 8891
rect 13127 8888 13139 8891
rect 13541 8891 13599 8897
rect 13541 8888 13553 8891
rect 13127 8860 13553 8888
rect 13127 8857 13139 8860
rect 13081 8851 13139 8857
rect 13541 8857 13553 8860
rect 13587 8857 13599 8891
rect 13541 8851 13599 8857
rect 12802 8820 12808 8832
rect 12406 8792 12808 8820
rect 6917 8783 6975 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 12986 8820 12992 8832
rect 12947 8792 12992 8820
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13449 8823 13507 8829
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 13740 8820 13768 8928
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 16132 8956 16160 8996
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16390 9024 16396 9036
rect 16351 8996 16396 9024
rect 16209 8987 16267 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 17144 8956 17172 9064
rect 19610 9052 19616 9064
rect 19668 9092 19674 9104
rect 19668 9064 20116 9092
rect 19668 9052 19674 9064
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 17276 8996 18337 9024
rect 17276 8984 17282 8996
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18656 8996 19073 9024
rect 18656 8984 18662 8996
rect 19061 8993 19073 8996
rect 19107 8993 19119 9027
rect 19061 8987 19119 8993
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19518 9024 19524 9036
rect 19475 8996 19524 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 16132 8928 17172 8956
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 18966 8956 18972 8968
rect 18187 8928 18972 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19076 8956 19104 8987
rect 19518 8984 19524 8996
rect 19576 8984 19582 9036
rect 20088 9033 20116 9064
rect 20162 9052 20168 9104
rect 20220 9092 20226 9104
rect 20346 9092 20352 9104
rect 20220 9064 20352 9092
rect 20220 9052 20226 9064
rect 20346 9052 20352 9064
rect 20404 9092 20410 9104
rect 21453 9095 21511 9101
rect 21453 9092 21465 9095
rect 20404 9064 21465 9092
rect 20404 9052 20410 9064
rect 21453 9061 21465 9064
rect 21499 9061 21511 9095
rect 21453 9055 21511 9061
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 8993 20131 9027
rect 20622 9024 20628 9036
rect 20073 8987 20131 8993
rect 20180 8996 20484 9024
rect 20583 8996 20628 9024
rect 19889 8959 19947 8965
rect 19889 8956 19901 8959
rect 19076 8928 19901 8956
rect 19889 8925 19901 8928
rect 19935 8956 19947 8959
rect 20180 8956 20208 8996
rect 20346 8956 20352 8968
rect 19935 8928 20208 8956
rect 20307 8928 20352 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20456 8956 20484 8996
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 20806 8956 20812 8968
rect 20456 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 13872 8860 14565 8888
rect 13872 8848 13878 8860
rect 14553 8857 14565 8860
rect 14599 8888 14611 8891
rect 15102 8888 15108 8900
rect 14599 8860 15108 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 16485 8891 16543 8897
rect 16485 8857 16497 8891
rect 16531 8857 16543 8891
rect 16485 8851 16543 8857
rect 18233 8891 18291 8897
rect 18233 8857 18245 8891
rect 18279 8888 18291 8891
rect 18279 8860 19012 8888
rect 18279 8857 18291 8860
rect 18233 8851 18291 8857
rect 14090 8820 14096 8832
rect 13495 8792 13768 8820
rect 14051 8792 14096 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 14734 8820 14740 8832
rect 14695 8792 14740 8820
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 16500 8820 16528 8851
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 16500 8792 17785 8820
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 18984 8820 19012 8860
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 21085 8891 21143 8897
rect 21085 8888 21097 8891
rect 20496 8860 21097 8888
rect 20496 8848 20502 8860
rect 21085 8857 21097 8860
rect 21131 8857 21143 8891
rect 21085 8851 21143 8857
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 18984 8792 19533 8820
rect 17773 8783 17831 8789
rect 19521 8789 19533 8792
rect 19567 8789 19579 8823
rect 19521 8783 19579 8789
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 20162 8820 20168 8832
rect 20027 8792 20168 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20588 8792 20913 8820
rect 20588 8780 20594 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1452 8588 1961 8616
rect 1452 8576 1458 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 1949 8579 2007 8585
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 3743 8588 4997 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 6086 8616 6092 8628
rect 5224 8588 5856 8616
rect 5999 8588 6092 8616
rect 5224 8576 5230 8588
rect 2317 8551 2375 8557
rect 2317 8517 2329 8551
rect 2363 8548 2375 8551
rect 3510 8548 3516 8560
rect 2363 8520 3516 8548
rect 2363 8517 2375 8520
rect 2317 8511 2375 8517
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2332 8480 2360 8511
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 4246 8548 4252 8560
rect 3651 8520 4252 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 4430 8548 4436 8560
rect 4391 8520 4436 8548
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 5718 8548 5724 8560
rect 4488 8520 5724 8548
rect 4488 8508 4494 8520
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 5828 8548 5856 8588
rect 6086 8576 6092 8588
rect 6144 8616 6150 8628
rect 7742 8616 7748 8628
rect 6144 8588 7748 8616
rect 6144 8576 6150 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 13722 8616 13728 8628
rect 11204 8588 13308 8616
rect 13683 8588 13728 8616
rect 11204 8576 11210 8588
rect 7006 8548 7012 8560
rect 5828 8520 7012 8548
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 7708 8520 12940 8548
rect 7708 8508 7714 8520
rect 4062 8480 4068 8492
rect 2179 8452 2360 8480
rect 3896 8452 4068 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 3896 8421 3924 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5132 8452 5365 8480
rect 5132 8440 5138 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5491 8452 5917 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5905 8449 5917 8452
rect 5951 8480 5963 8483
rect 12710 8480 12716 8492
rect 5951 8452 12716 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 4614 8412 4620 8424
rect 4571 8384 4620 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5166 8412 5172 8424
rect 4755 8384 5172 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5316 8384 5641 8412
rect 5316 8372 5322 8384
rect 5629 8381 5641 8384
rect 5675 8412 5687 8415
rect 6086 8412 6092 8424
rect 5675 8384 6092 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6454 8412 6460 8424
rect 6367 8384 6460 8412
rect 6454 8372 6460 8384
rect 6512 8412 6518 8424
rect 7466 8412 7472 8424
rect 6512 8384 7472 8412
rect 6512 8372 6518 8384
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 12912 8421 12940 8520
rect 13280 8421 13308 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14507 8588 14933 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 18874 8616 18880 8628
rect 18835 8588 18880 8616
rect 14921 8579 14979 8585
rect 13357 8551 13415 8557
rect 13357 8517 13369 8551
rect 13403 8548 13415 8551
rect 13906 8548 13912 8560
rect 13403 8520 13912 8548
rect 13403 8517 13415 8520
rect 13357 8511 13415 8517
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 14108 8548 14136 8579
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 20993 8619 21051 8625
rect 20993 8616 21005 8619
rect 20772 8588 21005 8616
rect 20772 8576 20778 8588
rect 20993 8585 21005 8588
rect 21039 8585 21051 8619
rect 20993 8579 21051 8585
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21634 8616 21640 8628
rect 21407 8588 21640 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 14550 8548 14556 8560
rect 14108 8520 14556 8548
rect 14550 8508 14556 8520
rect 14608 8508 14614 8560
rect 14734 8508 14740 8560
rect 14792 8548 14798 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14792 8520 15393 8548
rect 14792 8508 14798 8520
rect 15381 8517 15393 8520
rect 15427 8548 15439 8551
rect 18598 8548 18604 8560
rect 15427 8520 18604 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 18785 8551 18843 8557
rect 18785 8517 18797 8551
rect 18831 8548 18843 8551
rect 19426 8548 19432 8560
rect 18831 8520 19432 8548
rect 18831 8517 18843 8520
rect 18785 8511 18843 8517
rect 19426 8508 19432 8520
rect 19484 8548 19490 8560
rect 19886 8548 19892 8560
rect 19484 8520 19892 8548
rect 19484 8508 19490 8520
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 15289 8483 15347 8489
rect 14148 8452 14688 8480
rect 14148 8440 14154 8452
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 12943 8384 13185 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13722 8412 13728 8424
rect 13311 8384 13728 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 4065 8347 4123 8353
rect 4065 8313 4077 8347
rect 4111 8344 4123 8347
rect 4338 8344 4344 8356
rect 4111 8316 4344 8344
rect 4111 8313 4123 8316
rect 4065 8307 4123 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 13188 8344 13216 8375
rect 13722 8372 13728 8384
rect 13780 8412 13786 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 13780 8384 13829 8412
rect 13780 8372 13786 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 14550 8412 14556 8424
rect 14511 8384 14556 8412
rect 13817 8375 13875 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14660 8421 14688 8452
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15335 8452 15761 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 19150 8480 19156 8492
rect 15988 8452 19156 8480
rect 15988 8440 15994 8452
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 19978 8480 19984 8492
rect 19291 8452 19984 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20456 8452 20821 8480
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8381 14703 8415
rect 15194 8412 15200 8424
rect 14645 8375 14703 8381
rect 14752 8384 15200 8412
rect 14752 8344 14780 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 5920 8316 6500 8344
rect 13188 8316 14780 8344
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 5920 8276 5948 8316
rect 4028 8248 5948 8276
rect 6472 8276 6500 8316
rect 15102 8304 15108 8356
rect 15160 8344 15166 8356
rect 15488 8344 15516 8375
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 19058 8412 19064 8424
rect 17920 8384 19064 8412
rect 17920 8372 17926 8384
rect 19058 8372 19064 8384
rect 19116 8412 19122 8424
rect 19337 8415 19395 8421
rect 19337 8412 19349 8415
rect 19116 8384 19349 8412
rect 19116 8372 19122 8384
rect 19337 8381 19349 8384
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 15160 8316 15516 8344
rect 19352 8344 19380 8375
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19484 8384 19529 8412
rect 19484 8372 19490 8384
rect 19705 8347 19763 8353
rect 19705 8344 19717 8347
rect 19352 8316 19717 8344
rect 15160 8304 15166 8316
rect 19705 8313 19717 8316
rect 19751 8313 19763 8347
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19705 8307 19763 8313
rect 19812 8316 20085 8344
rect 13538 8276 13544 8288
rect 6472 8248 13544 8276
rect 4028 8236 4034 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 14642 8276 14648 8288
rect 13688 8248 14648 8276
rect 13688 8236 13694 8248
rect 14642 8236 14648 8248
rect 14700 8276 14706 8288
rect 18598 8276 18604 8288
rect 14700 8248 18604 8276
rect 14700 8236 14706 8248
rect 18598 8236 18604 8248
rect 18656 8276 18662 8288
rect 19812 8276 19840 8316
rect 20073 8313 20085 8316
rect 20119 8344 20131 8347
rect 20456 8344 20484 8452
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 21192 8412 21220 8443
rect 20579 8384 21220 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20119 8316 20484 8344
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 18656 8248 19840 8276
rect 18656 8236 18662 8248
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20622 8276 20628 8288
rect 20036 8248 20628 8276
rect 20036 8236 20042 8248
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2096 8044 2237 8072
rect 2096 8032 2102 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 13630 8072 13636 8084
rect 4120 8044 13636 8072
rect 4120 8032 4126 8044
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 13814 8072 13820 8084
rect 13775 8044 13820 8072
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14608 8044 14841 8072
rect 14608 8032 14614 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 18322 8072 18328 8084
rect 15243 8044 18328 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 3234 7964 3240 8016
rect 3292 8004 3298 8016
rect 14734 8004 14740 8016
rect 3292 7976 14740 8004
rect 3292 7964 3298 7976
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2590 7936 2596 7948
rect 1995 7908 2596 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 4154 7936 4160 7948
rect 2915 7908 4160 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4522 7936 4528 7948
rect 4483 7908 4528 7936
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5902 7936 5908 7948
rect 5215 7908 5908 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6914 7936 6920 7948
rect 6503 7908 6920 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 10318 7936 10324 7948
rect 9631 7908 10324 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13872 7908 14197 7936
rect 13872 7896 13878 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14458 7936 14464 7948
rect 14185 7899 14243 7905
rect 14292 7908 14464 7936
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 5261 7871 5319 7877
rect 2740 7840 3648 7868
rect 2740 7828 2746 7840
rect 3620 7809 3648 7840
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 6546 7868 6552 7880
rect 5307 7840 6552 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 14292 7868 14320 7908
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 12406 7840 14320 7868
rect 14369 7871 14427 7877
rect 2593 7803 2651 7809
rect 2593 7769 2605 7803
rect 2639 7800 2651 7803
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 2639 7772 3065 7800
rect 2639 7769 2651 7772
rect 2593 7763 2651 7769
rect 3053 7769 3065 7772
rect 3099 7769 3111 7803
rect 3053 7763 3111 7769
rect 3605 7803 3663 7809
rect 3605 7769 3617 7803
rect 3651 7800 3663 7803
rect 5353 7803 5411 7809
rect 3651 7772 4292 7800
rect 3651 7769 3663 7772
rect 3605 7763 3663 7769
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2038 7732 2044 7744
rect 1627 7704 2044 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2038 7692 2044 7704
rect 2096 7732 2102 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2096 7704 2697 7732
rect 2096 7692 2102 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 2685 7695 2743 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4264 7741 4292 7772
rect 5353 7769 5365 7803
rect 5399 7800 5411 7803
rect 5399 7772 5856 7800
rect 5399 7769 5411 7772
rect 5353 7763 5411 7769
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4430 7732 4436 7744
rect 4295 7704 4436 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7732 4951 7735
rect 5074 7732 5080 7744
rect 4939 7704 5080 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5828 7741 5856 7772
rect 5721 7735 5779 7741
rect 5721 7732 5733 7735
rect 5592 7704 5733 7732
rect 5592 7692 5598 7704
rect 5721 7701 5733 7704
rect 5767 7701 5779 7735
rect 5721 7695 5779 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 6052 7704 6193 7732
rect 6052 7692 6058 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6181 7695 6239 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6730 7732 6736 7744
rect 6319 7704 6736 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 9674 7732 9680 7744
rect 9635 7704 9680 7732
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10137 7735 10195 7741
rect 9824 7704 9869 7732
rect 9824 7692 9830 7704
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 12406 7732 12434 7840
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 15010 7868 15016 7880
rect 14415 7840 15016 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 12860 7772 14473 7800
rect 12860 7760 12866 7772
rect 14461 7769 14473 7772
rect 14507 7800 14519 7803
rect 15212 7800 15240 8035
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18598 8072 18604 8084
rect 18559 8044 18604 8072
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 19518 8072 19524 8084
rect 19479 8044 19524 8072
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21542 8072 21548 8084
rect 21407 8044 21548 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 17497 8007 17555 8013
rect 17497 7973 17509 8007
rect 17543 8004 17555 8007
rect 20346 8004 20352 8016
rect 17543 7976 20352 8004
rect 17543 7973 17555 7976
rect 17497 7967 17555 7973
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 20993 8007 21051 8013
rect 20993 7973 21005 8007
rect 21039 8004 21051 8007
rect 22094 8004 22100 8016
rect 21039 7976 22100 8004
rect 21039 7973 21051 7976
rect 20993 7967 21051 7973
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 16850 7936 16856 7948
rect 16811 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 18046 7936 18052 7948
rect 18007 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 19886 7936 19892 7948
rect 18196 7908 18241 7936
rect 18432 7908 19892 7936
rect 18196 7896 18202 7908
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16172 7840 17724 7868
rect 16172 7828 16178 7840
rect 14507 7772 15240 7800
rect 17037 7803 17095 7809
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 17037 7769 17049 7803
rect 17083 7800 17095 7803
rect 17696 7800 17724 7840
rect 18230 7800 18236 7812
rect 17083 7772 17632 7800
rect 17696 7772 18236 7800
rect 17083 7769 17095 7772
rect 17037 7763 17095 7769
rect 10183 7704 12434 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 15562 7732 15568 7744
rect 13596 7704 15568 7732
rect 13596 7692 13602 7704
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 17126 7732 17132 7744
rect 17087 7704 17132 7732
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17604 7741 17632 7772
rect 18230 7760 18236 7772
rect 18288 7800 18294 7812
rect 18432 7809 18460 7908
rect 19886 7896 19892 7908
rect 19944 7936 19950 7948
rect 19944 7908 20024 7936
rect 19944 7896 19950 7908
rect 18782 7868 18788 7880
rect 18743 7840 18788 7868
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 18984 7840 19349 7868
rect 18417 7803 18475 7809
rect 18417 7800 18429 7803
rect 18288 7772 18429 7800
rect 18288 7760 18294 7772
rect 18417 7769 18429 7772
rect 18463 7769 18475 7803
rect 18417 7763 18475 7769
rect 18984 7744 19012 7840
rect 19337 7837 19349 7840
rect 19383 7837 19395 7871
rect 19996 7868 20024 7908
rect 20070 7896 20076 7948
rect 20128 7936 20134 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 20128 7908 20177 7936
rect 20128 7896 20134 7908
rect 20165 7905 20177 7908
rect 20211 7905 20223 7939
rect 20165 7899 20223 7905
rect 20257 7939 20315 7945
rect 20257 7905 20269 7939
rect 20303 7905 20315 7939
rect 20257 7899 20315 7905
rect 20272 7868 20300 7899
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 19996 7840 20545 7868
rect 19337 7831 19395 7837
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20806 7868 20812 7880
rect 20767 7840 20812 7868
rect 20533 7831 20591 7837
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 21174 7868 21180 7880
rect 21135 7840 21180 7868
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 19978 7760 19984 7812
rect 20036 7800 20042 7812
rect 20073 7803 20131 7809
rect 20073 7800 20085 7803
rect 20036 7772 20085 7800
rect 20036 7760 20042 7772
rect 20073 7769 20085 7772
rect 20119 7769 20131 7803
rect 20073 7763 20131 7769
rect 17589 7735 17647 7741
rect 17589 7701 17601 7735
rect 17635 7701 17647 7735
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17589 7695 17647 7701
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18966 7732 18972 7744
rect 18927 7704 18972 7732
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 19668 7704 19717 7732
rect 19668 7692 19674 7704
rect 19705 7701 19717 7704
rect 19751 7701 19763 7735
rect 19705 7695 19763 7701
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2222 7528 2228 7540
rect 2087 7500 2228 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4304 7500 4353 7528
rect 4304 7488 4310 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 4341 7491 4399 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9824 7500 10333 7528
rect 9824 7488 9830 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10321 7491 10379 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15804 7500 15945 7528
rect 15804 7488 15810 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16439 7500 16957 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 16945 7491 17003 7497
rect 17037 7531 17095 7537
rect 17037 7497 17049 7531
rect 17083 7528 17095 7531
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 17083 7500 17509 7528
rect 17083 7497 17095 7500
rect 17037 7491 17095 7497
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 17957 7531 18015 7537
rect 17957 7497 17969 7531
rect 18003 7528 18015 7531
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 18003 7500 19165 7528
rect 18003 7497 18015 7500
rect 17957 7491 18015 7497
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 19153 7491 19211 7497
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 20346 7528 20352 7540
rect 19760 7500 20352 7528
rect 19760 7488 19766 7500
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20441 7531 20499 7537
rect 20441 7497 20453 7531
rect 20487 7528 20499 7531
rect 21082 7528 21088 7540
rect 20487 7500 21088 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 3326 7420 3332 7472
rect 3384 7460 3390 7472
rect 3973 7463 4031 7469
rect 3973 7460 3985 7463
rect 3384 7432 3985 7460
rect 3384 7420 3390 7432
rect 3973 7429 3985 7432
rect 4019 7429 4031 7463
rect 3973 7423 4031 7429
rect 7101 7463 7159 7469
rect 7101 7429 7113 7463
rect 7147 7460 7159 7463
rect 12066 7460 12072 7472
rect 7147 7432 12072 7460
rect 7147 7429 7159 7432
rect 7101 7423 7159 7429
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 18598 7460 18604 7472
rect 16071 7432 18604 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 18598 7420 18604 7432
rect 18656 7420 18662 7472
rect 18782 7460 18788 7472
rect 18743 7432 18788 7460
rect 18782 7420 18788 7432
rect 18840 7420 18846 7472
rect 20070 7420 20076 7472
rect 20128 7460 20134 7472
rect 20128 7432 20576 7460
rect 20128 7420 20134 7432
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 3418 7392 3424 7404
rect 2271 7364 3424 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 4246 7392 4252 7404
rect 4207 7364 4252 7392
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4706 7392 4712 7404
rect 4667 7364 4712 7392
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9398 7392 9404 7404
rect 8352 7364 9404 7392
rect 8352 7352 8358 7364
rect 9398 7352 9404 7364
rect 9456 7392 9462 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9456 7364 9965 7392
rect 9456 7352 9462 7364
rect 9953 7361 9965 7364
rect 9999 7392 10011 7395
rect 9999 7364 10916 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3384 7296 3709 7324
rect 3384 7284 3390 7296
rect 3697 7293 3709 7296
rect 3743 7324 3755 7327
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 3743 7296 4813 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7324 5043 7327
rect 5258 7324 5264 7336
rect 5031 7296 5264 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 8662 7324 8668 7336
rect 7423 7296 8668 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 5074 7216 5080 7268
rect 5132 7256 5138 7268
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 5132 7228 5641 7256
rect 5132 7216 5138 7228
rect 5629 7225 5641 7228
rect 5675 7256 5687 7259
rect 5994 7256 6000 7268
rect 5675 7228 6000 7256
rect 5675 7225 5687 7228
rect 5629 7219 5687 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 7208 7256 7236 7287
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 10778 7324 10784 7336
rect 10192 7296 10784 7324
rect 10192 7284 10198 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10888 7333 10916 7364
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 17862 7392 17868 7404
rect 11848 7364 15884 7392
rect 17823 7364 17868 7392
rect 11848 7352 11854 7364
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 15749 7327 15807 7333
rect 15749 7324 15761 7327
rect 14424 7296 15761 7324
rect 14424 7284 14430 7296
rect 15749 7293 15761 7296
rect 15795 7293 15807 7327
rect 15856 7324 15884 7364
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 20548 7392 20576 7432
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 21177 7463 21235 7469
rect 21177 7460 21189 7463
rect 20864 7432 21189 7460
rect 20864 7420 20870 7432
rect 21177 7429 21189 7432
rect 21223 7429 21235 7463
rect 21177 7423 21235 7429
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 19659 7364 20300 7392
rect 20548 7364 21005 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 15856 7296 16773 7324
rect 15749 7287 15807 7293
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 16761 7287 16819 7293
rect 16868 7296 18061 7324
rect 13170 7256 13176 7268
rect 7208 7228 13176 7256
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 15764 7256 15792 7287
rect 16868 7256 16896 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18288 7296 18889 7324
rect 18288 7284 18294 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 19300 7296 19717 7324
rect 19300 7284 19306 7296
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 20272 7324 20300 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 20533 7327 20591 7333
rect 20272 7296 20484 7324
rect 19705 7287 19763 7293
rect 15764 7228 16896 7256
rect 17405 7259 17463 7265
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 20254 7256 20260 7268
rect 17451 7228 20260 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 20254 7216 20260 7228
rect 20312 7216 20318 7268
rect 20456 7200 20484 7296
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20714 7324 20720 7336
rect 20579 7296 20720 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 20622 7216 20628 7268
rect 20680 7256 20686 7268
rect 21361 7259 21419 7265
rect 21361 7256 21373 7259
rect 20680 7228 21373 7256
rect 20680 7216 20686 7228
rect 21361 7225 21373 7228
rect 21407 7225 21419 7259
rect 21361 7219 21419 7225
rect 6730 7188 6736 7200
rect 6691 7160 6736 7188
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 10134 7188 10140 7200
rect 10095 7160 10140 7188
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 18138 7188 18144 7200
rect 15068 7160 18144 7188
rect 15068 7148 15074 7160
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 18322 7188 18328 7200
rect 18283 7160 18328 7188
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 19242 7188 19248 7200
rect 18472 7160 19248 7188
rect 18472 7148 18478 7160
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 19702 7148 19708 7200
rect 19760 7188 19766 7200
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19760 7160 19993 7188
rect 19760 7148 19766 7160
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20809 7191 20867 7197
rect 20809 7188 20821 7191
rect 20496 7160 20821 7188
rect 20496 7148 20502 7160
rect 20809 7157 20821 7160
rect 20855 7157 20867 7191
rect 20809 7151 20867 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 2593 6987 2651 6993
rect 2593 6984 2605 6987
rect 2188 6956 2605 6984
rect 2188 6944 2194 6956
rect 2593 6953 2605 6956
rect 2639 6953 2651 6987
rect 2593 6947 2651 6953
rect 17589 6987 17647 6993
rect 17589 6953 17601 6987
rect 17635 6984 17647 6987
rect 17862 6984 17868 6996
rect 17635 6956 17868 6984
rect 17635 6953 17647 6956
rect 17589 6947 17647 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 17954 6944 17960 6996
rect 18012 6984 18018 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18012 6956 19257 6984
rect 18012 6944 18018 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19886 6944 19892 6996
rect 19944 6984 19950 6996
rect 20073 6987 20131 6993
rect 20073 6984 20085 6987
rect 19944 6956 20085 6984
rect 19944 6944 19950 6956
rect 20073 6953 20085 6956
rect 20119 6984 20131 6987
rect 20714 6984 20720 6996
rect 20119 6956 20720 6984
rect 20119 6953 20131 6956
rect 20073 6947 20131 6953
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 20993 6919 21051 6925
rect 20993 6916 21005 6919
rect 4540 6888 4844 6916
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 3108 6820 3157 6848
rect 3108 6808 3114 6820
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3476 6820 4169 6848
rect 3476 6808 3482 6820
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 4540 6848 4568 6888
rect 4706 6848 4712 6860
rect 4157 6811 4215 6817
rect 4264 6820 4568 6848
rect 4667 6820 4712 6848
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4264 6780 4292 6820
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 4816 6848 4844 6888
rect 18156 6888 18552 6916
rect 5534 6848 5540 6860
rect 4816 6820 5212 6848
rect 5495 6820 5540 6848
rect 4120 6752 4292 6780
rect 4433 6783 4491 6789
rect 4120 6740 4126 6752
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 5184 6780 5212 6820
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 7190 6848 7196 6860
rect 5767 6820 7196 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 18156 6848 18184 6888
rect 10836 6820 18184 6848
rect 18233 6851 18291 6857
rect 10836 6808 10842 6820
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 18414 6848 18420 6860
rect 18279 6820 18420 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18524 6848 18552 6888
rect 19536 6888 21005 6916
rect 19536 6860 19564 6888
rect 20993 6885 21005 6888
rect 21039 6916 21051 6919
rect 21174 6916 21180 6928
rect 21039 6888 21180 6916
rect 21039 6885 21051 6888
rect 20993 6879 21051 6885
rect 21174 6876 21180 6888
rect 21232 6876 21238 6928
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 18524 6820 19073 6848
rect 19061 6817 19073 6820
rect 19107 6848 19119 6851
rect 19518 6848 19524 6860
rect 19107 6820 19524 6848
rect 19107 6817 19119 6820
rect 19061 6811 19119 6817
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 19886 6848 19892 6860
rect 19847 6820 19892 6848
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 20898 6848 20904 6860
rect 20811 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6848 20962 6860
rect 21082 6848 21088 6860
rect 20956 6820 21088 6848
rect 20956 6808 20962 6820
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 18966 6780 18972 6792
rect 4479 6752 5120 6780
rect 5184 6752 18972 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 2958 6644 2964 6656
rect 2919 6616 2964 6644
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3602 6644 3608 6656
rect 3099 6616 3608 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 5092 6653 5120 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19610 6780 19616 6792
rect 19571 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 17402 6712 17408 6724
rect 17363 6684 17408 6712
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 17957 6715 18015 6721
rect 17957 6681 17969 6715
rect 18003 6712 18015 6715
rect 18417 6715 18475 6721
rect 18417 6712 18429 6715
rect 18003 6684 18429 6712
rect 18003 6681 18015 6684
rect 17957 6675 18015 6681
rect 18417 6681 18429 6684
rect 18463 6681 18475 6715
rect 18417 6675 18475 6681
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6613 5135 6647
rect 5442 6644 5448 6656
rect 5403 6616 5448 6644
rect 5077 6607 5135 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 10502 6644 10508 6656
rect 7064 6616 10508 6644
rect 7064 6604 7070 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 14458 6644 14464 6656
rect 11756 6616 14464 6644
rect 11756 6604 11762 6616
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 17420 6644 17448 6672
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 17420 6616 18061 6644
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 18693 6647 18751 6653
rect 18693 6644 18705 6647
rect 18196 6616 18705 6644
rect 18196 6604 18202 6616
rect 18693 6613 18705 6616
rect 18739 6613 18751 6647
rect 18693 6607 18751 6613
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 20346 6644 20352 6656
rect 20220 6616 20352 6644
rect 20220 6604 20226 6616
rect 20346 6604 20352 6616
rect 20404 6644 20410 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 20404 6616 21189 6644
rect 20404 6604 20410 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3016 6412 3341 6440
rect 3016 6400 3022 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3602 6440 3608 6452
rect 3563 6412 3608 6440
rect 3329 6403 3387 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3936 6412 3985 6440
rect 3936 6400 3942 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 3973 6403 4031 6409
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4111 6412 4445 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4890 6440 4896 6452
rect 4851 6412 4896 6440
rect 4433 6403 4491 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5767 6412 6377 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6788 6412 6837 6440
rect 6788 6400 6794 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8294 6440 8300 6452
rect 8251 6412 8300 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 9674 6440 9680 6452
rect 9263 6412 9680 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6409 10011 6443
rect 12066 6440 12072 6452
rect 12027 6412 12072 6440
rect 9953 6403 10011 6409
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6372 4859 6375
rect 9968 6372 9996 6403
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12529 6443 12587 6449
rect 12529 6440 12541 6443
rect 12492 6412 12541 6440
rect 12492 6400 12498 6412
rect 12529 6409 12541 6412
rect 12575 6409 12587 6443
rect 12529 6403 12587 6409
rect 10778 6372 10784 6384
rect 4847 6344 9996 6372
rect 10336 6344 10784 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5224 6276 5641 6304
rect 5224 6264 5230 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 5629 6267 5687 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 10336 6313 10364 6344
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 11977 6375 12035 6381
rect 11977 6341 11989 6375
rect 12023 6372 12035 6375
rect 12158 6372 12164 6384
rect 12023 6344 12164 6372
rect 12023 6341 12035 6344
rect 11977 6335 12035 6341
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 12544 6372 12572 6403
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13044 6412 13921 6440
rect 13044 6400 13050 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 17126 6440 17132 6452
rect 16991 6412 17132 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17313 6443 17371 6449
rect 17313 6409 17325 6443
rect 17359 6440 17371 6443
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17359 6412 17785 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 18138 6440 18144 6452
rect 18099 6412 18144 6440
rect 17773 6403 17831 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 18322 6440 18328 6452
rect 18279 6412 18328 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 18598 6440 18604 6452
rect 18559 6412 18604 6440
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19061 6443 19119 6449
rect 19061 6409 19073 6443
rect 19107 6440 19119 6443
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19107 6412 19717 6440
rect 19107 6409 19119 6412
rect 19061 6403 19119 6409
rect 19705 6409 19717 6412
rect 19751 6440 19763 6443
rect 20622 6440 20628 6452
rect 19751 6412 20628 6440
rect 19751 6409 19763 6412
rect 19705 6403 19763 6409
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 13081 6375 13139 6381
rect 13081 6372 13093 6375
rect 12544 6344 13093 6372
rect 13081 6341 13093 6344
rect 13127 6341 13139 6375
rect 13081 6335 13139 6341
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 18046 6372 18052 6384
rect 13504 6344 18052 6372
rect 13504 6332 13510 6344
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8260 6276 8861 6304
rect 8260 6264 8266 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 8849 6267 8907 6273
rect 9324 6276 10333 6304
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 2866 6236 2872 6248
rect 2827 6208 2872 6236
rect 2685 6199 2743 6205
rect 2700 6168 2728 6199
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 4157 6239 4215 6245
rect 4157 6236 4169 6239
rect 3988 6208 4169 6236
rect 2774 6168 2780 6180
rect 2700 6140 2780 6168
rect 2774 6128 2780 6140
rect 2832 6168 2838 6180
rect 3988 6168 4016 6208
rect 4157 6205 4169 6208
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4580 6208 4997 6236
rect 4580 6196 4586 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 4985 6199 5043 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6638 6236 6644 6248
rect 6052 6208 6644 6236
rect 6052 6196 6058 6208
rect 6638 6196 6644 6208
rect 6696 6236 6702 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6696 6208 6929 6236
rect 6696 6196 6702 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8352 6208 8585 6236
rect 8352 6196 8358 6208
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 2832 6140 4016 6168
rect 2832 6128 2838 6140
rect 4246 6128 4252 6180
rect 4304 6168 4310 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 4304 6140 5273 6168
rect 4304 6128 4310 6140
rect 5261 6137 5273 6140
rect 5307 6137 5319 6171
rect 5261 6131 5319 6137
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 8772 6168 8800 6199
rect 9324 6177 9352 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 12437 6307 12495 6313
rect 10459 6276 11100 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10502 6236 10508 6248
rect 10463 6208 10508 6236
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 11072 6245 11100 6276
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12483 6276 13001 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12989 6273 13001 6276
rect 13035 6304 13047 6307
rect 13722 6304 13728 6316
rect 13035 6276 13728 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13832 6276 14289 6304
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 12526 6236 12532 6248
rect 11103 6208 12532 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 9309 6171 9367 6177
rect 9309 6168 9321 6171
rect 5592 6140 9321 6168
rect 5592 6128 5598 6140
rect 9309 6137 9321 6140
rect 9355 6137 9367 6171
rect 9309 6131 9367 6137
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8297 6103 8355 6109
rect 8297 6100 8309 6103
rect 8260 6072 8309 6100
rect 8260 6060 8266 6072
rect 8297 6069 8309 6072
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12636 6100 12664 6199
rect 13832 6112 13860 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 14384 6168 14412 6199
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 17402 6236 17408 6248
rect 14516 6208 14561 6236
rect 17363 6208 17408 6236
rect 14516 6196 14522 6208
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 17512 6245 17540 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 19978 6372 19984 6384
rect 19939 6344 19984 6372
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6304 19027 6307
rect 19518 6304 19524 6316
rect 19015 6276 19524 6304
rect 19015 6273 19027 6276
rect 18969 6267 19027 6273
rect 19518 6264 19524 6276
rect 19576 6304 19582 6316
rect 19794 6304 19800 6316
rect 19576 6276 19800 6304
rect 19576 6264 19582 6276
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 17828 6208 18337 6236
rect 17828 6196 17834 6208
rect 18325 6205 18337 6208
rect 18371 6205 18383 6239
rect 18325 6199 18383 6205
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 18472 6208 19165 6236
rect 18472 6196 18478 6208
rect 19153 6205 19165 6208
rect 19199 6205 19211 6239
rect 19153 6199 19211 6205
rect 14384 6140 14872 6168
rect 13814 6100 13820 6112
rect 12216 6072 12664 6100
rect 13775 6072 13820 6100
rect 12216 6060 12222 6072
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14844 6109 14872 6140
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15562 6100 15568 6112
rect 14875 6072 15568 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 19518 6100 19524 6112
rect 19479 6072 19524 6100
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 2958 5896 2964 5908
rect 2731 5868 2964 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 13814 5896 13820 5908
rect 4120 5868 13820 5896
rect 4120 5856 4126 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 17460 5868 19257 5896
rect 17460 5856 17466 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 5534 5828 5540 5840
rect 2556 5800 5540 5828
rect 2556 5788 2562 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6365 5831 6423 5837
rect 6365 5828 6377 5831
rect 5684 5800 6377 5828
rect 5684 5788 5690 5800
rect 6365 5797 6377 5800
rect 6411 5797 6423 5831
rect 6365 5791 6423 5797
rect 10778 5788 10784 5840
rect 10836 5828 10842 5840
rect 17954 5828 17960 5840
rect 10836 5800 17960 5828
rect 10836 5788 10842 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2832 5732 3341 5760
rect 2832 5720 2838 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 4522 5760 4528 5772
rect 3375 5732 4528 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5776 5732 6193 5760
rect 5776 5720 5782 5732
rect 6181 5729 6193 5732
rect 6227 5760 6239 5763
rect 6638 5760 6644 5772
rect 6227 5732 6644 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6880 5732 6929 5760
rect 6880 5720 6886 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 17770 5720 17776 5772
rect 17828 5760 17834 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 17828 5732 19809 5760
rect 17828 5720 17834 5732
rect 19797 5729 19809 5732
rect 19843 5760 19855 5763
rect 19886 5760 19892 5772
rect 19843 5732 19892 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 20625 5763 20683 5769
rect 20625 5760 20637 5763
rect 20036 5732 20637 5760
rect 20036 5720 20042 5732
rect 20625 5729 20637 5732
rect 20671 5729 20683 5763
rect 20625 5723 20683 5729
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5810 5692 5816 5704
rect 5408 5664 5816 5692
rect 5408 5652 5414 5664
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7190 5692 7196 5704
rect 6779 5664 7196 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 2593 5627 2651 5633
rect 2593 5593 2605 5627
rect 2639 5624 2651 5627
rect 3053 5627 3111 5633
rect 3053 5624 3065 5627
rect 2639 5596 3065 5624
rect 2639 5593 2651 5596
rect 2593 5587 2651 5593
rect 3053 5593 3065 5596
rect 3099 5593 3111 5627
rect 3053 5587 3111 5593
rect 6089 5627 6147 5633
rect 6089 5593 6101 5627
rect 6135 5624 6147 5627
rect 6546 5624 6552 5636
rect 6135 5596 6552 5624
rect 6135 5593 6147 5596
rect 6089 5587 6147 5593
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 10134 5624 10140 5636
rect 6748 5596 10140 5624
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5556 2286 5568
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 2280 5528 3157 5556
rect 2280 5516 2286 5528
rect 3145 5525 3157 5528
rect 3191 5556 3203 5559
rect 3786 5556 3792 5568
rect 3191 5528 3792 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 6748 5556 6776 5596
rect 10134 5584 10140 5596
rect 10192 5584 10198 5636
rect 19613 5627 19671 5633
rect 19613 5593 19625 5627
rect 19659 5624 19671 5627
rect 20438 5624 20444 5636
rect 19659 5596 20116 5624
rect 20351 5596 20444 5624
rect 19659 5593 19671 5596
rect 19613 5587 19671 5593
rect 4028 5528 6776 5556
rect 6825 5559 6883 5565
rect 4028 5516 4034 5528
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 7098 5556 7104 5568
rect 6871 5528 7104 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 20088 5565 20116 5596
rect 20438 5584 20444 5596
rect 20496 5624 20502 5636
rect 20496 5596 21220 5624
rect 20496 5584 20502 5596
rect 21192 5568 21220 5596
rect 20073 5559 20131 5565
rect 20073 5525 20085 5559
rect 20119 5525 20131 5559
rect 20073 5519 20131 5525
rect 20254 5516 20260 5568
rect 20312 5556 20318 5568
rect 20533 5559 20591 5565
rect 20533 5556 20545 5559
rect 20312 5528 20545 5556
rect 20312 5516 20318 5528
rect 20533 5525 20545 5528
rect 20579 5556 20591 5559
rect 20901 5559 20959 5565
rect 20901 5556 20913 5559
rect 20579 5528 20913 5556
rect 20579 5525 20591 5528
rect 20533 5519 20591 5525
rect 20901 5525 20913 5528
rect 20947 5525 20959 5559
rect 21174 5556 21180 5568
rect 21135 5528 21180 5556
rect 20901 5519 20959 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 2924 5324 3249 5352
rect 2924 5312 2930 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 6181 5355 6239 5361
rect 4120 5324 6132 5352
rect 4120 5312 4126 5324
rect 2777 5287 2835 5293
rect 2777 5253 2789 5287
rect 2823 5284 2835 5287
rect 2823 5256 4936 5284
rect 2823 5253 2835 5256
rect 2777 5247 2835 5253
rect 2130 5176 2136 5228
rect 2188 5216 2194 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2188 5188 2881 5216
rect 2188 5176 2194 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 2225 5083 2283 5089
rect 2225 5049 2237 5083
rect 2271 5080 2283 5083
rect 2700 5080 2728 5111
rect 2774 5080 2780 5092
rect 2271 5052 2452 5080
rect 2700 5052 2780 5080
rect 2271 5049 2283 5052
rect 2225 5043 2283 5049
rect 2130 4972 2136 5024
rect 2188 5012 2194 5024
rect 2317 5015 2375 5021
rect 2317 5012 2329 5015
rect 2188 4984 2329 5012
rect 2188 4972 2194 4984
rect 2317 4981 2329 4984
rect 2363 4981 2375 5015
rect 2424 5012 2452 5052
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 2976 5012 3004 5256
rect 3786 5216 3792 5228
rect 3699 5188 3792 5216
rect 3786 5176 3792 5188
rect 3844 5216 3850 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 3844 5188 4445 5216
rect 3844 5176 3850 5188
rect 4433 5185 4445 5188
rect 4479 5216 4491 5219
rect 4908 5216 4936 5256
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 5813 5287 5871 5293
rect 5813 5284 5825 5287
rect 5776 5256 5825 5284
rect 5776 5244 5782 5256
rect 5813 5253 5825 5256
rect 5859 5253 5871 5287
rect 6104 5284 6132 5324
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6730 5352 6736 5364
rect 6227 5324 6736 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 7098 5352 7104 5364
rect 7059 5324 7104 5352
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7248 5324 7293 5352
rect 7248 5312 7254 5324
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 17954 5352 17960 5364
rect 15620 5324 17960 5352
rect 15620 5312 15626 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 19429 5355 19487 5361
rect 19429 5321 19441 5355
rect 19475 5352 19487 5355
rect 19702 5352 19708 5364
rect 19475 5324 19708 5352
rect 19475 5321 19487 5324
rect 19429 5315 19487 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 8202 5284 8208 5296
rect 6104 5256 8208 5284
rect 5813 5247 5871 5253
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 19337 5287 19395 5293
rect 19337 5253 19349 5287
rect 19383 5284 19395 5287
rect 19978 5284 19984 5296
rect 19383 5256 19984 5284
rect 19383 5253 19395 5256
rect 19337 5247 19395 5253
rect 19978 5244 19984 5256
rect 20036 5244 20042 5296
rect 6546 5216 6552 5228
rect 4479 5188 4844 5216
rect 4908 5188 6552 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4525 5151 4583 5157
rect 4525 5148 4537 5151
rect 3896 5120 4537 5148
rect 3234 5040 3240 5092
rect 3292 5080 3298 5092
rect 3896 5089 3924 5120
rect 4525 5117 4537 5120
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 3881 5083 3939 5089
rect 3881 5080 3893 5083
rect 3292 5052 3893 5080
rect 3292 5040 3298 5052
rect 3881 5049 3893 5052
rect 3927 5049 3939 5083
rect 3881 5043 3939 5049
rect 3050 5012 3056 5024
rect 2424 4984 3056 5012
rect 2317 4975 2375 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4246 5012 4252 5024
rect 4111 4984 4252 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4724 5012 4752 5111
rect 4816 5080 4844 5188
rect 6546 5176 6552 5188
rect 6604 5216 6610 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6604 5188 6745 5216
rect 6604 5176 6610 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7607 5188 8033 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19576 5188 19809 5216
rect 19576 5176 19582 5188
rect 19797 5185 19809 5188
rect 19843 5216 19855 5219
rect 20530 5216 20536 5228
rect 19843 5188 20536 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5408 5120 5549 5148
rect 5408 5108 5414 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6362 5148 6368 5160
rect 5767 5120 6368 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6638 5148 6644 5160
rect 6512 5120 6557 5148
rect 6599 5120 6644 5148
rect 6512 5108 6518 5120
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 7650 5148 7656 5160
rect 7611 5120 7656 5148
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 19889 5151 19947 5157
rect 7800 5120 7845 5148
rect 7800 5108 7806 5120
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 7668 5080 7696 5108
rect 4816 5052 7696 5080
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4724 4984 4997 5012
rect 4985 4981 4997 4984
rect 5031 5012 5043 5015
rect 6086 5012 6092 5024
rect 5031 4984 6092 5012
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 19904 5012 19932 5111
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20036 5120 20081 5148
rect 20036 5108 20042 5120
rect 20346 5012 20352 5024
rect 19904 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20530 5012 20536 5024
rect 20491 4984 20536 5012
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3384 4780 3985 4808
rect 3384 4768 3390 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 3973 4771 4031 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3988 4604 4016 4771
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 7650 4808 7656 4820
rect 7331 4780 7656 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 5350 4700 5356 4752
rect 5408 4740 5414 4752
rect 8662 4740 8668 4752
rect 5408 4712 8668 4740
rect 5408 4700 5414 4712
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 5534 4672 5540 4684
rect 4663 4644 5540 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5902 4672 5908 4684
rect 5863 4644 5908 4672
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6546 4672 6552 4684
rect 6144 4644 6552 4672
rect 6144 4632 6150 4644
rect 6546 4632 6552 4644
rect 6604 4672 6610 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6604 4644 7021 4672
rect 6604 4632 6610 4644
rect 7009 4641 7021 4644
rect 7055 4672 7067 4675
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 7055 4644 7481 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7469 4641 7481 4644
rect 7515 4672 7527 4675
rect 12158 4672 12164 4684
rect 7515 4644 12164 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 3988 4576 4813 4604
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6696 4576 6745 4604
rect 6696 4564 6702 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 4709 4539 4767 4545
rect 4709 4536 4721 4539
rect 3191 4508 4721 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 3896 4480 3924 4508
rect 4709 4505 4721 4508
rect 4755 4505 4767 4539
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 4709 4499 4767 4505
rect 5184 4508 5733 4536
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4338 4468 4344 4480
rect 4299 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 5184 4477 5212 4508
rect 5721 4505 5733 4508
rect 5767 4505 5779 4539
rect 5721 4499 5779 4505
rect 6825 4539 6883 4545
rect 6825 4505 6837 4539
rect 6871 4536 6883 4539
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 6871 4508 7665 4536
rect 6871 4505 6883 4508
rect 6825 4499 6883 4505
rect 7653 4505 7665 4508
rect 7699 4536 7711 4539
rect 18690 4536 18696 4548
rect 7699 4508 18696 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 18690 4496 18696 4508
rect 18748 4496 18754 4548
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4437 5227 4471
rect 5626 4468 5632 4480
rect 5587 4440 5632 4468
rect 5169 4431 5227 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 5868 4440 6101 4468
rect 5868 4428 5874 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3292 4236 3801 4264
rect 3292 4224 3298 4236
rect 3789 4233 3801 4236
rect 3835 4264 3847 4267
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 3835 4236 5273 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5810 4264 5816 4276
rect 5771 4236 5816 4264
rect 5261 4227 5319 4233
rect 4709 4199 4767 4205
rect 4709 4196 4721 4199
rect 3988 4168 4721 4196
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4029 2743 4063
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2685 4023 2743 4029
rect 2700 3992 2728 4023
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3878 4060 3884 4072
rect 3839 4032 3884 4060
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 2774 3992 2780 4004
rect 2700 3964 2780 3992
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 3329 3995 3387 4001
rect 3329 3961 3341 3995
rect 3375 3992 3387 3995
rect 3988 3992 4016 4168
rect 4709 4165 4721 4168
rect 4755 4165 4767 4199
rect 4709 4159 4767 4165
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4080 4100 4353 4128
rect 4080 4069 4108 4100
rect 4341 4097 4353 4100
rect 4387 4128 4399 4131
rect 4614 4128 4620 4140
rect 4387 4100 4620 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4798 4128 4804 4140
rect 4759 4100 4804 4128
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5276 4128 5304 4227
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6052 4236 6469 4264
rect 6052 4224 6058 4236
rect 6457 4233 6469 4236
rect 6503 4264 6515 4267
rect 6638 4264 6644 4276
rect 6503 4236 6644 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 6822 4196 6828 4208
rect 5592 4168 6828 4196
rect 5592 4156 5598 4168
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5276 4100 5917 4128
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4060 4583 4063
rect 5810 4060 5816 4072
rect 4571 4032 5816 4060
rect 4571 4029 4583 4032
rect 4525 4023 4583 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6012 4069 6040 4168
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 5166 3992 5172 4004
rect 3375 3964 4016 3992
rect 5127 3964 5172 3992
rect 3375 3961 3387 3964
rect 3329 3955 3387 3961
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 5445 3995 5503 4001
rect 5445 3961 5457 3995
rect 5491 3992 5503 3995
rect 5626 3992 5632 4004
rect 5491 3964 5632 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 3200 3896 3433 3924
rect 3200 3884 3206 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2130 3720 2136 3732
rect 2091 3692 2136 3720
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3237 3723 3295 3729
rect 3237 3720 3249 3723
rect 3016 3692 3249 3720
rect 3016 3680 3022 3692
rect 3237 3689 3249 3692
rect 3283 3689 3295 3723
rect 3237 3683 3295 3689
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3720 4767 3723
rect 4798 3720 4804 3732
rect 4755 3692 4804 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3720 5963 3723
rect 6546 3720 6552 3732
rect 5951 3692 6552 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 2332 3448 2360 3680
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 5350 3652 5356 3664
rect 2832 3624 5356 3652
rect 2832 3612 2838 3624
rect 4080 3593 4108 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 4065 3587 4123 3593
rect 2731 3556 3464 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 2464 3488 2881 3516
rect 2464 3476 2470 3488
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 2777 3451 2835 3457
rect 2777 3448 2789 3451
rect 2332 3420 2789 3448
rect 2777 3417 2789 3420
rect 2823 3448 2835 3451
rect 3326 3448 3332 3460
rect 2823 3420 3332 3448
rect 2823 3417 2835 3420
rect 2777 3411 2835 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 3436 3457 3464 3556
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4246 3584 4252 3596
rect 4207 3556 4252 3584
rect 4065 3547 4123 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5534 3584 5540 3596
rect 5215 3556 5540 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 4338 3516 4344 3528
rect 4299 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4672 3488 5365 3516
rect 4672 3476 4678 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 3421 3451 3479 3457
rect 3421 3417 3433 3451
rect 3467 3448 3479 3451
rect 5460 3448 5488 3556
rect 5534 3544 5540 3556
rect 5592 3584 5598 3596
rect 5920 3584 5948 3683
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 5592 3556 5948 3584
rect 5592 3544 5598 3556
rect 3467 3420 5488 3448
rect 3467 3417 3479 3420
rect 3421 3411 3479 3417
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 4212 3352 4813 3380
rect 4212 3340 4218 3352
rect 4801 3349 4813 3352
rect 4847 3380 4859 3383
rect 5074 3380 5080 3392
rect 4847 3352 5080 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 5074 3340 5080 3352
rect 5132 3380 5138 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 5132 3352 5273 3380
rect 5132 3340 5138 3352
rect 5261 3349 5273 3352
rect 5307 3349 5319 3383
rect 5261 3343 5319 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 3605 3179 3663 3185
rect 3605 3176 3617 3179
rect 2924 3148 3617 3176
rect 2924 3136 2930 3148
rect 3605 3145 3617 3148
rect 3651 3145 3663 3179
rect 5534 3176 5540 3188
rect 3605 3139 3663 3145
rect 5092 3148 5540 3176
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3237 3111 3295 3117
rect 3237 3108 3249 3111
rect 3108 3080 3249 3108
rect 3108 3068 3114 3080
rect 3237 3077 3249 3080
rect 3283 3108 3295 3111
rect 3973 3111 4031 3117
rect 3973 3108 3985 3111
rect 3283 3080 3985 3108
rect 3283 3077 3295 3080
rect 3237 3071 3295 3077
rect 3973 3077 3985 3080
rect 4019 3077 4031 3111
rect 3973 3071 4031 3077
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 5092 3108 5120 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5258 3108 5264 3120
rect 4571 3080 5120 3108
rect 5219 3080 5264 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2972 3482 2984
rect 3878 2972 3884 2984
rect 3476 2944 3884 2972
rect 3476 2932 3482 2944
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3936 2944 4077 2972
rect 3936 2932 3942 2944
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2972 4307 2975
rect 4540 2972 4568 3071
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 18877 3111 18935 3117
rect 18877 3108 18889 3111
rect 7616 3080 18889 3108
rect 7616 3068 7622 3080
rect 18877 3077 18889 3080
rect 18923 3077 18935 3111
rect 18877 3071 18935 3077
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 12250 3040 12256 3052
rect 5583 3012 5764 3040
rect 12211 3012 12256 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 4295 2944 4568 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 2222 2864 2228 2916
rect 2280 2904 2286 2916
rect 4982 2904 4988 2916
rect 2280 2876 4988 2904
rect 2280 2864 2286 2876
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5736 2845 5764 3012
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 19153 3043 19211 3049
rect 12575 3012 12756 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 5721 2839 5779 2845
rect 5721 2805 5733 2839
rect 5767 2836 5779 2839
rect 11238 2836 11244 2848
rect 5767 2808 11244 2836
rect 5767 2805 5779 2808
rect 5721 2799 5779 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 12728 2845 12756 3012
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19199 3012 19380 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 12713 2839 12771 2845
rect 12713 2805 12725 2839
rect 12759 2836 12771 2839
rect 16022 2836 16028 2848
rect 12759 2808 16028 2836
rect 12759 2805 12771 2808
rect 12713 2799 12771 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 19352 2845 19380 3012
rect 19337 2839 19395 2845
rect 19337 2805 19349 2839
rect 19383 2836 19395 2839
rect 20622 2836 20628 2848
rect 19383 2808 20628 2836
rect 19383 2805 19395 2808
rect 19337 2799 19395 2805
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 5994 2632 6000 2644
rect 4120 2604 6000 2632
rect 4120 2592 4126 2604
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
<< via1 >>
rect 5172 21020 5224 21072
rect 7380 21020 7432 21072
rect 3884 20952 3936 21004
rect 11060 20952 11112 21004
rect 2964 20884 3016 20936
rect 16212 20884 16264 20936
rect 1676 20816 1728 20868
rect 5816 20816 5868 20868
rect 6828 20816 6880 20868
rect 13820 20816 13872 20868
rect 15108 20816 15160 20868
rect 20168 20748 20220 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 2872 20587 2924 20596
rect 2872 20553 2881 20587
rect 2881 20553 2915 20587
rect 2915 20553 2924 20587
rect 2872 20544 2924 20553
rect 4436 20587 4488 20596
rect 4436 20553 4445 20587
rect 4445 20553 4479 20587
rect 4479 20553 4488 20587
rect 4436 20544 4488 20553
rect 2044 20476 2096 20528
rect 6184 20544 6236 20596
rect 7196 20544 7248 20596
rect 7380 20587 7432 20596
rect 7380 20553 7389 20587
rect 7389 20553 7423 20587
rect 7423 20553 7432 20587
rect 7380 20544 7432 20553
rect 9312 20544 9364 20596
rect 9588 20544 9640 20596
rect 10048 20544 10100 20596
rect 6736 20476 6788 20528
rect 4252 20408 4304 20460
rect 4988 20451 5040 20460
rect 4988 20417 4997 20451
rect 4997 20417 5031 20451
rect 5031 20417 5040 20451
rect 4988 20408 5040 20417
rect 7012 20476 7064 20528
rect 7472 20519 7524 20528
rect 7472 20485 7481 20519
rect 7481 20485 7515 20519
rect 7515 20485 7524 20519
rect 7472 20476 7524 20485
rect 7748 20476 7800 20528
rect 8208 20519 8260 20528
rect 8208 20485 8217 20519
rect 8217 20485 8251 20519
rect 8251 20485 8260 20519
rect 8208 20476 8260 20485
rect 15568 20544 15620 20596
rect 16028 20544 16080 20596
rect 16396 20544 16448 20596
rect 19340 20544 19392 20596
rect 11060 20519 11112 20528
rect 4160 20383 4212 20392
rect 4160 20349 4169 20383
rect 4169 20349 4203 20383
rect 4203 20349 4212 20383
rect 4160 20340 4212 20349
rect 5172 20340 5224 20392
rect 7656 20408 7708 20460
rect 8024 20383 8076 20392
rect 4436 20272 4488 20324
rect 8024 20349 8033 20383
rect 8033 20349 8067 20383
rect 8067 20349 8076 20383
rect 8024 20340 8076 20349
rect 8116 20340 8168 20392
rect 11060 20485 11069 20519
rect 11069 20485 11103 20519
rect 11103 20485 11112 20519
rect 11060 20476 11112 20485
rect 12900 20476 12952 20528
rect 12992 20476 13044 20528
rect 13452 20476 13504 20528
rect 13544 20476 13596 20528
rect 14740 20476 14792 20528
rect 8668 20408 8720 20460
rect 9128 20408 9180 20460
rect 9312 20451 9364 20460
rect 9312 20417 9321 20451
rect 9321 20417 9355 20451
rect 9355 20417 9364 20451
rect 9312 20408 9364 20417
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 7472 20272 7524 20324
rect 8208 20272 8260 20324
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 10876 20340 10928 20392
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 12440 20408 12492 20460
rect 15016 20408 15068 20460
rect 15844 20408 15896 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 14372 20340 14424 20392
rect 14648 20340 14700 20392
rect 6552 20204 6604 20256
rect 6920 20247 6972 20256
rect 6920 20213 6929 20247
rect 6929 20213 6963 20247
rect 6963 20213 6972 20247
rect 6920 20204 6972 20213
rect 7380 20204 7432 20256
rect 7840 20204 7892 20256
rect 9496 20272 9548 20324
rect 13084 20272 13136 20324
rect 13452 20315 13504 20324
rect 13452 20281 13461 20315
rect 13461 20281 13495 20315
rect 13495 20281 13504 20315
rect 13452 20272 13504 20281
rect 14832 20272 14884 20324
rect 16396 20272 16448 20324
rect 9404 20204 9456 20256
rect 11520 20204 11572 20256
rect 11980 20204 12032 20256
rect 12440 20204 12492 20256
rect 13176 20204 13228 20256
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13268 20204 13320 20213
rect 13544 20204 13596 20256
rect 13820 20204 13872 20256
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 16580 20204 16632 20256
rect 17960 20247 18012 20256
rect 17960 20213 17969 20247
rect 17969 20213 18003 20247
rect 18003 20213 18012 20247
rect 17960 20204 18012 20213
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 21272 20204 21324 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2780 20000 2832 20052
rect 2964 20000 3016 20052
rect 4252 20000 4304 20052
rect 5540 20000 5592 20052
rect 5632 20000 5684 20052
rect 7472 20000 7524 20052
rect 10232 20000 10284 20052
rect 10876 20000 10928 20052
rect 11520 20000 11572 20052
rect 6828 19932 6880 19984
rect 11060 19975 11112 19984
rect 4436 19796 4488 19848
rect 7380 19864 7432 19916
rect 9496 19864 9548 19916
rect 11060 19941 11069 19975
rect 11069 19941 11103 19975
rect 11103 19941 11112 19975
rect 11060 19932 11112 19941
rect 11152 19932 11204 19984
rect 4252 19728 4304 19780
rect 2688 19703 2740 19712
rect 2688 19669 2697 19703
rect 2697 19669 2731 19703
rect 2731 19669 2740 19703
rect 2688 19660 2740 19669
rect 3976 19660 4028 19712
rect 6920 19796 6972 19848
rect 7196 19796 7248 19848
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9220 19796 9272 19848
rect 14096 20043 14148 20052
rect 12164 19932 12216 19984
rect 12348 19932 12400 19984
rect 5540 19660 5592 19712
rect 6644 19660 6696 19712
rect 6736 19660 6788 19712
rect 8208 19728 8260 19780
rect 7380 19660 7432 19712
rect 7472 19660 7524 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 8760 19703 8812 19712
rect 7656 19660 7708 19669
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 8944 19660 8996 19712
rect 9496 19660 9548 19712
rect 12348 19796 12400 19848
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 13452 19932 13504 19984
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 14556 20000 14608 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 15108 19975 15160 19984
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 13820 19864 13872 19916
rect 14556 19864 14608 19916
rect 14832 19864 14884 19916
rect 15108 19941 15117 19975
rect 15117 19941 15151 19975
rect 15151 19941 15160 19975
rect 15108 19932 15160 19941
rect 15200 19932 15252 19984
rect 17408 19932 17460 19984
rect 17868 20000 17920 20052
rect 18604 20000 18656 20052
rect 19708 20000 19760 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 21180 20000 21232 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 18144 19932 18196 19984
rect 20996 19975 21048 19984
rect 15476 19864 15528 19916
rect 15568 19864 15620 19916
rect 13636 19796 13688 19848
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16764 19839 16816 19848
rect 16212 19796 16264 19805
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 16948 19796 17000 19848
rect 12900 19728 12952 19780
rect 10876 19660 10928 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 12440 19660 12492 19669
rect 13176 19660 13228 19712
rect 14096 19728 14148 19780
rect 14372 19728 14424 19780
rect 16028 19728 16080 19780
rect 17684 19728 17736 19780
rect 18236 19864 18288 19916
rect 20996 19941 21005 19975
rect 21005 19941 21039 19975
rect 21039 19941 21048 19975
rect 20996 19932 21048 19941
rect 17960 19796 18012 19848
rect 18420 19839 18472 19848
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 18236 19728 18288 19780
rect 20168 19796 20220 19848
rect 20720 19796 20772 19848
rect 20996 19796 21048 19848
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 15752 19660 15804 19712
rect 17224 19660 17276 19712
rect 17500 19660 17552 19712
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 3056 19456 3108 19508
rect 3976 19456 4028 19508
rect 4436 19499 4488 19508
rect 4436 19465 4445 19499
rect 4445 19465 4479 19499
rect 4479 19465 4488 19499
rect 4436 19456 4488 19465
rect 6184 19499 6236 19508
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 6736 19499 6788 19508
rect 6736 19465 6745 19499
rect 6745 19465 6779 19499
rect 6779 19465 6788 19499
rect 6736 19456 6788 19465
rect 7012 19456 7064 19508
rect 7196 19456 7248 19508
rect 8944 19456 8996 19508
rect 9404 19456 9456 19508
rect 6920 19388 6972 19440
rect 10232 19456 10284 19508
rect 12624 19456 12676 19508
rect 12900 19456 12952 19508
rect 13268 19456 13320 19508
rect 13728 19456 13780 19508
rect 14924 19499 14976 19508
rect 9956 19431 10008 19440
rect 5540 19320 5592 19372
rect 7380 19320 7432 19372
rect 8024 19320 8076 19372
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 9588 19320 9640 19372
rect 9956 19397 9990 19431
rect 9990 19397 10008 19431
rect 9956 19388 10008 19397
rect 12348 19388 12400 19440
rect 14924 19465 14933 19499
rect 14933 19465 14967 19499
rect 14967 19465 14976 19499
rect 14924 19456 14976 19465
rect 15200 19456 15252 19508
rect 15384 19456 15436 19508
rect 16396 19499 16448 19508
rect 16396 19465 16405 19499
rect 16405 19465 16439 19499
rect 16439 19465 16448 19499
rect 16396 19456 16448 19465
rect 16948 19456 17000 19508
rect 11244 19320 11296 19372
rect 12072 19320 12124 19372
rect 12808 19320 12860 19372
rect 4068 19252 4120 19304
rect 15660 19388 15712 19440
rect 13360 19320 13412 19372
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 15108 19363 15160 19372
rect 14372 19320 14424 19329
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 15568 19363 15620 19372
rect 15568 19329 15577 19363
rect 15577 19329 15611 19363
rect 15611 19329 15620 19363
rect 15568 19320 15620 19329
rect 4620 19116 4672 19168
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 6920 19116 6972 19168
rect 10968 19116 11020 19168
rect 11152 19116 11204 19168
rect 11704 19116 11756 19168
rect 12532 19116 12584 19168
rect 13820 19252 13872 19304
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 16948 19320 17000 19372
rect 17224 19388 17276 19440
rect 21088 19456 21140 19508
rect 17960 19388 18012 19440
rect 15752 19252 15804 19261
rect 16396 19252 16448 19304
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 17684 19252 17736 19304
rect 18236 19388 18288 19440
rect 18328 19363 18380 19372
rect 18328 19329 18337 19363
rect 18337 19329 18371 19363
rect 18371 19329 18380 19363
rect 18328 19320 18380 19329
rect 18604 19320 18656 19372
rect 13176 19184 13228 19236
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 15476 19116 15528 19168
rect 17316 19184 17368 19236
rect 18972 19116 19024 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 22376 19116 22428 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 4436 18955 4488 18964
rect 4436 18921 4445 18955
rect 4445 18921 4479 18955
rect 4479 18921 4488 18955
rect 4436 18912 4488 18921
rect 4988 18912 5040 18964
rect 6552 18912 6604 18964
rect 7012 18912 7064 18964
rect 9312 18912 9364 18964
rect 9588 18912 9640 18964
rect 7380 18887 7432 18896
rect 7380 18853 7389 18887
rect 7389 18853 7423 18887
rect 7423 18853 7432 18887
rect 7380 18844 7432 18853
rect 9220 18844 9272 18896
rect 12440 18912 12492 18964
rect 12624 18912 12676 18964
rect 14372 18912 14424 18964
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 20628 18912 20680 18964
rect 11060 18887 11112 18896
rect 11060 18853 11069 18887
rect 11069 18853 11103 18887
rect 11103 18853 11112 18887
rect 11060 18844 11112 18853
rect 12808 18844 12860 18896
rect 7196 18776 7248 18828
rect 7564 18776 7616 18828
rect 8944 18776 8996 18828
rect 6000 18708 6052 18760
rect 6368 18751 6420 18760
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 7104 18708 7156 18760
rect 8208 18708 8260 18760
rect 12532 18776 12584 18828
rect 13176 18819 13228 18828
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 15752 18776 15804 18828
rect 3976 18640 4028 18692
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 4988 18683 5040 18692
rect 4988 18649 5022 18683
rect 5022 18649 5040 18683
rect 4988 18640 5040 18649
rect 8392 18640 8444 18692
rect 5540 18572 5592 18624
rect 6552 18572 6604 18624
rect 7380 18572 7432 18624
rect 7932 18572 7984 18624
rect 8944 18572 8996 18624
rect 9036 18572 9088 18624
rect 9312 18572 9364 18624
rect 9680 18572 9732 18624
rect 9864 18683 9916 18692
rect 9864 18649 9898 18683
rect 9898 18649 9916 18683
rect 9864 18640 9916 18649
rect 9956 18572 10008 18624
rect 10876 18708 10928 18760
rect 10508 18640 10560 18692
rect 11152 18640 11204 18692
rect 11704 18708 11756 18760
rect 12164 18751 12216 18760
rect 12164 18717 12182 18751
rect 12182 18717 12216 18751
rect 12164 18708 12216 18717
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 16212 18708 16264 18760
rect 17684 18844 17736 18896
rect 20720 18844 20772 18896
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 13728 18640 13780 18692
rect 15200 18640 15252 18692
rect 16396 18683 16448 18692
rect 11888 18572 11940 18624
rect 12716 18572 12768 18624
rect 12808 18572 12860 18624
rect 15660 18572 15712 18624
rect 16396 18649 16405 18683
rect 16405 18649 16439 18683
rect 16439 18649 16448 18683
rect 16396 18640 16448 18649
rect 18788 18640 18840 18692
rect 16304 18572 16356 18624
rect 21088 18572 21140 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 2780 18368 2832 18420
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 6184 18411 6236 18420
rect 6184 18377 6193 18411
rect 6193 18377 6227 18411
rect 6227 18377 6236 18411
rect 6184 18368 6236 18377
rect 6828 18368 6880 18420
rect 7656 18368 7708 18420
rect 12348 18368 12400 18420
rect 12624 18368 12676 18420
rect 13176 18368 13228 18420
rect 14004 18368 14056 18420
rect 15568 18411 15620 18420
rect 5540 18343 5592 18352
rect 5540 18309 5558 18343
rect 5558 18309 5592 18343
rect 5540 18300 5592 18309
rect 2412 18232 2464 18284
rect 4252 18232 4304 18284
rect 7288 18300 7340 18352
rect 6644 18275 6696 18284
rect 6644 18241 6678 18275
rect 6678 18241 6696 18275
rect 6644 18232 6696 18241
rect 8024 18232 8076 18284
rect 11244 18232 11296 18284
rect 12164 18300 12216 18352
rect 12532 18232 12584 18284
rect 12808 18300 12860 18352
rect 13360 18300 13412 18352
rect 13636 18343 13688 18352
rect 13636 18309 13645 18343
rect 13645 18309 13679 18343
rect 13679 18309 13688 18343
rect 13636 18300 13688 18309
rect 15108 18343 15160 18352
rect 14188 18232 14240 18284
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 2504 18096 2556 18148
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 4712 18028 4764 18080
rect 6184 18028 6236 18080
rect 7380 18028 7432 18080
rect 7656 18028 7708 18080
rect 7840 18028 7892 18080
rect 10232 18164 10284 18216
rect 9864 18096 9916 18148
rect 10324 18096 10376 18148
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10048 18028 10100 18080
rect 13728 18164 13780 18216
rect 11704 18096 11756 18148
rect 15108 18309 15117 18343
rect 15117 18309 15151 18343
rect 15151 18309 15160 18343
rect 15108 18300 15160 18309
rect 15568 18377 15577 18411
rect 15577 18377 15611 18411
rect 15611 18377 15620 18411
rect 15568 18368 15620 18377
rect 16396 18368 16448 18420
rect 20536 18368 20588 18420
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 18328 18300 18380 18352
rect 19064 18232 19116 18284
rect 20720 18232 20772 18284
rect 14648 18164 14700 18216
rect 15108 18164 15160 18216
rect 15752 18164 15804 18216
rect 16304 18164 16356 18216
rect 17408 18164 17460 18216
rect 11888 18028 11940 18080
rect 12992 18028 13044 18080
rect 14004 18028 14056 18080
rect 17316 18096 17368 18148
rect 17224 18028 17276 18080
rect 19708 18028 19760 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 2872 17824 2924 17876
rect 2596 17756 2648 17808
rect 4068 17688 4120 17740
rect 4436 17731 4488 17740
rect 2504 17620 2556 17672
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 6368 17824 6420 17876
rect 6644 17824 6696 17876
rect 9864 17824 9916 17876
rect 4712 17663 4764 17672
rect 4712 17629 4746 17663
rect 4746 17629 4764 17663
rect 4712 17620 4764 17629
rect 4988 17552 5040 17604
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 12900 17824 12952 17876
rect 11060 17756 11112 17808
rect 14004 17824 14056 17876
rect 14372 17824 14424 17876
rect 14832 17824 14884 17876
rect 15200 17824 15252 17876
rect 16488 17824 16540 17876
rect 17132 17824 17184 17876
rect 18236 17867 18288 17876
rect 18236 17833 18245 17867
rect 18245 17833 18279 17867
rect 18279 17833 18288 17867
rect 18236 17824 18288 17833
rect 20628 17824 20680 17876
rect 17040 17756 17092 17808
rect 2596 17484 2648 17536
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 3332 17484 3384 17536
rect 6736 17552 6788 17604
rect 6828 17552 6880 17604
rect 9772 17620 9824 17672
rect 13360 17731 13412 17740
rect 13360 17697 13369 17731
rect 13369 17697 13403 17731
rect 13403 17697 13412 17731
rect 13544 17731 13596 17740
rect 13360 17688 13412 17697
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 16120 17688 16172 17740
rect 16488 17731 16540 17740
rect 8300 17484 8352 17536
rect 10692 17552 10744 17604
rect 11980 17552 12032 17604
rect 13176 17552 13228 17604
rect 16488 17697 16497 17731
rect 16497 17697 16531 17731
rect 16531 17697 16540 17731
rect 19892 17756 19944 17808
rect 17776 17731 17828 17740
rect 16488 17688 16540 17697
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 18788 17731 18840 17740
rect 18788 17697 18797 17731
rect 18797 17697 18831 17731
rect 18831 17697 18840 17731
rect 18788 17688 18840 17697
rect 19800 17731 19852 17740
rect 19800 17697 19809 17731
rect 19809 17697 19843 17731
rect 19843 17697 19852 17731
rect 19800 17688 19852 17697
rect 16672 17663 16724 17672
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 11244 17484 11296 17536
rect 13820 17484 13872 17536
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14464 17484 14516 17493
rect 14832 17484 14884 17536
rect 15016 17484 15068 17536
rect 16120 17484 16172 17536
rect 18420 17552 18472 17604
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 18328 17484 18380 17536
rect 19156 17484 19208 17536
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 21180 17484 21232 17536
rect 22468 17484 22520 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 2780 17280 2832 17332
rect 3332 17280 3384 17332
rect 2228 17144 2280 17196
rect 3332 17144 3384 17196
rect 4252 17144 4304 17196
rect 5632 17144 5684 17196
rect 5908 17187 5960 17196
rect 5908 17153 5926 17187
rect 5926 17153 5960 17187
rect 5908 17144 5960 17153
rect 6276 17144 6328 17196
rect 7288 17280 7340 17332
rect 7380 17280 7432 17332
rect 9220 17280 9272 17332
rect 9772 17323 9824 17332
rect 9772 17289 9781 17323
rect 9781 17289 9815 17323
rect 9815 17289 9824 17323
rect 9772 17280 9824 17289
rect 9864 17280 9916 17332
rect 10048 17212 10100 17264
rect 10232 17280 10284 17332
rect 10876 17280 10928 17332
rect 11152 17280 11204 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 17408 17280 17460 17332
rect 17592 17280 17644 17332
rect 18328 17323 18380 17332
rect 18328 17289 18337 17323
rect 18337 17289 18371 17323
rect 18371 17289 18380 17323
rect 18328 17280 18380 17289
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 19616 17280 19668 17332
rect 20444 17280 20496 17332
rect 21364 17323 21416 17332
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 11888 17212 11940 17264
rect 12992 17255 13044 17264
rect 12992 17221 13001 17255
rect 13001 17221 13035 17255
rect 13035 17221 13044 17255
rect 12992 17212 13044 17221
rect 7840 17144 7892 17196
rect 8024 17144 8076 17196
rect 8668 17144 8720 17196
rect 9772 17144 9824 17196
rect 11704 17144 11756 17196
rect 12808 17144 12860 17196
rect 13268 17212 13320 17264
rect 15292 17212 15344 17264
rect 16212 17255 16264 17264
rect 16212 17221 16221 17255
rect 16221 17221 16255 17255
rect 16255 17221 16264 17255
rect 16212 17212 16264 17221
rect 18604 17212 18656 17264
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 13912 17144 13964 17153
rect 14096 17144 14148 17196
rect 16488 17187 16540 17196
rect 16488 17153 16497 17187
rect 16497 17153 16531 17187
rect 16531 17153 16540 17187
rect 16488 17144 16540 17153
rect 18512 17144 18564 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 20260 17144 20312 17196
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 6828 16940 6880 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 12440 17008 12492 17060
rect 17040 17119 17092 17128
rect 17040 17085 17049 17119
rect 17049 17085 17083 17119
rect 17083 17085 17092 17119
rect 17040 17076 17092 17085
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 18144 17076 18196 17128
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12992 16940 13044 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 19800 17119 19852 17128
rect 19800 17085 19809 17119
rect 19809 17085 19843 17119
rect 19843 17085 19852 17119
rect 19800 17076 19852 17085
rect 20536 17076 20588 17128
rect 19248 17008 19300 17060
rect 21088 17008 21140 17060
rect 17868 16940 17920 16992
rect 18972 16940 19024 16992
rect 20260 16983 20312 16992
rect 20260 16949 20269 16983
rect 20269 16949 20303 16983
rect 20303 16949 20312 16983
rect 20260 16940 20312 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 6276 16779 6328 16788
rect 1676 16600 1728 16652
rect 2596 16532 2648 16584
rect 3056 16600 3108 16652
rect 4068 16600 4120 16652
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 6920 16736 6972 16788
rect 8668 16736 8720 16788
rect 9220 16668 9272 16720
rect 11152 16668 11204 16720
rect 13728 16668 13780 16720
rect 15936 16668 15988 16720
rect 4436 16532 4488 16584
rect 4528 16532 4580 16584
rect 11060 16600 11112 16652
rect 13820 16600 13872 16652
rect 14556 16600 14608 16652
rect 16488 16736 16540 16788
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 18696 16736 18748 16788
rect 17960 16668 18012 16720
rect 18972 16711 19024 16720
rect 18972 16677 18981 16711
rect 18981 16677 19015 16711
rect 19015 16677 19024 16711
rect 18972 16668 19024 16677
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 2964 16464 3016 16516
rect 4252 16507 4304 16516
rect 4252 16473 4261 16507
rect 4261 16473 4295 16507
rect 4295 16473 4304 16507
rect 4252 16464 4304 16473
rect 2872 16396 2924 16448
rect 3332 16396 3384 16448
rect 4988 16507 5040 16516
rect 4988 16473 5022 16507
rect 5022 16473 5040 16507
rect 4988 16464 5040 16473
rect 8024 16464 8076 16516
rect 4436 16396 4488 16448
rect 7012 16396 7064 16448
rect 7840 16396 7892 16448
rect 9772 16396 9824 16448
rect 12164 16532 12216 16584
rect 14464 16532 14516 16584
rect 14924 16532 14976 16584
rect 15292 16532 15344 16584
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 10784 16396 10836 16448
rect 12440 16464 12492 16516
rect 15200 16464 15252 16516
rect 17316 16600 17368 16652
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 15108 16396 15160 16448
rect 16304 16396 16356 16448
rect 16396 16396 16448 16448
rect 16948 16464 17000 16516
rect 17316 16396 17368 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2320 16192 2372 16244
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 2412 16056 2464 16108
rect 5908 16192 5960 16244
rect 4252 16124 4304 16176
rect 9588 16192 9640 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 14464 16235 14516 16244
rect 3148 16056 3200 16108
rect 5724 16099 5776 16108
rect 5724 16065 5742 16099
rect 5742 16065 5776 16099
rect 5724 16056 5776 16065
rect 6920 16056 6972 16108
rect 7012 16056 7064 16108
rect 7840 16124 7892 16176
rect 10324 16124 10376 16176
rect 12164 16124 12216 16176
rect 14464 16201 14473 16235
rect 14473 16201 14507 16235
rect 14507 16201 14516 16235
rect 14464 16192 14516 16201
rect 15108 16192 15160 16244
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 16396 16192 16448 16244
rect 17684 16192 17736 16244
rect 17960 16235 18012 16244
rect 9772 16056 9824 16108
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 10232 16099 10284 16108
rect 10232 16065 10266 16099
rect 10266 16065 10284 16099
rect 10232 16056 10284 16065
rect 12348 16056 12400 16108
rect 12624 16099 12676 16108
rect 12624 16065 12642 16099
rect 12642 16065 12676 16099
rect 12624 16056 12676 16065
rect 1952 15852 2004 15904
rect 3424 15852 3476 15904
rect 9680 15988 9732 16040
rect 15200 16124 15252 16176
rect 17592 16124 17644 16176
rect 17960 16201 17969 16235
rect 17969 16201 18003 16235
rect 18003 16201 18012 16235
rect 17960 16192 18012 16201
rect 20720 16167 20772 16176
rect 20720 16133 20729 16167
rect 20729 16133 20763 16167
rect 20763 16133 20772 16167
rect 20720 16124 20772 16133
rect 15660 16056 15712 16108
rect 16028 16056 16080 16108
rect 16488 16056 16540 16108
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17960 16056 18012 16108
rect 19616 16056 19668 16108
rect 4252 15963 4304 15972
rect 4252 15929 4261 15963
rect 4261 15929 4295 15963
rect 4295 15929 4304 15963
rect 4252 15920 4304 15929
rect 4804 15920 4856 15972
rect 4344 15852 4396 15904
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 4988 15852 5040 15904
rect 5356 15852 5408 15904
rect 7932 15852 7984 15904
rect 8116 15852 8168 15904
rect 9220 15852 9272 15904
rect 11704 15920 11756 15972
rect 15936 16031 15988 16040
rect 15936 15997 15945 16031
rect 15945 15997 15979 16031
rect 15979 15997 15988 16031
rect 15936 15988 15988 15997
rect 16856 15988 16908 16040
rect 17316 16031 17368 16040
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 18236 15988 18288 16040
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 11888 15852 11940 15904
rect 17408 15920 17460 15972
rect 15568 15852 15620 15904
rect 15660 15852 15712 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 4528 15648 4580 15700
rect 6920 15648 6972 15700
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 5356 15444 5408 15496
rect 9956 15648 10008 15700
rect 10232 15580 10284 15632
rect 7104 15444 7156 15496
rect 9220 15487 9272 15496
rect 9220 15453 9254 15487
rect 9254 15453 9272 15487
rect 9220 15444 9272 15453
rect 11888 15444 11940 15496
rect 2136 15376 2188 15428
rect 4344 15376 4396 15428
rect 5632 15376 5684 15428
rect 6460 15376 6512 15428
rect 7656 15376 7708 15428
rect 3976 15308 4028 15360
rect 7012 15308 7064 15360
rect 9312 15308 9364 15360
rect 9588 15308 9640 15360
rect 10692 15376 10744 15428
rect 12624 15648 12676 15700
rect 13820 15648 13872 15700
rect 14832 15648 14884 15700
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 15568 15648 15620 15700
rect 16396 15648 16448 15700
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 17408 15691 17460 15700
rect 17408 15657 17417 15691
rect 17417 15657 17451 15691
rect 17451 15657 17460 15691
rect 17408 15648 17460 15657
rect 13728 15580 13780 15632
rect 12624 15512 12676 15564
rect 16488 15555 16540 15564
rect 12348 15444 12400 15496
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 16580 15512 16632 15564
rect 17040 15444 17092 15496
rect 17224 15444 17276 15496
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 20536 15555 20588 15564
rect 20536 15521 20545 15555
rect 20545 15521 20579 15555
rect 20579 15521 20588 15555
rect 20536 15512 20588 15521
rect 13820 15419 13872 15428
rect 11520 15308 11572 15360
rect 12256 15308 12308 15360
rect 13268 15308 13320 15360
rect 13820 15385 13829 15419
rect 13829 15385 13863 15419
rect 13863 15385 13872 15419
rect 13820 15376 13872 15385
rect 14832 15419 14884 15428
rect 14832 15385 14841 15419
rect 14841 15385 14875 15419
rect 14875 15385 14884 15419
rect 14832 15376 14884 15385
rect 15476 15376 15528 15428
rect 15660 15419 15712 15428
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 16948 15376 17000 15428
rect 20536 15376 20588 15428
rect 15936 15308 15988 15360
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 17040 15308 17092 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 18880 15308 18932 15360
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 19708 15308 19760 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 3240 15104 3292 15156
rect 3792 15079 3844 15088
rect 3792 15045 3801 15079
rect 3801 15045 3835 15079
rect 3835 15045 3844 15079
rect 3792 15036 3844 15045
rect 4528 15036 4580 15088
rect 6920 15104 6972 15156
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 4252 14968 4304 15020
rect 4068 14900 4120 14952
rect 4804 14832 4856 14884
rect 7012 14832 7064 14884
rect 5816 14764 5868 14816
rect 7656 14764 7708 14816
rect 9312 15104 9364 15156
rect 9956 15104 10008 15156
rect 7932 15036 7984 15088
rect 13268 15104 13320 15156
rect 15108 15104 15160 15156
rect 16948 15104 17000 15156
rect 19064 15104 19116 15156
rect 19524 15104 19576 15156
rect 19708 15147 19760 15156
rect 19708 15113 19717 15147
rect 19717 15113 19751 15147
rect 19751 15113 19760 15147
rect 19708 15104 19760 15113
rect 20352 15104 20404 15156
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 8116 15011 8168 15020
rect 8116 14977 8150 15011
rect 8150 14977 8168 15011
rect 8116 14968 8168 14977
rect 8576 14968 8628 15020
rect 9220 14900 9272 14952
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 11060 14832 11112 14884
rect 8576 14764 8628 14816
rect 10968 14764 11020 14816
rect 12992 14900 13044 14952
rect 14004 14968 14056 15020
rect 15292 15036 15344 15088
rect 16304 15036 16356 15088
rect 14188 14900 14240 14952
rect 14648 14900 14700 14952
rect 15108 14900 15160 14952
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 16396 14943 16448 14952
rect 14648 14764 14700 14816
rect 15200 14764 15252 14816
rect 16396 14909 16405 14943
rect 16405 14909 16439 14943
rect 16439 14909 16448 14943
rect 16396 14900 16448 14909
rect 17684 15036 17736 15088
rect 18236 15036 18288 15088
rect 19984 15036 20036 15088
rect 20536 15036 20588 15088
rect 17316 14968 17368 15020
rect 19064 14968 19116 15020
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 20352 14968 20404 15020
rect 21180 15011 21232 15020
rect 21180 14977 21189 15011
rect 21189 14977 21223 15011
rect 21223 14977 21232 15011
rect 21180 14968 21232 14977
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 17592 14832 17644 14884
rect 17224 14764 17276 14816
rect 17868 14764 17920 14816
rect 18788 14807 18840 14816
rect 18788 14773 18797 14807
rect 18797 14773 18831 14807
rect 18831 14773 18840 14807
rect 18788 14764 18840 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 4160 14560 4212 14612
rect 5448 14560 5500 14612
rect 3332 14467 3384 14476
rect 3332 14433 3341 14467
rect 3341 14433 3375 14467
rect 3375 14433 3384 14467
rect 3332 14424 3384 14433
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 6920 14560 6972 14612
rect 7472 14424 7524 14476
rect 7748 14424 7800 14476
rect 9956 14560 10008 14612
rect 10968 14560 11020 14612
rect 10876 14492 10928 14544
rect 12440 14560 12492 14612
rect 12532 14560 12584 14612
rect 15384 14560 15436 14612
rect 18328 14560 18380 14612
rect 20628 14560 20680 14612
rect 13636 14535 13688 14544
rect 13636 14501 13645 14535
rect 13645 14501 13679 14535
rect 13679 14501 13688 14535
rect 13636 14492 13688 14501
rect 15108 14492 15160 14544
rect 16028 14492 16080 14544
rect 16396 14492 16448 14544
rect 5816 14356 5868 14408
rect 6552 14356 6604 14408
rect 11428 14424 11480 14476
rect 14372 14424 14424 14476
rect 10968 14356 11020 14408
rect 12808 14356 12860 14408
rect 14832 14424 14884 14476
rect 16212 14424 16264 14476
rect 20536 14492 20588 14544
rect 17500 14424 17552 14476
rect 18144 14424 18196 14476
rect 5356 14288 5408 14340
rect 5448 14288 5500 14340
rect 2964 14220 3016 14272
rect 3240 14263 3292 14272
rect 3240 14229 3249 14263
rect 3249 14229 3283 14263
rect 3283 14229 3292 14263
rect 3240 14220 3292 14229
rect 4344 14220 4396 14272
rect 8392 14288 8444 14340
rect 10324 14288 10376 14340
rect 10508 14288 10560 14340
rect 12348 14288 12400 14340
rect 12900 14288 12952 14340
rect 8116 14220 8168 14272
rect 10048 14220 10100 14272
rect 10876 14220 10928 14272
rect 11428 14220 11480 14272
rect 18052 14356 18104 14408
rect 18236 14356 18288 14408
rect 18604 14424 18656 14476
rect 21180 14424 21232 14476
rect 18788 14356 18840 14408
rect 13636 14220 13688 14272
rect 15200 14220 15252 14272
rect 18144 14220 18196 14272
rect 18696 14220 18748 14272
rect 20628 14220 20680 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2780 14016 2832 14068
rect 3424 14016 3476 14068
rect 4068 14016 4120 14068
rect 1952 13880 2004 13932
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 5540 13948 5592 14000
rect 7472 14016 7524 14068
rect 5816 13948 5868 14000
rect 9220 14016 9272 14068
rect 3976 13880 4028 13932
rect 8576 13948 8628 14000
rect 9956 14016 10008 14068
rect 11152 14016 11204 14068
rect 12440 14016 12492 14068
rect 16580 14016 16632 14068
rect 17408 14016 17460 14068
rect 18604 14016 18656 14068
rect 19892 14016 19944 14068
rect 20076 14016 20128 14068
rect 20628 14059 20680 14068
rect 20628 14025 20637 14059
rect 20637 14025 20671 14059
rect 20671 14025 20680 14059
rect 20628 14016 20680 14025
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 8392 13880 8444 13932
rect 10048 13948 10100 14000
rect 14372 13948 14424 14000
rect 16396 13948 16448 14000
rect 18052 13991 18104 14000
rect 10508 13880 10560 13932
rect 10968 13880 11020 13932
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 5172 13676 5224 13728
rect 6368 13787 6420 13796
rect 6368 13753 6377 13787
rect 6377 13753 6411 13787
rect 6411 13753 6420 13787
rect 6368 13744 6420 13753
rect 9496 13812 9548 13864
rect 11244 13812 11296 13864
rect 12164 13880 12216 13932
rect 18052 13957 18061 13991
rect 18061 13957 18095 13991
rect 18095 13957 18104 13991
rect 18052 13948 18104 13957
rect 19708 13948 19760 14000
rect 18696 13880 18748 13932
rect 19432 13880 19484 13932
rect 20812 13948 20864 14000
rect 12900 13812 12952 13864
rect 17592 13812 17644 13864
rect 18972 13855 19024 13864
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 20444 13812 20496 13864
rect 12808 13744 12860 13796
rect 17776 13744 17828 13796
rect 20628 13744 20680 13796
rect 21272 13812 21324 13864
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 18052 13676 18104 13728
rect 18696 13676 18748 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 5080 13472 5132 13524
rect 7564 13472 7616 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9956 13472 10008 13524
rect 2780 13404 2832 13456
rect 3148 13404 3200 13456
rect 6828 13404 6880 13456
rect 15752 13472 15804 13524
rect 17132 13472 17184 13524
rect 17316 13472 17368 13524
rect 17776 13472 17828 13524
rect 19064 13472 19116 13524
rect 19984 13472 20036 13524
rect 12716 13404 12768 13456
rect 12992 13404 13044 13456
rect 18052 13404 18104 13456
rect 10968 13336 11020 13388
rect 12164 13336 12216 13388
rect 15752 13336 15804 13388
rect 16580 13379 16632 13388
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 16580 13336 16632 13345
rect 3148 13268 3200 13320
rect 3884 13268 3936 13320
rect 9312 13268 9364 13320
rect 12256 13268 12308 13320
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 15844 13268 15896 13320
rect 16304 13268 16356 13320
rect 17408 13268 17460 13320
rect 5172 13200 5224 13252
rect 5632 13132 5684 13184
rect 9588 13200 9640 13252
rect 11980 13200 12032 13252
rect 17776 13336 17828 13388
rect 18512 13404 18564 13456
rect 19524 13336 19576 13388
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 20444 13336 20496 13388
rect 20536 13336 20588 13388
rect 18696 13200 18748 13252
rect 20812 13200 20864 13252
rect 8668 13132 8720 13184
rect 12532 13132 12584 13184
rect 15844 13132 15896 13184
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 17316 13132 17368 13184
rect 17408 13132 17460 13184
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 19432 13132 19484 13184
rect 20260 13132 20312 13184
rect 20536 13175 20588 13184
rect 20536 13141 20545 13175
rect 20545 13141 20579 13175
rect 20579 13141 20588 13175
rect 20536 13132 20588 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2596 12928 2648 12980
rect 6736 12928 6788 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 7012 12860 7064 12912
rect 2044 12792 2096 12844
rect 4988 12792 5040 12844
rect 6828 12835 6880 12844
rect 6828 12801 6862 12835
rect 6862 12801 6880 12835
rect 6828 12792 6880 12801
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 5172 12588 5224 12640
rect 9956 12928 10008 12980
rect 11060 12928 11112 12980
rect 10876 12860 10928 12912
rect 10968 12860 11020 12912
rect 12532 12928 12584 12980
rect 13636 12928 13688 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17776 12928 17828 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20260 12971 20312 12980
rect 20260 12937 20269 12971
rect 20269 12937 20303 12971
rect 20303 12937 20312 12971
rect 20260 12928 20312 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 10692 12792 10744 12844
rect 13544 12903 13596 12912
rect 13544 12869 13553 12903
rect 13553 12869 13587 12903
rect 13587 12869 13596 12903
rect 13544 12860 13596 12869
rect 15568 12860 15620 12912
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 16120 12860 16172 12912
rect 18052 12860 18104 12912
rect 12808 12656 12860 12708
rect 15752 12724 15804 12776
rect 16212 12724 16264 12776
rect 17776 12792 17828 12844
rect 18420 12792 18472 12844
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19800 12835 19852 12844
rect 16948 12656 17000 12708
rect 11244 12588 11296 12640
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 15660 12588 15712 12640
rect 17592 12724 17644 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 17868 12656 17920 12708
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 19524 12724 19576 12776
rect 20352 12588 20404 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 3424 12384 3476 12436
rect 5724 12316 5776 12368
rect 10968 12384 11020 12436
rect 14280 12384 14332 12436
rect 14740 12384 14792 12436
rect 14464 12316 14516 12368
rect 9956 12248 10008 12300
rect 5172 12180 5224 12232
rect 10968 12180 11020 12232
rect 12808 12248 12860 12300
rect 14372 12248 14424 12300
rect 15200 12384 15252 12436
rect 17868 12427 17920 12436
rect 17868 12393 17877 12427
rect 17877 12393 17911 12427
rect 17911 12393 17920 12427
rect 17868 12384 17920 12393
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 21456 12384 21508 12436
rect 15476 12316 15528 12368
rect 16212 12316 16264 12368
rect 17316 12316 17368 12368
rect 20260 12316 20312 12368
rect 22376 12316 22428 12368
rect 15752 12248 15804 12300
rect 16396 12180 16448 12232
rect 17500 12248 17552 12300
rect 18052 12248 18104 12300
rect 18972 12248 19024 12300
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 20628 12248 20680 12300
rect 17684 12180 17736 12232
rect 19524 12180 19576 12232
rect 4252 12112 4304 12164
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 5632 12044 5684 12096
rect 5816 12044 5868 12096
rect 7472 12112 7524 12164
rect 9036 12112 9088 12164
rect 11060 12112 11112 12164
rect 12532 12112 12584 12164
rect 16948 12112 17000 12164
rect 18880 12112 18932 12164
rect 19432 12112 19484 12164
rect 21272 12112 21324 12164
rect 9496 12044 9548 12096
rect 9956 12044 10008 12096
rect 10784 12044 10836 12096
rect 11796 12044 11848 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 14740 12044 14792 12096
rect 15384 12044 15436 12096
rect 15660 12044 15712 12096
rect 16028 12044 16080 12096
rect 18052 12044 18104 12096
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 18696 12044 18748 12096
rect 20352 12044 20404 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1952 11815 2004 11824
rect 1952 11781 1961 11815
rect 1961 11781 1995 11815
rect 1995 11781 2004 11815
rect 1952 11772 2004 11781
rect 1768 11704 1820 11756
rect 3056 11840 3108 11892
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 5540 11840 5592 11892
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 9128 11840 9180 11892
rect 10968 11840 11020 11892
rect 13544 11883 13596 11892
rect 7840 11704 7892 11756
rect 8484 11704 8536 11756
rect 9496 11704 9548 11756
rect 9772 11747 9824 11756
rect 9772 11713 9801 11747
rect 9801 11713 9824 11747
rect 9772 11704 9824 11713
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 10968 11704 11020 11756
rect 12164 11772 12216 11824
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 15016 11883 15068 11892
rect 15016 11849 15025 11883
rect 15025 11849 15059 11883
rect 15059 11849 15068 11883
rect 15016 11840 15068 11849
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 16396 11840 16448 11892
rect 11796 11747 11848 11756
rect 11796 11713 11830 11747
rect 11830 11713 11848 11747
rect 11796 11704 11848 11713
rect 12716 11704 12768 11756
rect 13820 11772 13872 11824
rect 17224 11840 17276 11892
rect 18328 11840 18380 11892
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 20812 11883 20864 11892
rect 20812 11849 20821 11883
rect 20821 11849 20855 11883
rect 20855 11849 20864 11883
rect 20812 11840 20864 11849
rect 20996 11840 21048 11892
rect 14280 11747 14332 11756
rect 12900 11636 12952 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 18052 11772 18104 11824
rect 18696 11772 18748 11824
rect 19800 11772 19852 11824
rect 20260 11772 20312 11824
rect 17960 11704 18012 11756
rect 19616 11747 19668 11756
rect 5448 11568 5500 11620
rect 7472 11568 7524 11620
rect 2780 11500 2832 11552
rect 4252 11500 4304 11552
rect 6644 11500 6696 11552
rect 9036 11500 9088 11552
rect 11520 11568 11572 11620
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 16396 11636 16448 11688
rect 18052 11636 18104 11688
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 10324 11500 10376 11552
rect 17040 11568 17092 11620
rect 17776 11568 17828 11620
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 20812 11704 20864 11756
rect 19708 11636 19760 11688
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 20260 11568 20312 11620
rect 12992 11500 13044 11552
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 15200 11500 15252 11552
rect 17500 11500 17552 11552
rect 17684 11500 17736 11552
rect 19616 11500 19668 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2872 11296 2924 11348
rect 3792 11296 3844 11348
rect 8852 11296 8904 11348
rect 3148 11228 3200 11280
rect 7196 11271 7248 11280
rect 7196 11237 7205 11271
rect 7205 11237 7239 11271
rect 7239 11237 7248 11271
rect 7196 11228 7248 11237
rect 10968 11339 11020 11348
rect 10968 11305 10977 11339
rect 10977 11305 11011 11339
rect 11011 11305 11020 11339
rect 10968 11296 11020 11305
rect 11060 11296 11112 11348
rect 17040 11339 17092 11348
rect 10324 11271 10376 11280
rect 10324 11237 10333 11271
rect 10333 11237 10367 11271
rect 10367 11237 10376 11271
rect 10324 11228 10376 11237
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 12532 11271 12584 11280
rect 12532 11237 12541 11271
rect 12541 11237 12575 11271
rect 12575 11237 12584 11271
rect 12532 11228 12584 11237
rect 12900 11271 12952 11280
rect 12900 11237 12909 11271
rect 12909 11237 12943 11271
rect 12943 11237 12952 11271
rect 12900 11228 12952 11237
rect 13544 11228 13596 11280
rect 13820 11228 13872 11280
rect 12716 11160 12768 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 16212 11228 16264 11280
rect 15476 11160 15528 11212
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 18236 11296 18288 11348
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 6920 11092 6972 11144
rect 9496 11092 9548 11144
rect 4252 11024 4304 11076
rect 5632 11024 5684 11076
rect 5908 11024 5960 11076
rect 7196 11024 7248 11076
rect 7840 11024 7892 11076
rect 10692 11024 10744 11076
rect 9772 10956 9824 11008
rect 9864 10956 9916 11008
rect 10140 10956 10192 11008
rect 10508 10956 10560 11008
rect 11244 11024 11296 11076
rect 11704 11024 11756 11076
rect 11152 10956 11204 11008
rect 11888 10956 11940 11008
rect 12440 11092 12492 11144
rect 16028 11092 16080 11144
rect 16120 11092 16172 11144
rect 17316 11092 17368 11144
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18512 11092 18564 11144
rect 12072 11024 12124 11076
rect 15660 11024 15712 11076
rect 18328 11067 18380 11076
rect 18328 11033 18337 11067
rect 18337 11033 18371 11067
rect 18371 11033 18380 11067
rect 18328 11024 18380 11033
rect 19064 11296 19116 11348
rect 20536 11296 20588 11348
rect 19800 11228 19852 11280
rect 20628 11228 20680 11280
rect 18880 11160 18932 11212
rect 20168 11160 20220 11212
rect 20536 11092 20588 11144
rect 20812 11092 20864 11144
rect 19064 11024 19116 11076
rect 13084 10956 13136 11008
rect 15844 10999 15896 11008
rect 15844 10965 15853 10999
rect 15853 10965 15887 10999
rect 15887 10965 15896 10999
rect 15844 10956 15896 10965
rect 16028 10956 16080 11008
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 19984 10956 20036 11008
rect 20812 10956 20864 11008
rect 20996 10999 21048 11008
rect 20996 10965 21005 10999
rect 21005 10965 21039 10999
rect 21039 10965 21048 10999
rect 20996 10956 21048 10965
rect 21456 10999 21508 11008
rect 21456 10965 21465 10999
rect 21465 10965 21499 10999
rect 21499 10965 21508 10999
rect 21456 10956 21508 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 3884 10752 3936 10804
rect 10508 10752 10560 10804
rect 10784 10752 10836 10804
rect 3424 10616 3476 10668
rect 5724 10684 5776 10736
rect 5356 10616 5408 10668
rect 6828 10616 6880 10668
rect 9864 10616 9916 10668
rect 10968 10684 11020 10736
rect 13268 10752 13320 10804
rect 13820 10752 13872 10804
rect 14832 10752 14884 10804
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 15936 10752 15988 10804
rect 20996 10752 21048 10804
rect 10232 10659 10284 10668
rect 10232 10625 10266 10659
rect 10266 10625 10284 10659
rect 10232 10616 10284 10625
rect 10692 10616 10744 10668
rect 11152 10616 11204 10668
rect 11888 10616 11940 10668
rect 12348 10616 12400 10668
rect 12808 10616 12860 10668
rect 12992 10616 13044 10668
rect 15568 10684 15620 10736
rect 16856 10616 16908 10668
rect 17960 10616 18012 10668
rect 19524 10684 19576 10736
rect 20168 10684 20220 10736
rect 19616 10616 19668 10668
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 22468 10616 22520 10668
rect 16488 10548 16540 10600
rect 16580 10548 16632 10600
rect 17776 10548 17828 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 9496 10480 9548 10532
rect 2780 10412 2832 10464
rect 5448 10412 5500 10464
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 7748 10412 7800 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 11060 10412 11112 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 17224 10480 17276 10532
rect 19892 10480 19944 10532
rect 12992 10412 13044 10421
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 18052 10412 18104 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2688 10251 2740 10260
rect 2688 10217 2697 10251
rect 2697 10217 2731 10251
rect 2731 10217 2740 10251
rect 2688 10208 2740 10217
rect 2872 10208 2924 10260
rect 6920 10251 6972 10260
rect 3976 10072 4028 10124
rect 4160 10004 4212 10056
rect 4528 10004 4580 10056
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 6000 10004 6052 10056
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 6552 10140 6604 10192
rect 10968 10208 11020 10260
rect 12808 10251 12860 10260
rect 10140 10140 10192 10192
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 12992 10208 13044 10260
rect 14372 10208 14424 10260
rect 15292 10208 15344 10260
rect 16396 10208 16448 10260
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 17960 10251 18012 10260
rect 16948 10208 17000 10217
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 19984 10208 20036 10260
rect 21088 10208 21140 10260
rect 17132 10140 17184 10192
rect 12808 10072 12860 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 14096 10072 14148 10124
rect 14648 10072 14700 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 16120 10072 16172 10124
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 10508 10004 10560 10056
rect 10876 10047 10928 10056
rect 10876 10013 10905 10047
rect 10905 10013 10928 10047
rect 10876 10004 10928 10013
rect 15200 10004 15252 10056
rect 19708 10140 19760 10192
rect 20444 10140 20496 10192
rect 20536 10140 20588 10192
rect 18144 10072 18196 10124
rect 19524 10072 19576 10124
rect 19616 10072 19668 10124
rect 19892 10072 19944 10124
rect 5540 9936 5592 9988
rect 2596 9868 2648 9920
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3516 9868 3568 9920
rect 3976 9868 4028 9920
rect 6828 9868 6880 9920
rect 10048 9936 10100 9988
rect 13084 9936 13136 9988
rect 13820 9936 13872 9988
rect 9496 9868 9548 9920
rect 10416 9868 10468 9920
rect 10508 9868 10560 9920
rect 11060 9868 11112 9920
rect 11796 9868 11848 9920
rect 12716 9868 12768 9920
rect 12900 9868 12952 9920
rect 14740 9936 14792 9988
rect 14924 9911 14976 9920
rect 14924 9877 14933 9911
rect 14933 9877 14967 9911
rect 14967 9877 14976 9911
rect 15292 9911 15344 9920
rect 14924 9868 14976 9877
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 16120 9868 16172 9920
rect 17592 9936 17644 9988
rect 19616 9979 19668 9988
rect 19616 9945 19625 9979
rect 19625 9945 19659 9979
rect 19659 9945 19668 9979
rect 19616 9936 19668 9945
rect 17868 9911 17920 9920
rect 17868 9877 17877 9911
rect 17877 9877 17911 9911
rect 17911 9877 17920 9911
rect 17868 9868 17920 9877
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 19708 9868 19760 9920
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 20444 10004 20496 10056
rect 20812 9868 20864 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 3056 9664 3108 9716
rect 4252 9707 4304 9716
rect 4252 9673 4261 9707
rect 4261 9673 4295 9707
rect 4295 9673 4304 9707
rect 4252 9664 4304 9673
rect 4436 9664 4488 9716
rect 4712 9664 4764 9716
rect 5356 9664 5408 9716
rect 3700 9639 3752 9648
rect 3700 9605 3709 9639
rect 3709 9605 3743 9639
rect 3743 9605 3752 9639
rect 3700 9596 3752 9605
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2688 9528 2740 9580
rect 1676 9460 1728 9512
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 2780 9460 2832 9512
rect 3056 9460 3108 9512
rect 5540 9596 5592 9648
rect 4436 9528 4488 9580
rect 5448 9571 5500 9580
rect 4160 9392 4212 9444
rect 4620 9460 4672 9512
rect 4712 9460 4764 9512
rect 4988 9460 5040 9512
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 6000 9664 6052 9716
rect 6552 9664 6604 9716
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7012 9528 7064 9580
rect 10968 9664 11020 9716
rect 12348 9664 12400 9716
rect 14096 9664 14148 9716
rect 14924 9664 14976 9716
rect 15200 9664 15252 9716
rect 18144 9664 18196 9716
rect 18420 9664 18472 9716
rect 19616 9664 19668 9716
rect 9864 9639 9916 9648
rect 9864 9605 9898 9639
rect 9898 9605 9916 9639
rect 9864 9596 9916 9605
rect 5632 9392 5684 9444
rect 6920 9392 6972 9444
rect 2780 9324 2832 9376
rect 3516 9324 3568 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 8392 9324 8444 9376
rect 9128 9324 9180 9376
rect 12624 9571 12676 9580
rect 12624 9537 12642 9571
rect 12642 9537 12676 9571
rect 12624 9528 12676 9537
rect 12808 9528 12860 9580
rect 10876 9324 10928 9376
rect 15292 9596 15344 9648
rect 16948 9596 17000 9648
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 18604 9596 18656 9648
rect 19524 9596 19576 9648
rect 20260 9639 20312 9648
rect 20260 9605 20269 9639
rect 20269 9605 20303 9639
rect 20303 9605 20312 9639
rect 20260 9596 20312 9605
rect 20812 9664 20864 9716
rect 15200 9528 15252 9580
rect 15476 9528 15528 9580
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17408 9528 17460 9580
rect 18880 9528 18932 9580
rect 16396 9503 16448 9512
rect 13728 9392 13780 9444
rect 14832 9392 14884 9444
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 20076 9528 20128 9580
rect 20536 9528 20588 9580
rect 20628 9528 20680 9580
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 17408 9392 17460 9444
rect 20904 9392 20956 9444
rect 21364 9435 21416 9444
rect 21364 9401 21373 9435
rect 21373 9401 21407 9435
rect 21407 9401 21416 9435
rect 21364 9392 21416 9401
rect 13452 9324 13504 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 16396 9324 16448 9376
rect 16856 9324 16908 9376
rect 17592 9324 17644 9376
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 17868 9324 17920 9333
rect 18604 9324 18656 9376
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1860 9120 1912 9172
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3332 9120 3384 9172
rect 4252 9120 4304 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5448 9120 5500 9172
rect 7380 9120 7432 9172
rect 13636 9120 13688 9172
rect 13912 9120 13964 9172
rect 15936 9120 15988 9172
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 3976 9052 4028 9104
rect 9680 9052 9732 9104
rect 10232 9052 10284 9104
rect 5172 8984 5224 9036
rect 5724 8984 5776 9036
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 6828 8984 6880 9036
rect 6920 8984 6972 9036
rect 12532 8984 12584 9036
rect 14280 8984 14332 9036
rect 16488 9052 16540 9104
rect 18420 9120 18472 9172
rect 20076 9120 20128 9172
rect 20260 9120 20312 9172
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 4712 8916 4764 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 12716 8916 12768 8968
rect 13360 8916 13412 8968
rect 3332 8848 3384 8900
rect 3516 8848 3568 8900
rect 4436 8780 4488 8832
rect 4988 8780 5040 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 6552 8780 6604 8832
rect 12808 8780 12860 8832
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 15660 8916 15712 8968
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 19616 9052 19668 9104
rect 17224 8984 17276 9036
rect 18604 8984 18656 9036
rect 18972 8916 19024 8968
rect 19524 8984 19576 9036
rect 20168 9052 20220 9104
rect 20352 9052 20404 9104
rect 20628 9027 20680 9036
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 20628 8993 20637 9027
rect 20637 8993 20671 9027
rect 20671 8993 20680 9027
rect 20628 8984 20680 8993
rect 20812 8916 20864 8968
rect 13820 8848 13872 8900
rect 15108 8848 15160 8900
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 20444 8848 20496 8900
rect 20168 8780 20220 8832
rect 20536 8780 20588 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1400 8576 1452 8628
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 5172 8576 5224 8628
rect 6092 8619 6144 8628
rect 3516 8508 3568 8560
rect 4252 8508 4304 8560
rect 4436 8551 4488 8560
rect 4436 8517 4445 8551
rect 4445 8517 4479 8551
rect 4479 8517 4488 8551
rect 4436 8508 4488 8517
rect 5724 8508 5776 8560
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7748 8576 7800 8628
rect 11152 8576 11204 8628
rect 13728 8619 13780 8628
rect 7012 8508 7064 8560
rect 7656 8508 7708 8560
rect 4068 8440 4120 8492
rect 5080 8440 5132 8492
rect 12716 8440 12768 8492
rect 4620 8372 4672 8424
rect 5172 8372 5224 8424
rect 5264 8372 5316 8424
rect 6092 8372 6144 8424
rect 6460 8415 6512 8424
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 6460 8372 6512 8381
rect 7472 8372 7524 8424
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 18880 8619 18932 8628
rect 13912 8508 13964 8560
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 20720 8576 20772 8628
rect 21640 8576 21692 8628
rect 14556 8508 14608 8560
rect 14740 8508 14792 8560
rect 18604 8508 18656 8560
rect 19432 8508 19484 8560
rect 19892 8508 19944 8560
rect 14096 8440 14148 8492
rect 4344 8304 4396 8356
rect 13728 8372 13780 8424
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 15936 8440 15988 8492
rect 19156 8440 19208 8492
rect 19984 8440 20036 8492
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 15200 8372 15252 8424
rect 3976 8236 4028 8288
rect 15108 8304 15160 8356
rect 17868 8372 17920 8424
rect 19064 8372 19116 8424
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 13544 8236 13596 8288
rect 13636 8236 13688 8288
rect 14648 8236 14700 8288
rect 18604 8236 18656 8288
rect 19984 8279 20036 8288
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 20628 8236 20680 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2044 8032 2096 8084
rect 4068 8032 4120 8084
rect 13636 8032 13688 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 14556 8032 14608 8084
rect 3240 7964 3292 8016
rect 14740 7964 14792 8016
rect 2596 7896 2648 7948
rect 4160 7896 4212 7948
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 5908 7896 5960 7948
rect 6920 7896 6972 7948
rect 10324 7896 10376 7948
rect 13820 7896 13872 7948
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 2688 7828 2740 7880
rect 6552 7828 6604 7880
rect 14464 7896 14516 7948
rect 2044 7692 2096 7744
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 4436 7692 4488 7744
rect 5080 7692 5132 7744
rect 5540 7692 5592 7744
rect 6000 7692 6052 7744
rect 6736 7735 6788 7744
rect 6736 7701 6745 7735
rect 6745 7701 6779 7735
rect 6779 7701 6788 7735
rect 6736 7692 6788 7701
rect 9680 7735 9732 7744
rect 9680 7701 9689 7735
rect 9689 7701 9723 7735
rect 9723 7701 9732 7735
rect 9680 7692 9732 7701
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 12808 7760 12860 7812
rect 18328 8032 18380 8084
rect 18604 8075 18656 8084
rect 18604 8041 18613 8075
rect 18613 8041 18647 8075
rect 18647 8041 18656 8075
rect 18604 8032 18656 8041
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 21548 8032 21600 8084
rect 20352 7964 20404 8016
rect 22100 7964 22152 8016
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 18144 7939 18196 7948
rect 18144 7905 18153 7939
rect 18153 7905 18187 7939
rect 18187 7905 18196 7939
rect 18144 7896 18196 7905
rect 16120 7828 16172 7880
rect 13544 7692 13596 7744
rect 15568 7692 15620 7744
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 18236 7760 18288 7812
rect 19892 7896 19944 7948
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 20076 7896 20128 7948
rect 20812 7871 20864 7880
rect 20812 7837 20821 7871
rect 20821 7837 20855 7871
rect 20855 7837 20864 7871
rect 20812 7828 20864 7837
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 19984 7760 20036 7812
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18972 7735 19024 7744
rect 18972 7701 18981 7735
rect 18981 7701 19015 7735
rect 19015 7701 19024 7735
rect 18972 7692 19024 7701
rect 19616 7692 19668 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2228 7488 2280 7540
rect 4252 7488 4304 7540
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 9772 7488 9824 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 15752 7488 15804 7540
rect 19708 7488 19760 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 21088 7488 21140 7540
rect 3332 7420 3384 7472
rect 12072 7420 12124 7472
rect 18604 7420 18656 7472
rect 18788 7463 18840 7472
rect 18788 7429 18797 7463
rect 18797 7429 18831 7463
rect 18831 7429 18840 7463
rect 18788 7420 18840 7429
rect 20076 7420 20128 7472
rect 3424 7352 3476 7404
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 8300 7352 8352 7404
rect 9404 7352 9456 7404
rect 3332 7284 3384 7336
rect 5264 7284 5316 7336
rect 5080 7216 5132 7268
rect 6000 7216 6052 7268
rect 8668 7284 8720 7336
rect 10140 7284 10192 7336
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11796 7352 11848 7404
rect 17868 7395 17920 7404
rect 14372 7284 14424 7336
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 20812 7420 20864 7472
rect 13176 7216 13228 7268
rect 18236 7284 18288 7336
rect 19248 7284 19300 7336
rect 20260 7216 20312 7268
rect 20720 7284 20772 7336
rect 20628 7216 20680 7268
rect 6736 7191 6788 7200
rect 6736 7157 6745 7191
rect 6745 7157 6779 7191
rect 6779 7157 6788 7191
rect 6736 7148 6788 7157
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 15016 7148 15068 7200
rect 18144 7148 18196 7200
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 18420 7148 18472 7200
rect 19248 7148 19300 7200
rect 19708 7148 19760 7200
rect 20444 7148 20496 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2136 6944 2188 6996
rect 17868 6944 17920 6996
rect 17960 6944 18012 6996
rect 19892 6944 19944 6996
rect 20720 6944 20772 6996
rect 3056 6808 3108 6860
rect 3424 6808 3476 6860
rect 4712 6851 4764 6860
rect 4068 6740 4120 6792
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 7196 6808 7248 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 10784 6808 10836 6860
rect 18420 6808 18472 6860
rect 21180 6876 21232 6928
rect 19524 6808 19576 6860
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 21088 6808 21140 6860
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 3608 6604 3660 6656
rect 18972 6740 19024 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 7012 6604 7064 6656
rect 10508 6604 10560 6656
rect 11704 6604 11756 6656
rect 14464 6604 14516 6656
rect 18144 6604 18196 6656
rect 20168 6604 20220 6656
rect 20352 6604 20404 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2964 6400 3016 6452
rect 3608 6443 3660 6452
rect 3608 6409 3617 6443
rect 3617 6409 3651 6443
rect 3651 6409 3660 6443
rect 3608 6400 3660 6409
rect 3884 6400 3936 6452
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 6736 6400 6788 6452
rect 8300 6400 8352 6452
rect 9680 6400 9732 6452
rect 12072 6443 12124 6452
rect 12072 6409 12081 6443
rect 12081 6409 12115 6443
rect 12115 6409 12124 6443
rect 12072 6400 12124 6409
rect 12440 6400 12492 6452
rect 10784 6375 10836 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 5172 6264 5224 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 8208 6264 8260 6316
rect 10784 6341 10793 6375
rect 10793 6341 10827 6375
rect 10827 6341 10836 6375
rect 10784 6332 10836 6341
rect 12164 6332 12216 6384
rect 12992 6400 13044 6452
rect 17132 6400 17184 6452
rect 18144 6443 18196 6452
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 18328 6400 18380 6452
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 20628 6400 20680 6452
rect 13452 6332 13504 6384
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 2780 6128 2832 6180
rect 4528 6196 4580 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6000 6196 6052 6248
rect 6644 6196 6696 6248
rect 8300 6196 8352 6248
rect 4252 6128 4304 6180
rect 5540 6128 5592 6180
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 13728 6264 13780 6316
rect 12532 6196 12584 6248
rect 8208 6060 8260 6112
rect 12164 6060 12216 6112
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 17408 6239 17460 6248
rect 14464 6196 14516 6205
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 18052 6332 18104 6384
rect 19984 6375 20036 6384
rect 19984 6341 19993 6375
rect 19993 6341 20027 6375
rect 20027 6341 20036 6375
rect 19984 6332 20036 6341
rect 19524 6264 19576 6316
rect 19800 6264 19852 6316
rect 17776 6196 17828 6248
rect 18420 6196 18472 6248
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 15568 6060 15620 6112
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 2964 5856 3016 5908
rect 4068 5856 4120 5908
rect 13820 5856 13872 5908
rect 17408 5856 17460 5908
rect 2504 5788 2556 5840
rect 5540 5788 5592 5840
rect 5632 5788 5684 5840
rect 10784 5788 10836 5840
rect 17960 5788 18012 5840
rect 2780 5720 2832 5772
rect 4528 5720 4580 5772
rect 5724 5720 5776 5772
rect 6644 5720 6696 5772
rect 6828 5720 6880 5772
rect 17776 5720 17828 5772
rect 19892 5720 19944 5772
rect 19984 5720 20036 5772
rect 5356 5652 5408 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 7196 5652 7248 5704
rect 6552 5584 6604 5636
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 3792 5516 3844 5568
rect 3976 5516 4028 5568
rect 10140 5584 10192 5636
rect 20444 5627 20496 5636
rect 7104 5516 7156 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 20444 5593 20453 5627
rect 20453 5593 20487 5627
rect 20487 5593 20496 5627
rect 20444 5584 20496 5593
rect 20260 5516 20312 5568
rect 21180 5559 21232 5568
rect 21180 5525 21189 5559
rect 21189 5525 21223 5559
rect 21223 5525 21232 5559
rect 21180 5516 21232 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2872 5312 2924 5364
rect 4068 5312 4120 5364
rect 2136 5176 2188 5228
rect 2136 4972 2188 5024
rect 2780 5040 2832 5092
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 5724 5244 5776 5296
rect 6736 5312 6788 5364
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 15568 5312 15620 5364
rect 17960 5312 18012 5364
rect 19708 5312 19760 5364
rect 8208 5244 8260 5296
rect 19984 5244 20036 5296
rect 3240 5040 3292 5092
rect 3056 4972 3108 5024
rect 4252 4972 4304 5024
rect 6552 5176 6604 5228
rect 19524 5176 19576 5228
rect 20536 5176 20588 5228
rect 5356 5108 5408 5160
rect 6368 5108 6420 5160
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6644 5151 6696 5160
rect 6460 5108 6512 5117
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 6092 4972 6144 5024
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 3332 4768 3384 4820
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 5448 4768 5500 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 7656 4768 7708 4820
rect 5356 4700 5408 4752
rect 8668 4700 8720 4752
rect 5540 4632 5592 4684
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 6092 4632 6144 4684
rect 6552 4632 6604 4684
rect 12164 4632 12216 4684
rect 6644 4564 6696 4616
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 18696 4496 18748 4548
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 5816 4428 5868 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 3240 4224 3292 4276
rect 5816 4267 5868 4276
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 2780 3952 2832 4004
rect 4620 4088 4672 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 6000 4224 6052 4276
rect 6644 4224 6696 4276
rect 5540 4156 5592 4208
rect 5816 4020 5868 4072
rect 6828 4156 6880 4208
rect 5172 3995 5224 4004
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 5632 3952 5684 4004
rect 3148 3884 3200 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 2964 3680 3016 3732
rect 4804 3680 4856 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 2780 3612 2832 3664
rect 5356 3612 5408 3664
rect 2412 3476 2464 3528
rect 3332 3408 3384 3460
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4620 3476 4672 3528
rect 5540 3544 5592 3596
rect 6552 3680 6604 3732
rect 4160 3340 4212 3392
rect 5080 3340 5132 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 2872 3136 2924 3188
rect 3056 3068 3108 3120
rect 5540 3136 5592 3188
rect 5264 3111 5316 3120
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 3884 2932 3936 2984
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 7564 3068 7616 3120
rect 12256 3043 12308 3052
rect 2228 2864 2280 2916
rect 4988 2864 5040 2916
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 11244 2796 11296 2848
rect 16028 2796 16080 2848
rect 20628 2796 20680 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 4068 2592 4120 2644
rect 6000 2592 6052 2644
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
<< metal2 >>
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2516 22222 2728 22250
rect 1688 20874 1716 22200
rect 1950 20904 2006 20913
rect 1676 20868 1728 20874
rect 1950 20839 2006 20848
rect 1676 20810 1728 20816
rect 1582 20088 1638 20097
rect 1964 20058 1992 20839
rect 2056 20534 2084 22200
rect 2424 22114 2452 22200
rect 2516 22114 2544 22222
rect 2424 22086 2544 22114
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 1582 20023 1638 20032
rect 1952 20052 2004 20058
rect 1398 15600 1454 15609
rect 1398 15535 1454 15544
rect 1412 8634 1440 15535
rect 1596 14074 1624 20023
rect 1952 19994 2004 20000
rect 2700 19938 2728 22222
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5092 22222 5304 22250
rect 2792 21434 2820 22200
rect 2792 21406 2912 21434
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 2792 20058 2820 21247
rect 2884 20602 2912 21406
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2872 20596 2924 20602
rect 2872 20538 2924 20544
rect 2870 20496 2926 20505
rect 2870 20431 2926 20440
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2778 19952 2834 19961
rect 2700 19910 2778 19938
rect 2778 19887 2834 19896
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2778 19680 2834 19689
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 18086 2452 18226
rect 2700 18193 2728 19654
rect 2778 19615 2834 19624
rect 2792 18426 2820 19615
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2686 18184 2742 18193
rect 2504 18148 2556 18154
rect 2686 18119 2742 18128
rect 2504 18090 2556 18096
rect 2412 18080 2464 18086
rect 1950 18048 2006 18057
rect 1950 17983 2006 17992
rect 2410 18048 2412 18057
rect 2464 18048 2466 18057
rect 2410 17983 2466 17992
rect 1964 17338 1992 17983
rect 2516 17678 2544 18090
rect 2884 17882 2912 20431
rect 2976 20058 3004 20878
rect 3160 20369 3188 22200
rect 3528 20505 3556 22200
rect 3896 21010 3924 22200
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 4264 20618 4292 22200
rect 4434 20904 4490 20913
rect 4434 20839 4490 20848
rect 4264 20590 4384 20618
rect 4448 20602 4476 20839
rect 3514 20496 3570 20505
rect 3514 20431 3570 20440
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20392 4212 20398
rect 3146 20360 3202 20369
rect 4160 20334 4212 20340
rect 3146 20295 3202 20304
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19514 4016 19654
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2596 17808 2648 17814
rect 2596 17750 2648 17756
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2332 17241 2360 17274
rect 2318 17232 2374 17241
rect 2228 17196 2280 17202
rect 2318 17167 2374 17176
rect 2228 17138 2280 17144
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1688 9518 1716 16594
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1964 15502 1992 15846
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11762 1808 12038
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1872 9178 1900 15127
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1964 11830 1992 13874
rect 2056 12850 2084 16050
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15026 2176 15370
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2240 14929 2268 17138
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16250 2360 16390
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2226 14920 2282 14929
rect 2226 14855 2282 14864
rect 2318 14376 2374 14385
rect 2318 14311 2374 14320
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 2226 9616 2282 9625
rect 2044 9580 2096 9586
rect 2226 9551 2282 9560
rect 2044 9522 2096 9528
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 2056 8090 2084 9522
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 6882 2084 7686
rect 2148 7002 2176 7822
rect 2240 7546 2268 9551
rect 2332 9178 2360 14311
rect 2424 9450 2452 16050
rect 2516 13025 2544 17614
rect 2608 17542 2636 17750
rect 2778 17640 2834 17649
rect 2976 17626 3004 19207
rect 2778 17575 2834 17584
rect 2884 17598 3004 17626
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2792 17338 2820 17575
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2778 16824 2834 16833
rect 2778 16759 2834 16768
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2502 13016 2558 13025
rect 2608 12986 2636 16526
rect 2792 14074 2820 16759
rect 2884 16454 2912 17598
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 16522 3004 17478
rect 3068 16658 3096 19450
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3146 18864 3202 18873
rect 3146 18799 3202 18808
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 3160 16114 3188 18799
rect 3988 18698 4016 19314
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3238 18456 3294 18465
rect 3238 18391 3294 18400
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3146 16008 3202 16017
rect 3146 15943 3202 15952
rect 2870 14784 2926 14793
rect 2870 14719 2926 14728
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 13954 2912 14719
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2792 13926 2912 13954
rect 2976 13938 3004 14214
rect 2964 13932 3016 13938
rect 2792 13546 2820 13926
rect 2964 13874 3016 13880
rect 2962 13832 3018 13841
rect 2962 13767 3018 13776
rect 2792 13518 2912 13546
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2502 12951 2558 12960
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2056 6854 2176 6882
rect 2148 5234 2176 6854
rect 2516 5846 2544 11086
rect 2700 10266 2728 11698
rect 2792 11558 2820 13398
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2884 11354 2912 13518
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2870 10704 2926 10713
rect 2870 10639 2926 10648
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2608 9674 2636 9862
rect 2608 9646 2728 9674
rect 2700 9586 2728 9646
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 7954 2636 8910
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2700 7886 2728 9522
rect 2792 9518 2820 10406
rect 2884 10266 2912 10639
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2976 9697 3004 13767
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 11898 3096 13670
rect 3160 13462 3188 15943
rect 3252 15162 3280 18391
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 4080 17746 4108 19246
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3344 17338 3372 17478
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3344 17202 3372 17274
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3882 16416 3938 16425
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3344 14482 3372 16390
rect 3882 16351 3938 16360
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3054 11792 3110 11801
rect 3054 11727 3110 11736
rect 3068 10713 3096 11727
rect 3160 11286 3188 13262
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3054 10704 3110 10713
rect 3054 10639 3110 10648
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3068 9722 3096 9862
rect 3056 9716 3108 9722
rect 2962 9688 3018 9697
rect 3056 9658 3108 9664
rect 2962 9623 3018 9632
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2792 6186 2820 9318
rect 3068 6866 3096 9454
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6458 3004 6598
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2148 5030 2176 5170
rect 2136 5024 2188 5030
rect 2240 5001 2268 5510
rect 2792 5098 2820 5714
rect 2884 5370 2912 6190
rect 2976 5914 3004 6258
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 3056 5024 3108 5030
rect 2136 4966 2188 4972
rect 2226 4992 2282 5001
rect 2148 4185 2176 4966
rect 3056 4966 3108 4972
rect 2226 4927 2282 4936
rect 2134 4176 2190 4185
rect 2134 4111 2190 4120
rect 2964 4140 3016 4146
rect 2148 3738 2176 4111
rect 2964 4082 3016 4088
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2318 3768 2374 3777
rect 2136 3732 2188 3738
rect 2188 3692 2268 3720
rect 2318 3703 2320 3712
rect 2136 3674 2188 3680
rect 2240 3618 2268 3692
rect 2372 3703 2374 3712
rect 2320 3674 2372 3680
rect 2792 3670 2820 3946
rect 2780 3664 2832 3670
rect 2240 3590 2452 3618
rect 2780 3606 2832 3612
rect 2424 3534 2452 3590
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2884 3194 2912 4014
rect 2976 3738 3004 4082
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3068 3369 3096 4966
rect 3160 3942 3188 9862
rect 3252 8634 3280 14214
rect 3436 14074 3464 15846
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3792 15088 3844 15094
rect 3790 15056 3792 15065
rect 3844 15056 3846 15065
rect 3790 14991 3846 15000
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3330 13560 3386 13569
rect 3549 13563 3857 13572
rect 3330 13495 3386 13504
rect 3344 9178 3372 13495
rect 3896 13326 3924 16351
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3988 13938 4016 15302
rect 4080 14958 4108 16594
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14074 4108 14894
rect 4172 14618 4200 20334
rect 4264 20058 4292 20402
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4250 19816 4306 19825
rect 4250 19751 4252 19760
rect 4304 19751 4306 19760
rect 4252 19722 4304 19728
rect 4252 18624 4304 18630
rect 4356 18612 4384 20590
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4436 20324 4488 20330
rect 4436 20266 4488 20272
rect 4448 19854 4476 20266
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4448 19514 4476 19790
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4448 18970 4476 19450
rect 4632 19174 4660 22200
rect 5000 20466 5028 22200
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4436 18964 4488 18970
rect 4436 18906 4488 18912
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4304 18584 4384 18612
rect 4252 18566 4304 18572
rect 4264 18290 4292 18566
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4342 18184 4398 18193
rect 4342 18119 4398 18128
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4264 16522 4292 17138
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4264 15978 4292 16118
rect 4356 16096 4384 18119
rect 4448 17746 4476 18906
rect 5000 18698 5028 18906
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4724 17678 4752 18022
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4988 17604 5040 17610
rect 4988 17546 5040 17552
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4448 16454 4476 16526
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4356 16068 4476 16096
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4356 15434 4384 15846
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4342 15056 4398 15065
rect 4252 15020 4304 15026
rect 4342 14991 4398 15000
rect 4252 14962 4304 14968
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4264 14482 4292 14962
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4356 14278 4384 14991
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 11529 3464 12378
rect 3422 11520 3478 11529
rect 3422 11455 3478 11464
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3804 11121 3832 11290
rect 3790 11112 3846 11121
rect 3790 11047 3846 11056
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 10248 3464 10610
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3436 10220 3556 10248
rect 3528 9926 3556 10220
rect 3516 9920 3568 9926
rect 3896 9897 3924 10746
rect 3988 10130 4016 13874
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3976 9920 4028 9926
rect 3516 9862 3568 9868
rect 3882 9888 3938 9897
rect 3528 9382 3556 9862
rect 3976 9862 4028 9868
rect 3882 9823 3938 9832
rect 3700 9648 3752 9654
rect 3698 9616 3700 9625
rect 3752 9616 3754 9625
rect 3698 9551 3754 9560
rect 3988 9489 4016 9862
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3252 7041 3280 7958
rect 3344 7478 3372 8842
rect 3528 8566 3556 8842
rect 3988 8673 4016 9046
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 4080 8498 4108 14010
rect 4448 12889 4476 16068
rect 4540 15706 4568 16526
rect 4816 15978 4844 16934
rect 5000 16522 5028 17546
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4540 15094 4568 15642
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4434 12880 4490 12889
rect 4434 12815 4490 12824
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 10062 4200 12582
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11558 4292 12106
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4356 11150 4384 11630
rect 4448 11257 4476 12815
rect 4526 12336 4582 12345
rect 4526 12271 4582 12280
rect 4434 11248 4490 11257
rect 4434 11183 4490 11192
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4264 9722 4292 11018
rect 4540 10146 4568 12271
rect 4448 10118 4568 10146
rect 4448 9722 4476 10118
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3988 7857 4016 8230
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 4622 3280 5034
rect 3344 4826 3372 7278
rect 3436 6866 3464 7346
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6458 3648 6598
rect 3896 6458 3924 7686
rect 4080 7449 4108 8026
rect 4172 7954 4200 9386
rect 4264 9178 4292 9658
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4448 9466 4476 9522
rect 4356 9438 4476 9466
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4356 9081 4384 9438
rect 4342 9072 4398 9081
rect 4342 9007 4398 9016
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8566 4476 8774
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4264 7546 4292 8502
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7954 4384 8298
rect 4540 7954 4568 9998
rect 4632 9518 4660 15846
rect 4816 15042 4844 15914
rect 5000 15910 5028 16458
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4724 15014 4844 15042
rect 4724 12434 4752 15014
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 13682 4844 14826
rect 4816 13654 4936 13682
rect 4724 12406 4844 12434
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4724 9518 4752 9658
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8974 4752 9318
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8424 4672 8430
rect 4618 8392 4620 8401
rect 4672 8392 4674 8401
rect 4618 8327 4674 8336
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4066 7440 4122 7449
rect 4066 7375 4122 7384
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4080 6633 4108 6734
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3974 6216 4030 6225
rect 4264 6186 4292 7346
rect 3974 6151 4030 6160
rect 4252 6180 4304 6186
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3988 5574 4016 6151
rect 4252 6122 4304 6128
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4080 5817 4108 5850
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3804 5234 3832 5510
rect 4066 5400 4122 5409
rect 4066 5335 4068 5344
rect 4120 5335 4122 5344
rect 4068 5306 4120 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3240 4616 3292 4622
rect 3238 4584 3240 4593
rect 3292 4584 3294 4593
rect 3238 4519 3294 4528
rect 3252 4282 3280 4519
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3344 3466 3372 4762
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 4078 3924 4422
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3054 3360 3110 3369
rect 3054 3295 3110 3304
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3068 3126 3096 3295
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3896 2990 3924 4014
rect 4264 3602 4292 4966
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4356 3534 4384 4422
rect 4344 3528 4396 3534
rect 4448 3516 4476 7686
rect 4540 6254 4568 7890
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4724 6866 4752 7346
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4540 5778 4568 6190
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4816 4298 4844 12406
rect 4908 6458 4936 13654
rect 5092 13530 5120 22222
rect 5276 22114 5304 22222
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8666 22200 8722 23000
rect 8772 22222 8984 22250
rect 5368 22114 5396 22200
rect 5276 22086 5396 22114
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5184 20398 5212 21014
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5538 20088 5594 20097
rect 5538 20023 5540 20032
rect 5592 20023 5594 20032
rect 5632 20052 5684 20058
rect 5540 19994 5592 20000
rect 5632 19994 5684 20000
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5552 19378 5580 19654
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5552 18873 5580 19314
rect 5538 18864 5594 18873
rect 5538 18799 5594 18808
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5552 18358 5580 18566
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5644 17202 5672 19994
rect 5736 18057 5764 22200
rect 6104 20890 6132 22200
rect 5816 20868 5868 20874
rect 5816 20810 5868 20816
rect 5920 20862 6132 20890
rect 5722 18048 5778 18057
rect 5722 17983 5778 17992
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5828 17082 5856 20810
rect 5920 17377 5948 20862
rect 6472 20856 6500 22200
rect 6840 20874 6868 22200
rect 6828 20868 6880 20874
rect 6472 20828 6592 20856
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6184 20596 6236 20602
rect 6564 20584 6592 20828
rect 6828 20810 6880 20816
rect 6184 20538 6236 20544
rect 6472 20556 6592 20584
rect 6734 20632 6790 20641
rect 7208 20602 7236 22200
rect 7380 21072 7432 21078
rect 7380 21014 7432 21020
rect 7392 20602 7420 21014
rect 7470 20904 7526 20913
rect 7470 20839 7526 20848
rect 6734 20567 6790 20576
rect 7196 20596 7248 20602
rect 6196 20505 6224 20538
rect 6182 20496 6238 20505
rect 6182 20431 6238 20440
rect 6472 19700 6500 20556
rect 6748 20534 6776 20567
rect 7196 20538 7248 20544
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 7102 20496 7158 20505
rect 6552 20256 6604 20262
rect 6920 20256 6972 20262
rect 6552 20198 6604 20204
rect 6918 20224 6920 20233
rect 6972 20224 6974 20233
rect 6472 19672 6531 19700
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6184 19508 6236 19514
rect 6503 19496 6531 19672
rect 6184 19450 6236 19456
rect 6472 19468 6531 19496
rect 6196 19417 6224 19450
rect 6182 19408 6238 19417
rect 6182 19343 6238 19352
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18766 6408 19110
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6368 18760 6420 18766
rect 6472 18737 6500 19468
rect 6564 18970 6592 20198
rect 6918 20159 6974 20168
rect 6828 19984 6880 19990
rect 6828 19926 6880 19932
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6368 18702 6420 18708
rect 6458 18728 6514 18737
rect 6012 18426 6040 18702
rect 6458 18663 6514 18672
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6196 18086 6224 18362
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6380 17524 6408 17818
rect 6564 17785 6592 18566
rect 6656 18290 6684 19654
rect 6748 19514 6776 19654
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6748 19281 6776 19450
rect 6734 19272 6790 19281
rect 6734 19207 6790 19216
rect 6734 18728 6790 18737
rect 6734 18663 6790 18672
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6656 17882 6684 18226
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6550 17776 6606 17785
rect 6748 17762 6776 18663
rect 6840 18426 6868 19926
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6932 19446 6960 19790
rect 7024 19514 7052 20470
rect 7102 20431 7158 20440
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6932 19174 6960 19382
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7024 18612 7052 18906
rect 7116 18766 7144 20431
rect 7208 19854 7236 20538
rect 7392 20262 7420 20538
rect 7484 20534 7512 20839
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7484 20058 7512 20266
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7392 19718 7420 19858
rect 7484 19718 7512 19994
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7472 19712 7524 19718
rect 7576 19700 7604 22200
rect 7748 20528 7800 20534
rect 7654 20496 7710 20505
rect 7748 20470 7800 20476
rect 7654 20431 7656 20440
rect 7708 20431 7710 20440
rect 7656 20402 7708 20408
rect 7656 19712 7708 19718
rect 7576 19672 7656 19700
rect 7472 19654 7524 19660
rect 7656 19654 7708 19660
rect 7392 19530 7420 19654
rect 7196 19508 7248 19514
rect 7392 19502 7512 19530
rect 7196 19450 7248 19456
rect 7208 18834 7236 19450
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7392 18902 7420 19314
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7380 18624 7432 18630
rect 7024 18584 7144 18612
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6550 17711 6606 17720
rect 6656 17734 6776 17762
rect 6380 17496 6592 17524
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 5906 17368 5962 17377
rect 6148 17371 6456 17380
rect 5906 17303 5962 17312
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 5644 17054 5856 17082
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15502 5396 15846
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5644 15434 5672 17054
rect 5920 16250 5948 17138
rect 6288 16794 6316 17138
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5724 16108 5776 16114
rect 5776 16068 5856 16096
rect 5724 16050 5776 16056
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5828 14822 5856 16068
rect 6458 15464 6514 15473
rect 6458 15399 6460 15408
rect 6512 15399 6514 15408
rect 6460 15370 6512 15376
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5460 14346 5488 14554
rect 5828 14414 5856 14758
rect 6564 14414 6592 17496
rect 6656 15065 6684 17734
rect 6734 17640 6790 17649
rect 6734 17575 6736 17584
rect 6788 17575 6790 17584
rect 6828 17604 6880 17610
rect 6736 17546 6788 17552
rect 6828 17546 6880 17552
rect 6840 16998 6868 17546
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6642 15056 6698 15065
rect 6642 14991 6698 15000
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5184 13258 5212 13670
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5000 12434 5028 12786
rect 5184 12646 5212 13194
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5000 12406 5120 12434
rect 5092 12084 5120 12406
rect 5184 12238 5212 12582
rect 5368 12434 5396 14282
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 5540 14000 5592 14006
rect 5816 14000 5868 14006
rect 5592 13948 5816 13954
rect 5540 13942 5868 13948
rect 5552 13926 5856 13942
rect 6366 13832 6422 13841
rect 6366 13767 6368 13776
rect 6420 13767 6422 13776
rect 6368 13738 6420 13744
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5276 12406 5396 12434
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5092 12056 5212 12084
rect 5078 11112 5134 11121
rect 5078 11047 5134 11056
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5000 8838 5028 9454
rect 5092 9178 5120 11047
rect 5184 9625 5212 12056
rect 5170 9616 5226 9625
rect 5170 9551 5226 9560
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5184 9042 5212 9454
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4988 8832 5040 8838
rect 5276 8786 5304 12406
rect 5644 12102 5672 13126
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5538 11928 5594 11937
rect 5736 11914 5764 12310
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5538 11863 5540 11872
rect 5592 11863 5594 11872
rect 5644 11886 5764 11914
rect 5540 11834 5592 11840
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 10062 5396 10610
rect 5460 10470 5488 11562
rect 5644 11082 5672 11886
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9722 5396 9998
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5552 9654 5580 9930
rect 5540 9648 5592 9654
rect 5354 9616 5410 9625
rect 5540 9590 5592 9596
rect 5354 9551 5410 9560
rect 5448 9580 5500 9586
rect 4988 8774 5040 8780
rect 5092 8758 5304 8786
rect 5092 8650 5120 8758
rect 5000 8622 5120 8650
rect 5172 8628 5224 8634
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4632 4270 4844 4298
rect 4632 4146 4660 4270
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4620 3528 4672 3534
rect 4448 3488 4620 3516
rect 4344 3470 4396 3476
rect 4620 3470 4672 3476
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3424 2984 3476 2990
rect 3422 2952 3424 2961
rect 3884 2984 3936 2990
rect 3476 2952 3478 2961
rect 2228 2916 2280 2922
rect 3884 2926 3936 2932
rect 3422 2887 3478 2896
rect 2228 2858 2280 2864
rect 2240 800 2268 2858
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4080 1737 4108 2586
rect 4172 2145 4200 3334
rect 4632 2854 4660 3470
rect 5000 2922 5028 8622
rect 5172 8570 5224 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 7750 5120 8434
rect 5184 8430 5212 8570
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5264 8424 5316 8430
rect 5368 8401 5396 9551
rect 5448 9522 5500 9528
rect 5460 9178 5488 9522
rect 5644 9450 5672 11018
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5736 9042 5764 10678
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5264 8366 5316 8372
rect 5354 8392 5410 8401
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 7274 5120 7686
rect 5276 7546 5304 8366
rect 5354 8327 5410 8336
rect 5354 7848 5410 7857
rect 5354 7783 5410 7792
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 7342 5304 7482
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5092 3398 5120 7210
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5184 4010 5212 6258
rect 5368 5710 5396 7783
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 6866 5580 7686
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4758 5396 5102
rect 5460 4826 5488 6598
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5552 5846 5580 6122
rect 5644 5846 5672 8774
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5736 5778 5764 8502
rect 5828 6254 5856 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5920 7954 5948 11018
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6564 10198 6592 14350
rect 6840 13462 6868 16934
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6932 16114 6960 16730
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16114 7052 16390
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6932 15706 6960 16050
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6932 15162 6960 15642
rect 7116 15502 7144 18584
rect 7380 18566 7432 18572
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7300 17746 7328 18294
rect 7392 18086 7420 18566
rect 7484 18193 7512 19502
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7576 18601 7604 18770
rect 7562 18592 7618 18601
rect 7562 18527 7618 18536
rect 7470 18184 7526 18193
rect 7470 18119 7526 18128
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 17338 7328 17682
rect 7392 17338 7420 18022
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6932 14618 6960 15098
rect 7024 14890 7052 15302
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6826 13152 6882 13161
rect 6826 13087 6882 13096
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9722 6040 9998
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9722 6592 10134
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5724 5296 5776 5302
rect 5828 5273 5856 5646
rect 5724 5238 5776 5244
rect 5814 5264 5870 5273
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5262 4040 5318 4049
rect 5172 4004 5224 4010
rect 5262 3975 5318 3984
rect 5172 3946 5224 3952
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5276 3126 5304 3975
rect 5368 3670 5396 4694
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4214 5580 4626
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5644 4010 5672 4422
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 3738 5764 5238
rect 5814 5199 5870 5208
rect 5920 4690 5948 7890
rect 6012 7857 6040 9658
rect 6550 9072 6606 9081
rect 6550 9007 6552 9016
rect 6604 9007 6606 9016
rect 6552 8978 6604 8984
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6104 8430 6132 8570
rect 6092 8424 6144 8430
rect 6460 8424 6512 8430
rect 6092 8366 6144 8372
rect 6458 8392 6460 8401
rect 6512 8392 6514 8401
rect 6458 8327 6514 8336
rect 6564 7886 6592 8774
rect 6552 7880 6604 7886
rect 5998 7848 6054 7857
rect 6552 7822 6604 7828
rect 5998 7783 6054 7792
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7274 6040 7686
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6656 6254 6684 11494
rect 6748 7750 6776 12922
rect 6840 12850 6868 13087
rect 7024 12918 7052 14826
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 7024 11744 7052 12854
rect 7116 12434 7144 15438
rect 7484 14482 7512 18119
rect 7576 18068 7604 18527
rect 7668 18426 7696 19654
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7656 18080 7708 18086
rect 7576 18040 7656 18068
rect 7656 18022 7708 18028
rect 7668 15434 7696 18022
rect 7760 17105 7788 20470
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 18086 7880 20198
rect 7944 18630 7972 22200
rect 8206 20632 8262 20641
rect 8206 20567 8262 20576
rect 8220 20534 8248 20567
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8036 20097 8064 20334
rect 8022 20088 8078 20097
rect 8022 20023 8078 20032
rect 8024 19372 8076 19378
rect 8128 19360 8156 20334
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8220 20233 8248 20266
rect 8206 20224 8262 20233
rect 8312 20210 8340 22200
rect 8680 20466 8708 22200
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8772 20244 8800 22222
rect 8956 22114 8984 22222
rect 9034 22200 9090 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12084 22222 12296 22250
rect 9048 22114 9076 22200
rect 8956 22086 9076 22114
rect 9232 20602 9352 20618
rect 9232 20596 9364 20602
rect 9232 20590 9312 20596
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8588 20216 8800 20244
rect 8312 20182 8524 20210
rect 8206 20159 8262 20168
rect 8298 20088 8354 20097
rect 8298 20023 8354 20032
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8220 19378 8248 19722
rect 8076 19332 8156 19360
rect 8208 19372 8260 19378
rect 8024 19314 8076 19320
rect 8208 19314 8260 19320
rect 8220 18766 8248 19314
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 8036 17202 8064 18226
rect 8312 17626 8340 20023
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 18698 8432 19790
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8312 17598 8432 17626
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7746 17096 7802 17105
rect 7746 17031 7802 17040
rect 7852 16454 7880 17138
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 16182 7880 16390
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 8036 15858 8064 16458
rect 8116 15904 8168 15910
rect 8036 15852 8116 15858
rect 8036 15846 8168 15852
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7668 14822 7696 15370
rect 7944 15094 7972 15846
rect 8036 15830 8156 15846
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7484 14074 7512 14418
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7116 12406 7420 12434
rect 7024 11716 7144 11744
rect 7010 11656 7066 11665
rect 7010 11591 7066 11600
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6840 9926 6868 10610
rect 6932 10470 6960 11086
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 10266 6960 10406
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9042 6868 9862
rect 6932 9586 6960 10202
rect 7024 9586 7052 11591
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7116 9466 7144 11716
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7208 11082 7236 11222
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7024 9438 7144 9466
rect 6932 9042 6960 9386
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7313 6776 7686
rect 6734 7304 6790 7313
rect 6734 7239 6790 7248
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6748 6458 6776 7142
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6012 4570 6040 6190
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6458 5264 6514 5273
rect 6564 5234 6592 5578
rect 6458 5199 6514 5208
rect 6552 5228 6604 5234
rect 6472 5166 6500 5199
rect 6552 5170 6604 5176
rect 6656 5166 6684 5714
rect 6748 5370 6776 6258
rect 6840 5778 6868 8978
rect 6932 7954 6960 8978
rect 7024 8566 7052 9438
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6932 5658 6960 7890
rect 7024 6662 7052 8502
rect 7208 6866 7236 11018
rect 7392 9178 7420 12406
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7484 11626 7512 12106
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7470 10160 7526 10169
rect 7470 10095 7526 10104
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7380 8968 7432 8974
rect 7378 8936 7380 8945
rect 7432 8936 7434 8945
rect 7378 8871 7434 8880
rect 7484 8430 7512 10095
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6840 5630 6960 5658
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4690 6132 4966
rect 6380 4826 6408 5102
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 5920 4542 6040 4570
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4282 5856 4422
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5920 4162 5948 4542
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5828 4134 5948 4162
rect 5828 4078 5856 4134
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5552 3194 5580 3538
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4632 2553 4660 2790
rect 6012 2650 6040 4218
rect 6564 3738 6592 4626
rect 6656 4622 6684 5102
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4282 6684 4558
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6840 4214 6868 5630
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5370 7144 5510
rect 7208 5370 7236 5646
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7300 5273 7328 5510
rect 7286 5264 7342 5273
rect 7286 5199 7342 5208
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6826 4040 6882 4049
rect 6826 3975 6882 3984
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 4618 2544 4674 2553
rect 4618 2479 4674 2488
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 4158 2136 4214 2145
rect 6148 2139 6456 2148
rect 4158 2071 4214 2080
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 6840 800 6868 3975
rect 7576 3126 7604 13466
rect 7668 8566 7696 14758
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 10470 7788 14418
rect 8036 12986 8064 15830
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14278 8156 14962
rect 8312 14385 8340 17478
rect 8298 14376 8354 14385
rect 8404 14346 8432 17598
rect 8496 14362 8524 20182
rect 8588 15026 8616 20216
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8772 19553 8800 19654
rect 8758 19544 8814 19553
rect 8956 19514 8984 19654
rect 8758 19479 8814 19488
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8956 18630 8984 18770
rect 8944 18624 8996 18630
rect 9036 18624 9088 18630
rect 8944 18566 8996 18572
rect 9034 18592 9036 18601
rect 9088 18592 9090 18601
rect 9034 18527 9090 18536
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 16998 8708 17138
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16794 8708 16934
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8588 14822 8616 14962
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8298 14311 8354 14320
rect 8392 14340 8444 14346
rect 8496 14334 8708 14362
rect 8392 14282 8444 14288
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8404 14226 8432 14282
rect 8404 14198 8524 14226
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11082 7880 11698
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 8634 7788 10406
rect 8404 9382 8432 13874
rect 8496 11762 8524 14198
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8588 13530 8616 13942
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8680 13190 8708 14334
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 6458 8340 7346
rect 8680 7342 8708 11834
rect 9048 11558 9076 12106
rect 9140 11898 9168 20402
rect 9232 19854 9260 20590
rect 9312 20538 9364 20544
rect 9416 20482 9444 22200
rect 9784 20618 9812 22200
rect 9600 20602 9812 20618
rect 9588 20596 9812 20602
rect 9640 20590 9812 20596
rect 10048 20596 10100 20602
rect 9588 20538 9640 20544
rect 10048 20538 10100 20544
rect 9312 20460 9364 20466
rect 9416 20454 9628 20482
rect 9312 20402 9364 20408
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 18902 9260 19790
rect 9324 18970 9352 20402
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9404 20256 9456 20262
rect 9508 20233 9536 20266
rect 9404 20198 9456 20204
rect 9494 20224 9550 20233
rect 9416 19514 9444 20198
rect 9494 20159 9550 20168
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9508 19718 9536 19858
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9220 18896 9272 18902
rect 9220 18838 9272 18844
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9232 16726 9260 17274
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 15502 9260 15846
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9324 15366 9352 18566
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9416 15178 9444 19450
rect 9324 15162 9444 15178
rect 9312 15156 9444 15162
rect 9364 15150 9444 15156
rect 9312 15098 9364 15104
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14074 9260 14894
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9324 13326 9352 15098
rect 9508 13870 9536 19654
rect 9600 19496 9628 20454
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 20233 9904 20334
rect 9862 20224 9918 20233
rect 9862 20159 9918 20168
rect 9770 19816 9826 19825
rect 9876 19802 9904 20159
rect 10060 19961 10088 20538
rect 10152 20482 10180 22200
rect 10152 20454 10272 20482
rect 10244 20058 10272 20454
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10046 19952 10102 19961
rect 10046 19887 10102 19896
rect 9826 19774 9904 19802
rect 9770 19751 9826 19760
rect 9600 19468 9720 19496
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9600 18970 9628 19314
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9692 18850 9720 19468
rect 9876 19360 9904 19774
rect 9954 19816 10010 19825
rect 9954 19751 10010 19760
rect 9968 19446 9996 19751
rect 10244 19514 10272 19994
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9600 18822 9720 18850
rect 9784 19332 9904 19360
rect 9600 16250 9628 18822
rect 9680 18624 9732 18630
rect 9784 18612 9812 19332
rect 10520 18698 10548 22200
rect 10888 20482 10916 22200
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11072 20534 11100 20946
rect 10796 20454 10916 20482
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10968 20460 11020 20466
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 9732 18584 9812 18612
rect 9680 18566 9732 18572
rect 9876 18154 9904 18634
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9968 18086 9996 18566
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10048 18080 10100 18086
rect 10244 18057 10272 18158
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10048 18022 10100 18028
rect 10230 18048 10286 18057
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17338 9812 17614
rect 9876 17338 9904 17818
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9784 17202 9812 17274
rect 9968 17241 9996 18022
rect 10060 17270 10088 18022
rect 10230 17983 10286 17992
rect 10232 17332 10284 17338
rect 10152 17292 10232 17320
rect 10048 17264 10100 17270
rect 9954 17232 10010 17241
rect 9772 17196 9824 17202
rect 10048 17206 10100 17212
rect 9954 17167 10010 17176
rect 9772 17138 9824 17144
rect 9784 16454 9812 17138
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16250 9812 16390
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9600 15745 9628 16186
rect 9784 16114 9812 16186
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9586 15736 9642 15745
rect 9586 15671 9642 15680
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8864 10577 8892 11290
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 9140 8129 9168 9318
rect 9324 8401 9352 13262
rect 9600 13258 9628 15302
rect 9692 14657 9720 15982
rect 9968 15706 9996 16050
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9968 15162 9996 15642
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9678 14648 9734 14657
rect 9968 14618 9996 15098
rect 9678 14583 9734 14592
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9968 14074 9996 14554
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9968 13530 9996 14010
rect 10060 14006 10088 14214
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11762 9536 12038
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11150 9536 11698
rect 9496 11144 9548 11150
rect 9416 11104 9496 11132
rect 9310 8392 9366 8401
rect 9310 8327 9366 8336
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9416 7410 9444 11104
rect 9496 11086 9548 11092
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 9926 9536 10474
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9600 8537 9628 13194
rect 9968 12986 9996 13466
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 12102 9996 12242
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11014 9812 11698
rect 10152 11014 10180 17292
rect 10232 17274 10284 17280
rect 10336 16182 10364 18090
rect 10690 17640 10746 17649
rect 10690 17575 10692 17584
rect 10744 17575 10746 17584
rect 10692 17546 10744 17552
rect 10796 16538 10824 20454
rect 10968 20402 11020 20408
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10888 20058 10916 20334
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 18766 10916 19654
rect 10980 19174 11008 20402
rect 11058 20360 11114 20369
rect 11058 20295 11114 20304
rect 11072 19990 11100 20295
rect 11150 20088 11206 20097
rect 11150 20023 11206 20032
rect 11164 19990 11192 20023
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11152 19984 11204 19990
rect 11152 19926 11204 19932
rect 11256 19378 11284 22200
rect 11624 20890 11652 22200
rect 11992 22114 12020 22200
rect 12084 22114 12112 22222
rect 11992 22086 12112 22114
rect 11624 20862 11836 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11532 20262 11560 20334
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 20058 11560 20198
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 11152 19168 11204 19174
rect 11704 19168 11756 19174
rect 11204 19128 11284 19156
rect 11152 19110 11204 19116
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10888 17338 10916 18702
rect 11072 17814 11100 18838
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11058 17640 11114 17649
rect 11058 17575 11114 17584
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 11072 16658 11100 17575
rect 11164 17338 11192 18634
rect 11256 18329 11284 19128
rect 11704 19110 11756 19116
rect 11716 18766 11744 19110
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11242 18320 11298 18329
rect 11242 18255 11244 18264
rect 11296 18255 11298 18264
rect 11244 18226 11296 18232
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11150 17096 11206 17105
rect 11150 17031 11206 17040
rect 11164 16726 11192 17031
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10796 16510 10916 16538
rect 10784 16448 10836 16454
rect 10704 16408 10784 16436
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 16017 10272 16050
rect 10230 16008 10286 16017
rect 10230 15943 10286 15952
rect 10244 15638 10272 15943
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10704 15434 10732 16408
rect 10784 16390 10836 16396
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10414 14648 10470 14657
rect 10414 14583 10470 14592
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 11558 10364 14282
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11286 10364 11494
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9876 10674 9904 10950
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 9654 9904 10406
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 10060 9994 10088 10231
rect 10140 10192 10192 10198
rect 10244 10146 10272 10610
rect 10192 10140 10272 10146
rect 10140 10134 10272 10140
rect 10152 10118 10272 10134
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9864 9648 9916 9654
rect 9678 9616 9734 9625
rect 9864 9590 9916 9596
rect 9678 9551 9734 9560
rect 9692 9110 9720 9551
rect 10244 9110 10272 10118
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9586 8528 9642 8537
rect 9586 8463 9642 8472
rect 10336 7954 10364 11222
rect 10428 9926 10456 14583
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10520 13938 10548 14282
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 12594 10548 13874
rect 10704 12850 10732 15370
rect 10888 14634 10916 16510
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10796 14606 10916 14634
rect 10980 14618 11008 14758
rect 10968 14612 11020 14618
rect 10796 14113 10824 14606
rect 10968 14554 11020 14560
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10888 14278 10916 14486
rect 10980 14414 11008 14554
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10782 14104 10838 14113
rect 10782 14039 10838 14048
rect 10888 12918 10916 14214
rect 10980 13938 11008 14350
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11072 13433 11100 14826
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11058 13424 11114 13433
rect 10968 13388 11020 13394
rect 11058 13359 11114 13368
rect 10968 13330 11020 13336
rect 10980 12918 11008 13330
rect 11072 12986 11100 13359
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10520 12566 10824 12594
rect 10796 12102 10824 12566
rect 10980 12442 11008 12854
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10980 12238 11008 12378
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10810 10548 10950
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10704 10674 10732 11018
rect 10796 10810 10824 12038
rect 10980 11898 11008 12174
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10980 11762 11008 11834
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 11354 11008 11698
rect 11072 11354 11100 12106
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10980 10742 11008 11290
rect 11058 11248 11114 11257
rect 11058 11183 11114 11192
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10980 10266 11008 10678
rect 11072 10470 11100 11183
rect 11164 11014 11192 14010
rect 11256 13870 11284 17478
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17202 11744 18090
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11716 15978 11744 17138
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15366 11560 15846
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 14278 11468 14418
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 11082 11284 12582
rect 11808 12434 11836 20862
rect 11980 20256 12032 20262
rect 11978 20224 11980 20233
rect 12032 20224 12034 20233
rect 11978 20159 12034 20168
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12176 19496 12204 19926
rect 11992 19468 12204 19496
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11900 18086 11928 18566
rect 11992 18465 12020 19468
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11978 18456 12034 18465
rect 11978 18391 12034 18400
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11992 17610 12020 18391
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11886 17504 11942 17513
rect 11886 17439 11942 17448
rect 11900 17270 11928 17439
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15586 11928 15846
rect 11900 15558 12020 15586
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 15337 11928 15438
rect 11886 15328 11942 15337
rect 11886 15263 11942 15272
rect 11992 13258 12020 15558
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11808 12406 11928 12434
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11808 11762 11836 12038
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11200 11560 11562
rect 11532 11172 11836 11200
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10520 9926 10548 9998
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10888 9382 10916 9998
rect 10980 9722 11008 10202
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11072 9489 11100 9862
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 11164 8634 11192 10610
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11348 10033 11376 10406
rect 11532 10305 11560 10406
rect 11518 10296 11574 10305
rect 11518 10231 11574 10240
rect 11334 10024 11390 10033
rect 11334 9959 11390 9968
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 6118 8248 6258
rect 8312 6254 8340 6394
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5302 8248 6054
rect 8208 5296 8260 5302
rect 7746 5264 7802 5273
rect 8208 5238 8260 5244
rect 7746 5199 7802 5208
rect 7760 5166 7788 5199
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 8680 4758 8708 7278
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9692 6458 9720 7686
rect 9784 7546 9812 7686
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10152 7206 10180 7278
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 10152 5642 10180 7142
rect 10704 6866 10732 7482
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10796 6866 10824 7278
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 11716 6662 11744 11018
rect 11808 9926 11836 11172
rect 11900 11121 11928 12406
rect 11978 12064 12034 12073
rect 11978 11999 12034 12008
rect 11992 11665 12020 11999
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 11886 11112 11942 11121
rect 12084 11082 12112 19314
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12176 18358 12204 18702
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16590 12204 16934
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 16182 12204 16526
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12268 15366 12296 22222
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13188 22222 13400 22250
rect 12360 19990 12388 22200
rect 12438 20496 12494 20505
rect 12438 20431 12440 20440
rect 12492 20431 12494 20440
rect 12440 20402 12492 20408
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12348 19848 12400 19854
rect 12452 19836 12480 20198
rect 12400 19808 12480 19836
rect 12532 19848 12584 19854
rect 12348 19790 12400 19796
rect 12532 19790 12584 19796
rect 12440 19712 12492 19718
rect 12438 19680 12440 19689
rect 12492 19680 12494 19689
rect 12544 19666 12572 19790
rect 12494 19638 12572 19666
rect 12438 19615 12494 19624
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12360 18426 12388 19382
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12452 18170 12480 18906
rect 12544 18834 12572 19110
rect 12636 18970 12664 19450
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12544 18290 12572 18770
rect 12728 18714 12756 22200
rect 13096 22114 13124 22200
rect 13188 22114 13216 22222
rect 13096 22086 13216 22114
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 12912 19786 12940 20470
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 18902 12848 19314
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12728 18686 12848 18714
rect 12820 18630 12848 18686
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12636 18193 12664 18362
rect 12622 18184 12678 18193
rect 12452 18142 12572 18170
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16522 12480 17002
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12544 16153 12572 18142
rect 12622 18119 12678 18128
rect 12728 17649 12756 18566
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12714 17640 12770 17649
rect 12714 17575 12770 17584
rect 12820 17202 12848 18294
rect 12912 17882 12940 19450
rect 13004 18193 13032 20470
rect 13174 20360 13230 20369
rect 13084 20324 13136 20330
rect 13174 20295 13230 20304
rect 13084 20266 13136 20272
rect 12990 18184 13046 18193
rect 12990 18119 13046 18128
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12912 16561 12940 17818
rect 13004 17377 13032 18022
rect 13096 17728 13124 20266
rect 13188 20262 13216 20295
rect 13176 20256 13228 20262
rect 13268 20256 13320 20262
rect 13176 20198 13228 20204
rect 13266 20224 13268 20233
rect 13320 20224 13322 20233
rect 13266 20159 13322 20168
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19242 13216 19654
rect 13280 19514 13308 19858
rect 13372 19530 13400 22222
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 13924 22222 14136 22250
rect 13464 20534 13492 22200
rect 13832 20874 13860 22200
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13464 19990 13492 20266
rect 13556 20262 13584 20470
rect 13924 20346 13952 22222
rect 14108 22114 14136 22222
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 16868 22222 17080 22250
rect 14200 22114 14228 22200
rect 14108 22086 14228 22114
rect 13740 20318 13952 20346
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13268 19508 13320 19514
rect 13372 19502 13492 19530
rect 13268 19450 13320 19456
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13188 18426 13216 18770
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13372 18358 13400 19314
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13360 17740 13412 17746
rect 13096 17700 13360 17728
rect 13360 17682 13412 17688
rect 13176 17604 13228 17610
rect 13228 17564 13308 17592
rect 13176 17546 13228 17552
rect 13174 17504 13230 17513
rect 13174 17439 13230 17448
rect 12990 17368 13046 17377
rect 12990 17303 13046 17312
rect 13004 17270 13032 17303
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 12990 17096 13046 17105
rect 13188 17082 13216 17439
rect 13280 17270 13308 17564
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13464 17184 13492 19502
rect 13648 18358 13676 19790
rect 13740 19514 13768 20318
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19922 13860 20198
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 14108 19786 14136 19994
rect 14384 19786 14412 20334
rect 14568 20058 14596 22200
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14660 20233 14688 20334
rect 14646 20224 14702 20233
rect 14646 20159 14702 20168
rect 14556 20052 14608 20058
rect 14752 20040 14780 20470
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14556 19994 14608 20000
rect 14660 20012 14780 20040
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13832 19174 13860 19246
rect 13820 19168 13872 19174
rect 13818 19136 13820 19145
rect 13872 19136 13874 19145
rect 13818 19071 13874 19080
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14384 18970 14412 19314
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13740 18222 13768 18634
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 17649 13584 17682
rect 13542 17640 13598 17649
rect 13542 17575 13598 17584
rect 13464 17156 13676 17184
rect 12990 17031 13046 17040
rect 13096 17054 13216 17082
rect 13450 17096 13506 17105
rect 13004 16998 13032 17031
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12898 16552 12954 16561
rect 12898 16487 12954 16496
rect 12530 16144 12586 16153
rect 12348 16108 12400 16114
rect 12530 16079 12586 16088
rect 12624 16108 12676 16114
rect 12348 16050 12400 16056
rect 12624 16050 12676 16056
rect 12360 15502 12388 16050
rect 12636 15706 12664 16050
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12346 14512 12402 14521
rect 12346 14447 12402 14456
rect 12360 14346 12388 14447
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12452 14074 12480 14554
rect 12544 14521 12572 14554
rect 12530 14512 12586 14521
rect 12530 14447 12586 14456
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13394 12204 13874
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12636 13326 12664 15506
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 14906 12940 14962
rect 12820 14878 12940 14906
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12820 14414 12848 14878
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13802 12848 14350
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12912 13870 12940 14282
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 11886 11047 11942 11056
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10674 11928 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11978 10568 12034 10577
rect 11978 10503 12034 10512
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11808 7410 11836 9862
rect 11992 7857 12020 10503
rect 11978 7848 12034 7857
rect 11978 7783 12034 7792
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 10520 6254 10548 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 12084 6458 12112 7414
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12176 6390 12204 11766
rect 12268 10033 12296 13262
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12438 13016 12494 13025
rect 12544 12986 12572 13126
rect 12438 12951 12494 12960
rect 12532 12980 12584 12986
rect 12452 11150 12480 12951
rect 12532 12922 12584 12928
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 11286 12572 12106
rect 12728 11914 12756 13398
rect 12820 12714 12848 13738
rect 12912 13734 12940 13806
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 13004 13462 13032 14894
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 13004 12730 13032 13398
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12912 12702 13032 12730
rect 12820 12306 12848 12650
rect 12912 12646 12940 12702
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12636 11886 12756 11914
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12254 10024 12310 10033
rect 12254 9959 12310 9968
rect 12360 9722 12388 10610
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12452 6458 12480 11086
rect 12544 9042 12572 11222
rect 12636 10577 12664 11886
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12728 11218 12756 11698
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12820 10674 12848 12242
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11286 12940 11630
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12898 11112 12954 11121
rect 12898 11047 12954 11056
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12622 10568 12678 10577
rect 12622 10503 12678 10512
rect 12636 9586 12664 10503
rect 12820 10266 12848 10610
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12820 10130 12848 10202
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12728 9466 12756 9862
rect 12820 9586 12848 10066
rect 12912 9926 12940 11047
rect 13004 10674 13032 11494
rect 13096 11014 13124 17054
rect 13450 17031 13506 17040
rect 13464 16697 13492 17031
rect 13450 16688 13506 16697
rect 13450 16623 13506 16632
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15162 13308 15302
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13648 14550 13676 17156
rect 13740 16726 13768 18158
rect 14016 18086 14044 18362
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14200 18136 14228 18226
rect 14200 18108 14320 18136
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13818 17912 13874 17921
rect 13945 17915 14253 17924
rect 13818 17847 13874 17856
rect 14004 17876 14056 17882
rect 13832 17649 13860 17847
rect 14004 17818 14056 17824
rect 13818 17640 13874 17649
rect 13818 17575 13874 17584
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13832 16658 13860 17478
rect 13910 17368 13966 17377
rect 14016 17338 14044 17818
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13910 17303 13966 17312
rect 14004 17332 14056 17338
rect 13924 17202 13952 17303
rect 14004 17274 14056 17280
rect 14108 17202 14136 17478
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 15638 13768 16390
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13818 15736 13874 15745
rect 13945 15739 14253 15748
rect 13818 15671 13820 15680
rect 13872 15671 13874 15680
rect 13820 15642 13872 15648
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13818 15464 13874 15473
rect 13818 15399 13820 15408
rect 13872 15399 13874 15408
rect 13820 15370 13872 15376
rect 14016 15026 14228 15042
rect 14004 15020 14228 15026
rect 14056 15014 14228 15020
rect 14004 14962 14056 14968
rect 14016 14929 14044 14962
rect 14200 14958 14228 15014
rect 14188 14952 14240 14958
rect 14002 14920 14058 14929
rect 14188 14894 14240 14900
rect 14002 14855 14058 14864
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 14278 13676 14486
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13818 13968 13874 13977
rect 13818 13903 13874 13912
rect 13542 13832 13598 13841
rect 13542 13767 13598 13776
rect 13450 13016 13506 13025
rect 13450 12951 13506 12960
rect 13464 12753 13492 12951
rect 13556 12918 13584 13767
rect 13832 13025 13860 13903
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13818 13016 13874 13025
rect 13636 12980 13688 12986
rect 13818 12951 13874 12960
rect 13636 12922 13688 12928
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13450 12744 13506 12753
rect 13450 12679 13506 12688
rect 13556 11898 13584 12854
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 13044 10220 13124 10248
rect 12992 10202 13044 10208
rect 13096 9994 13124 10220
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12636 9438 12756 9466
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12636 8922 12664 9438
rect 12544 8894 12664 8922
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10796 5846 10824 6326
rect 12176 6118 12204 6326
rect 12544 6254 12572 8894
rect 12728 8498 12756 8910
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12820 7818 12848 8774
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 13004 6458 13032 8774
rect 13188 7274 13216 11494
rect 13556 11286 13584 11834
rect 13648 11694 13676 12922
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14292 12442 14320 18108
rect 14384 17882 14412 18226
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 14482 14412 16934
rect 14476 16776 14504 17478
rect 14568 16969 14596 19858
rect 14660 18222 14688 20012
rect 14738 19952 14794 19961
rect 14844 19922 14872 20266
rect 14738 19887 14794 19896
rect 14832 19916 14884 19922
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14646 17776 14702 17785
rect 14646 17711 14648 17720
rect 14700 17711 14702 17720
rect 14648 17682 14700 17688
rect 14752 17626 14780 19887
rect 14832 19858 14884 19864
rect 14936 19514 14964 22200
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15028 18442 15056 20402
rect 15120 19990 15148 20810
rect 15108 19984 15160 19990
rect 15108 19926 15160 19932
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15304 19938 15332 22200
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15212 19514 15240 19926
rect 15304 19910 15424 19938
rect 15580 19922 15608 20538
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15198 19408 15254 19417
rect 15108 19372 15160 19378
rect 15198 19343 15254 19352
rect 15108 19314 15160 19320
rect 14936 18414 15056 18442
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14844 17882 14872 18226
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14752 17598 14872 17626
rect 14844 17542 14872 17598
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14554 16960 14610 16969
rect 14554 16895 14610 16904
rect 14476 16748 14780 16776
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14476 16250 14504 16526
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14462 14920 14518 14929
rect 14462 14855 14518 14864
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14384 12306 14412 13942
rect 14476 12374 14504 14855
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 14278 11792 14334 11801
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13832 11286 13860 11766
rect 14278 11727 14280 11736
rect 14332 11727 14334 11736
rect 14280 11698 14332 11704
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13358 11112 13414 11121
rect 13358 11047 13414 11056
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 10130 13308 10746
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13372 8974 13400 11047
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 9994 13860 10746
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 14108 9722 14136 10066
rect 14096 9716 14148 9722
rect 14148 9676 14320 9704
rect 14096 9658 14148 9664
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13464 6390 13492 9318
rect 13648 9178 13676 9318
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13740 8634 13768 9386
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13728 8424 13780 8430
rect 13832 8401 13860 8842
rect 13924 8566 13952 9114
rect 14292 9042 14320 9676
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13912 8560 13964 8566
rect 14108 8537 14136 8774
rect 13912 8502 13964 8508
rect 14094 8528 14150 8537
rect 14094 8463 14096 8472
rect 14148 8463 14150 8472
rect 14096 8434 14148 8440
rect 14108 8403 14136 8434
rect 13728 8366 13780 8372
rect 13818 8392 13874 8401
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13556 7750 13584 8230
rect 13648 8090 13676 8230
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13740 7449 13768 8366
rect 13818 8327 13874 8336
rect 13832 8090 13860 8327
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13832 7954 13860 8026
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13740 6322 13768 7375
rect 14384 7342 14412 10202
rect 14476 7954 14504 12038
rect 14568 8566 14596 16594
rect 14646 15464 14702 15473
rect 14646 15399 14702 15408
rect 14660 14958 14688 15399
rect 14752 15314 14780 16748
rect 14936 16590 14964 18414
rect 15120 18358 15148 19314
rect 15212 18834 15240 19343
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14844 15434 14872 15642
rect 14832 15428 14884 15434
rect 14832 15370 14884 15376
rect 14752 15286 14964 15314
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14660 10130 14688 14758
rect 14830 14648 14886 14657
rect 14830 14583 14886 14592
rect 14844 14482 14872 14583
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14830 13696 14886 13705
rect 14830 13631 14886 13640
rect 14738 12472 14794 12481
rect 14738 12407 14740 12416
rect 14792 12407 14794 12416
rect 14740 12378 14792 12384
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11898 14780 12038
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 10810 14872 13631
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14936 10690 14964 15286
rect 15028 11898 15056 17478
rect 15120 16454 15148 18158
rect 15212 17882 15240 18634
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15304 17270 15332 19790
rect 15396 19514 15424 19910
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15488 19258 15516 19858
rect 15672 19446 15700 22200
rect 16040 20602 16068 22200
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15764 19718 15792 19994
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15396 19230 15516 19258
rect 15396 17746 15424 19230
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18766 15516 19110
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15580 18426 15608 19314
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15764 18873 15792 19246
rect 15750 18864 15806 18873
rect 15750 18799 15752 18808
rect 15804 18799 15806 18808
rect 15752 18770 15804 18776
rect 15764 18739 15792 18770
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15382 16552 15438 16561
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15120 15162 15148 16186
rect 15212 16182 15240 16458
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15304 15706 15332 16526
rect 15382 16487 15438 16496
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15292 15088 15344 15094
rect 15106 15056 15162 15065
rect 15292 15030 15344 15036
rect 15396 15042 15424 16487
rect 15672 16114 15700 18566
rect 15752 18216 15804 18222
rect 15750 18184 15752 18193
rect 15804 18184 15806 18193
rect 15750 18119 15806 18128
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15580 15706 15608 15846
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 15434 15700 15846
rect 15476 15428 15528 15434
rect 15660 15428 15712 15434
rect 15528 15388 15608 15416
rect 15476 15370 15528 15376
rect 15106 14991 15162 15000
rect 15120 14958 15148 14991
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15120 14657 15148 14894
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15106 14648 15162 14657
rect 15106 14583 15162 14592
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15120 12322 15148 14486
rect 15212 14278 15240 14758
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 12442 15240 14214
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15120 12294 15240 12322
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15212 11642 15240 12294
rect 14844 10662 14964 10690
rect 15120 11614 15240 11642
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14752 9994 14780 10406
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14752 8922 14780 9930
rect 14844 9450 14872 10662
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9722 14964 9862
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 15120 9081 15148 11614
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15304 10266 15332 15030
rect 15396 15014 15516 15042
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15396 14618 15424 14894
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15488 12434 15516 15014
rect 15580 12918 15608 15388
rect 15660 15370 15712 15376
rect 15764 13530 15792 18119
rect 15856 16590 15884 20402
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19786 16068 20198
rect 16224 19854 16252 20878
rect 16408 20602 16436 22200
rect 16776 22114 16804 22200
rect 16868 22114 16896 22222
rect 16776 22086 16896 22114
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16684 20369 16712 20402
rect 16670 20360 16726 20369
rect 16396 20324 16448 20330
rect 16670 20295 16726 20304
rect 16396 20266 16448 20272
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 16408 19514 16436 20266
rect 16580 20256 16632 20262
rect 16578 20224 16580 20233
rect 16632 20224 16634 20233
rect 16578 20159 16634 20168
rect 16762 19952 16818 19961
rect 16762 19887 16818 19896
rect 16776 19854 16804 19887
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16960 19514 16988 19790
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16408 19310 16436 19450
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16394 18728 16450 18737
rect 16118 18456 16174 18465
rect 16118 18391 16174 18400
rect 16132 17746 16160 18391
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15948 16402 15976 16662
rect 16026 16552 16082 16561
rect 16026 16487 16082 16496
rect 15856 16374 15976 16402
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15764 13394 15792 13466
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15856 13326 15884 16374
rect 16040 16250 16068 16487
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15934 16144 15990 16153
rect 15934 16079 15990 16088
rect 16028 16108 16080 16114
rect 15948 16046 15976 16079
rect 16028 16050 16080 16056
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 13190 15884 13262
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15488 12406 15608 12434
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11898 15424 12038
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15488 11665 15516 12310
rect 15580 11694 15608 12406
rect 15672 12102 15700 12582
rect 15764 12306 15792 12718
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11688 15620 11694
rect 15474 11656 15530 11665
rect 15568 11630 15620 11636
rect 15474 11591 15530 11600
rect 15672 11506 15700 12038
rect 15580 11478 15700 11506
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 10810 15516 11154
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10742 15608 11478
rect 15856 11098 15884 12786
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15764 11070 15884 11098
rect 15672 10810 15700 11018
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15212 9722 15240 9998
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15304 9654 15332 9862
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15488 9586 15516 10066
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15106 9072 15162 9081
rect 15106 9007 15162 9016
rect 14660 8894 14780 8922
rect 15108 8900 15160 8906
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 8090 14596 8366
rect 14660 8294 14688 8894
rect 15108 8842 15160 8848
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8566 14780 8774
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14752 8022 14780 8502
rect 15120 8362 15148 8842
rect 15212 8430 15240 9522
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 15028 7206 15056 7822
rect 15580 7750 15608 10678
rect 15764 9466 15792 11070
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15672 9438 15792 9466
rect 15672 8974 15700 9438
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15764 7546 15792 9318
rect 15856 8945 15884 10950
rect 15948 10810 15976 15302
rect 16040 14550 16068 16050
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16026 14376 16082 14385
rect 16026 14311 16082 14320
rect 16040 12102 16068 14311
rect 16132 13274 16160 17478
rect 16224 17270 16252 18702
rect 16394 18663 16396 18672
rect 16448 18663 16450 18672
rect 16396 18634 16448 18640
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16316 18222 16344 18566
rect 16408 18426 16436 18634
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16394 17776 16450 17785
rect 16500 17746 16528 17818
rect 16394 17711 16450 17720
rect 16488 17740 16540 17746
rect 16408 17513 16436 17711
rect 16488 17682 16540 17688
rect 16672 17672 16724 17678
rect 16670 17640 16672 17649
rect 16724 17640 16726 17649
rect 16670 17575 16726 17584
rect 16394 17504 16450 17513
rect 16394 17439 16450 17448
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16500 16794 16528 17138
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16960 16522 16988 19314
rect 17052 18970 17080 22222
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 17144 19836 17172 22200
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17144 19808 17356 19836
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 19446 17264 19654
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17224 19304 17276 19310
rect 17222 19272 17224 19281
rect 17276 19272 17278 19281
rect 17328 19242 17356 19808
rect 17222 19207 17278 19216
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17420 18306 17448 19926
rect 17512 19718 17540 22200
rect 17590 20496 17646 20505
rect 17590 20431 17646 20440
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17132 18284 17184 18290
rect 17420 18278 17540 18306
rect 17132 18226 17184 18232
rect 17144 17882 17172 18226
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17052 17134 17080 17750
rect 17236 17218 17264 18022
rect 17144 17190 17264 17218
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 17144 16674 17172 17190
rect 17224 17128 17276 17134
rect 17222 17096 17224 17105
rect 17276 17096 17278 17105
rect 17222 17031 17278 17040
rect 17052 16646 17172 16674
rect 17222 16688 17278 16697
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16210 15328 16266 15337
rect 16210 15263 16266 15272
rect 16224 14482 16252 15263
rect 16316 15094 16344 16390
rect 16408 16250 16436 16390
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 17052 16266 17080 16646
rect 17328 16658 17356 18090
rect 17420 17338 17448 18158
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17222 16623 17278 16632
rect 17316 16652 17368 16658
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16960 16238 17080 16266
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16408 15450 16436 15642
rect 16500 15570 16528 16050
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 15450 16620 15506
rect 16408 15422 16620 15450
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16408 14958 16436 15422
rect 16868 15366 16896 15982
rect 16960 15609 16988 16238
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16946 15600 17002 15609
rect 16946 15535 17002 15544
rect 17052 15502 17080 16050
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15162 16988 15370
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16408 14006 16436 14486
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16592 13394 16620 14010
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16304 13320 16356 13326
rect 16132 13246 16252 13274
rect 16304 13262 16356 13268
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12918 16160 13126
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16224 12782 16252 13246
rect 16316 13190 16344 13262
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16118 12200 16174 12209
rect 16118 12135 16174 12144
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16132 11801 16160 12135
rect 16118 11792 16174 11801
rect 16118 11727 16174 11736
rect 16224 11370 16252 12310
rect 16132 11342 16252 11370
rect 16132 11150 16160 11342
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16040 11014 16068 11086
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16132 10033 16160 10066
rect 16118 10024 16174 10033
rect 16118 9959 16174 9968
rect 16132 9926 16160 9959
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15842 8936 15898 8945
rect 15842 8871 15898 8880
rect 15948 8498 15976 9114
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16132 7886 16160 9862
rect 16224 9586 16252 11222
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16316 8537 16344 13126
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16408 11898 16436 12174
rect 16960 12170 16988 12650
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16408 11694 16436 11834
rect 17052 11744 17080 15302
rect 17144 13530 17172 16526
rect 17236 15706 17264 16623
rect 17316 16594 17368 16600
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17328 16046 17356 16390
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17236 15502 17264 15642
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17328 15026 17356 15982
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17420 15706 17448 15914
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17406 15600 17462 15609
rect 17406 15535 17462 15544
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17236 11898 17264 14758
rect 17420 14634 17448 15535
rect 17328 14606 17448 14634
rect 17328 13530 17356 14606
rect 17406 14512 17462 14521
rect 17512 14482 17540 18278
rect 17604 17626 17632 20431
rect 17880 20058 17908 22200
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17972 19854 18000 20198
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 17960 19848 18012 19854
rect 17774 19816 17830 19825
rect 17684 19780 17736 19786
rect 17774 19751 17830 19760
rect 17880 19808 17960 19836
rect 17684 19722 17736 19728
rect 17696 19310 17724 19722
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17696 18902 17724 19246
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17788 17746 17816 19751
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17880 17626 17908 19808
rect 17960 19790 18012 19796
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17972 18834 18000 19382
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17604 17598 17724 17626
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17696 16250 17724 17598
rect 17788 17598 17908 17626
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17592 16176 17644 16182
rect 17788 16130 17816 17598
rect 18156 17134 18184 19926
rect 18248 19922 18276 22200
rect 18616 20058 18644 22200
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18248 19446 18276 19722
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 17882 18276 18702
rect 18340 18358 18368 19314
rect 18432 18834 18460 19790
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18340 17338 18368 17478
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17592 16118 17644 16124
rect 17604 14890 17632 16118
rect 17696 16102 17816 16130
rect 17696 15178 17724 16102
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17788 15366 17816 15399
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17696 15150 17816 15178
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17406 14447 17462 14456
rect 17500 14476 17552 14482
rect 17420 14074 17448 14447
rect 17500 14418 17552 14424
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17408 13320 17460 13326
rect 17460 13268 17540 13274
rect 17408 13262 17540 13268
rect 17420 13246 17540 13262
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17328 12374 17356 13126
rect 17420 12986 17448 13126
rect 17512 12986 17540 13246
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17498 12880 17554 12889
rect 17498 12815 17554 12824
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17512 12306 17540 12815
rect 17604 12782 17632 13806
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17696 12434 17724 15030
rect 17788 14634 17816 15150
rect 17880 14822 17908 16934
rect 18156 16794 18184 17070
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17972 16250 18000 16662
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18234 16144 18290 16153
rect 17960 16108 18012 16114
rect 18234 16079 18290 16088
rect 17960 16050 18012 16056
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17788 14606 17908 14634
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17788 13530 17816 13738
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 13394 17816 13466
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12986 17816 13126
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17880 12889 17908 14606
rect 17866 12880 17922 12889
rect 17776 12844 17828 12850
rect 17866 12815 17922 12824
rect 17776 12786 17828 12792
rect 17604 12406 17724 12434
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17052 11716 17448 11744
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 17052 11354 17080 11562
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17314 11248 17370 11257
rect 17314 11183 17370 11192
rect 17328 11150 17356 11183
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16488 10600 16540 10606
rect 16580 10600 16632 10606
rect 16488 10542 16540 10548
rect 16578 10568 16580 10577
rect 16632 10568 16634 10577
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16408 10130 16436 10202
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16500 10010 16528 10542
rect 16578 10503 16634 10512
rect 16868 10266 16896 10610
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16408 9982 16528 10010
rect 16408 9518 16436 9982
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 9654 16988 10202
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17144 9654 17172 10134
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17236 9518 17264 10474
rect 17420 10010 17448 11716
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 10130 17540 11494
rect 17604 10577 17632 12406
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11558 17724 12174
rect 17788 11626 17816 12786
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17880 12442 17908 12650
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17972 11914 18000 16050
rect 18248 16046 18276 16079
rect 18236 16040 18288 16046
rect 18142 16008 18198 16017
rect 18236 15982 18288 15988
rect 18142 15943 18198 15952
rect 18156 14958 18184 15943
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18248 15094 18276 15438
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 14006 18092 14350
rect 18156 14278 18184 14418
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18064 13734 18092 13942
rect 18052 13728 18104 13734
rect 18156 13705 18184 14214
rect 18052 13670 18104 13676
rect 18142 13696 18198 13705
rect 18142 13631 18198 13640
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18064 12918 18092 13398
rect 18052 12912 18104 12918
rect 18156 12889 18184 13631
rect 18052 12854 18104 12860
rect 18142 12880 18198 12889
rect 18142 12815 18198 12824
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12306 18092 12718
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17880 11886 18000 11914
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17590 10568 17646 10577
rect 17590 10503 17646 10512
rect 17604 10169 17632 10503
rect 17590 10160 17646 10169
rect 17500 10124 17552 10130
rect 17590 10095 17646 10104
rect 17500 10066 17552 10072
rect 17420 9982 17540 10010
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 16396 9512 16448 9518
rect 17224 9512 17276 9518
rect 16448 9460 16528 9466
rect 16396 9454 16528 9460
rect 17224 9454 17276 9460
rect 16408 9438 16528 9454
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 9042 16436 9318
rect 16500 9110 16528 9438
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 9178 16896 9318
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 17236 9042 17264 9454
rect 17420 9450 17448 9522
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16302 8528 16358 8537
rect 16302 8463 16358 8472
rect 16854 7984 16910 7993
rect 16854 7919 16856 7928
rect 16908 7919 16910 7928
rect 16856 7890 16908 7896
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 14476 6254 14504 6598
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 17144 6458 17172 7686
rect 17406 6760 17462 6769
rect 17512 6746 17540 9982
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17604 9382 17632 9930
rect 17696 9625 17724 11494
rect 17880 10826 17908 11886
rect 18064 11830 18092 12038
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11150 18000 11698
rect 18052 11688 18104 11694
rect 18248 11665 18276 14350
rect 18432 13274 18460 17546
rect 18616 17270 18644 19314
rect 18800 18698 18828 19790
rect 18984 19174 19012 22200
rect 19352 20602 19380 22200
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19720 20058 19748 22200
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18604 17264 18656 17270
rect 18800 17241 18828 17682
rect 18604 17206 18656 17212
rect 18786 17232 18842 17241
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18696 17196 18748 17202
rect 18786 17167 18842 17176
rect 18696 17138 18748 17144
rect 18524 13462 18552 17138
rect 18708 16969 18736 17138
rect 18972 16992 19024 16998
rect 18694 16960 18750 16969
rect 18972 16934 19024 16940
rect 18694 16895 18750 16904
rect 18708 16794 18736 16895
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18984 16726 19012 16934
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18616 14074 18644 14418
rect 18800 14414 18828 14758
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18708 13938 18736 14214
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18432 13246 18644 13274
rect 18708 13258 18736 13670
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11898 18368 12038
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18432 11665 18460 12786
rect 18052 11630 18104 11636
rect 18234 11656 18290 11665
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18064 11014 18092 11630
rect 18234 11591 18290 11600
rect 18418 11656 18474 11665
rect 18418 11591 18474 11600
rect 18248 11354 18276 11591
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18234 11248 18290 11257
rect 18234 11183 18290 11192
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17958 10840 18014 10849
rect 17880 10798 17958 10826
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17682 9616 17738 9625
rect 17682 9551 17738 9560
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17682 7984 17738 7993
rect 17682 7919 17738 7928
rect 17696 7313 17724 7919
rect 17682 7304 17738 7313
rect 17682 7239 17738 7248
rect 17462 6718 17540 6746
rect 17406 6695 17408 6704
rect 17460 6695 17462 6704
rect 17408 6666 17460 6672
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17788 6254 17816 10542
rect 17880 10146 17908 10798
rect 17958 10775 18014 10784
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10266 18000 10610
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17880 10118 18000 10146
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9382 17908 9862
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 8430 17908 9318
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17972 7993 18000 10118
rect 17958 7984 18014 7993
rect 18064 7954 18092 10406
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18156 9722 18184 10066
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18248 9489 18276 11183
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18340 10033 18368 11018
rect 18326 10024 18382 10033
rect 18326 9959 18382 9968
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9722 18460 9862
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18234 9480 18290 9489
rect 18234 9415 18290 9424
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 17958 7919 18014 7928
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18156 7834 18184 7890
rect 18064 7806 18184 7834
rect 18236 7812 18288 7818
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 7002 17908 7346
rect 17972 7002 18000 7686
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18064 6390 18092 7806
rect 18236 7754 18288 7760
rect 18248 7342 18276 7754
rect 18236 7336 18288 7342
rect 18340 7313 18368 8026
rect 18236 7278 18288 7284
rect 18326 7304 18382 7313
rect 18326 7239 18382 7248
rect 18432 7206 18460 9114
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18156 6769 18184 7142
rect 18142 6760 18198 6769
rect 18142 6695 18198 6704
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6458 18184 6598
rect 18340 6458 18368 7142
rect 18432 6866 18460 7142
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 18432 6254 18460 6802
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17776 6248 17828 6254
rect 18420 6248 18472 6254
rect 17776 6190 17828 6196
rect 17958 6216 18014 6225
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 12176 4690 12204 6054
rect 13832 5914 13860 6054
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 15580 5370 15608 6054
rect 17420 5914 17448 6190
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17788 5778 17816 6190
rect 18420 6190 18472 6196
rect 17958 6151 18014 6160
rect 17972 5846 18000 6151
rect 17960 5840 18012 5846
rect 18524 5817 18552 11086
rect 18616 9654 18644 13246
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18892 12434 18920 15302
rect 19076 15162 19104 18226
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19536 17785 19564 19654
rect 19798 18320 19854 18329
rect 19798 18255 19854 18264
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19522 17776 19578 17785
rect 19522 17711 19578 17720
rect 19720 17542 19748 18022
rect 19812 17746 19840 18255
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19168 17338 19196 17478
rect 19628 17338 19656 17478
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19812 17134 19840 17682
rect 19800 17128 19852 17134
rect 19246 17096 19302 17105
rect 19800 17070 19852 17076
rect 19246 17031 19248 17040
rect 19300 17031 19302 17040
rect 19248 17002 19300 17008
rect 19904 16980 19932 17750
rect 19812 16952 19932 16980
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 15162 19564 15302
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18972 13864 19024 13870
rect 18970 13832 18972 13841
rect 19024 13832 19026 13841
rect 18970 13767 19026 13776
rect 19076 13530 19104 14962
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19430 13968 19486 13977
rect 19628 13954 19656 16050
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 15162 19748 15302
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19430 13903 19432 13912
rect 19484 13903 19486 13912
rect 19536 13926 19656 13954
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19812 13954 19840 16952
rect 20088 15348 20116 22200
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20058 20208 20742
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20180 19854 20208 19994
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20456 19394 20484 22200
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20534 20088 20590 20097
rect 20534 20023 20590 20032
rect 20364 19366 20484 19394
rect 20364 19009 20392 19366
rect 20442 19272 20498 19281
rect 20442 19207 20498 19216
rect 20350 19000 20406 19009
rect 20350 18935 20406 18944
rect 20350 18864 20406 18873
rect 20350 18799 20406 18808
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20272 16998 20300 17138
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19904 15320 20116 15348
rect 19904 14074 19932 15320
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19432 13874 19484 13880
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19536 13394 19564 13926
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19720 13240 19748 13942
rect 19812 13926 19932 13954
rect 19798 13424 19854 13433
rect 19798 13359 19800 13368
rect 19852 13359 19854 13368
rect 19800 13330 19852 13336
rect 19628 13212 19748 13240
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12986 19472 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19628 12866 19656 13212
rect 18972 12844 19024 12850
rect 19628 12838 19748 12866
rect 18972 12786 19024 12792
rect 18800 12406 18920 12434
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11830 18736 12038
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18616 9382 18644 9415
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18708 9081 18736 11766
rect 18800 9489 18828 12406
rect 18984 12306 19012 12786
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18892 11694 18920 12106
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11218 18920 11630
rect 19076 11354 19104 12718
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19536 12442 19564 12718
rect 19524 12436 19576 12442
rect 19444 12406 19524 12434
rect 19444 12209 19472 12406
rect 19524 12378 19576 12384
rect 19524 12232 19576 12238
rect 19430 12200 19486 12209
rect 19524 12174 19576 12180
rect 19430 12135 19432 12144
rect 19484 12135 19486 12144
rect 19432 12106 19484 12112
rect 19444 12075 19472 12106
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18786 9480 18842 9489
rect 18786 9415 18842 9424
rect 18694 9072 18750 9081
rect 18604 9036 18656 9042
rect 18694 9007 18750 9016
rect 18604 8978 18656 8984
rect 18616 8566 18644 8978
rect 18892 8634 18920 9522
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 8974 19012 9318
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19076 8786 19104 11018
rect 19536 10742 19564 12174
rect 19720 11898 19748 12838
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19812 12306 19840 12786
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19628 11558 19656 11698
rect 19720 11694 19748 11834
rect 19800 11824 19852 11830
rect 19798 11792 19800 11801
rect 19852 11792 19854 11801
rect 19798 11727 19854 11736
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19536 10130 19564 10406
rect 19628 10130 19656 10610
rect 19708 10192 19760 10198
rect 19708 10134 19760 10140
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19628 9722 19656 9930
rect 19720 9926 19748 10134
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19524 9648 19576 9654
rect 19246 9616 19302 9625
rect 19302 9574 19472 9602
rect 19524 9590 19576 9596
rect 19246 9551 19302 9560
rect 19444 9518 19472 9574
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19536 9042 19564 9590
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19628 9110 19656 9454
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 18984 8758 19104 8786
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 8090 18644 8230
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18616 7698 18644 8026
rect 18788 7880 18840 7886
rect 18786 7848 18788 7857
rect 18984 7857 19012 8758
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19064 8424 19116 8430
rect 19168 8401 19196 8434
rect 19444 8430 19472 8502
rect 19432 8424 19484 8430
rect 19064 8366 19116 8372
rect 19154 8392 19210 8401
rect 18840 7848 18842 7857
rect 18970 7848 19026 7857
rect 18842 7806 18920 7834
rect 18786 7783 18842 7792
rect 18616 7670 18828 7698
rect 18800 7478 18828 7670
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18616 6458 18644 7414
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18708 7290 18736 7346
rect 18892 7290 18920 7806
rect 18970 7783 19026 7792
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18708 7262 18920 7290
rect 18694 7168 18750 7177
rect 18694 7103 18750 7112
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 17960 5782 18012 5788
rect 18510 5808 18566 5817
rect 17776 5772 17828 5778
rect 18510 5743 18566 5752
rect 17776 5714 17828 5720
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 5273 18000 5306
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 18708 4554 18736 7103
rect 18984 6798 19012 7686
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18696 4548 18748 4554
rect 18696 4490 18748 4496
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 12268 3058 12296 3431
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 11256 1442 11284 2790
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11256 1414 11468 1442
rect 11440 800 11468 1414
rect 16040 800 16068 2790
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 19076 1737 19104 8366
rect 19432 8366 19484 8372
rect 19154 8327 19210 8336
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19522 8120 19578 8129
rect 19522 8055 19524 8064
rect 19576 8055 19578 8064
rect 19524 8026 19576 8032
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19260 7206 19288 7278
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19536 6866 19564 7346
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19628 6798 19656 7686
rect 19720 7546 19748 9862
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19720 6866 19748 7142
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19812 6322 19840 11222
rect 19904 10538 19932 13926
rect 19996 13530 20024 15030
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14074 20116 14962
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20272 13954 20300 16934
rect 20364 15162 20392 18799
rect 20456 17338 20484 19207
rect 20548 18426 20576 20023
rect 20732 19854 20760 20198
rect 20720 19848 20772 19854
rect 20626 19816 20682 19825
rect 20720 19790 20772 19796
rect 20626 19751 20682 19760
rect 20640 18970 20668 19751
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20732 18902 20760 19110
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20536 18420 20588 18426
rect 20824 18408 20852 22200
rect 20994 21312 21050 21321
rect 20994 21247 21050 21256
rect 21008 19990 21036 21247
rect 21086 20904 21142 20913
rect 21086 20839 21142 20848
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20536 18362 20588 18368
rect 20640 18380 20852 18408
rect 20534 18048 20590 18057
rect 20534 17983 20590 17992
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20548 17218 20576 17983
rect 20640 17882 20668 18380
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20548 17190 20668 17218
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20548 15570 20576 17070
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20548 15094 20576 15370
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20088 13926 20300 13954
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 12345 20116 13926
rect 20364 13682 20392 14962
rect 20640 14618 20668 17190
rect 20732 16182 20760 18226
rect 21008 17626 21036 19790
rect 21100 19514 21128 20839
rect 21192 20058 21220 22200
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21362 20496 21418 20505
rect 21362 20431 21418 20440
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21180 19848 21232 19854
rect 21284 19836 21312 20198
rect 21376 20058 21404 20431
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21232 19808 21312 19836
rect 21180 19790 21232 19796
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20916 17598 21036 17626
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20824 16561 20852 17138
rect 20810 16552 20866 16561
rect 20810 16487 20866 16496
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20718 16008 20774 16017
rect 20718 15943 20774 15952
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20180 13654 20392 13682
rect 20180 12442 20208 13654
rect 20456 13394 20484 13806
rect 20548 13394 20576 14486
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 14074 20668 14214
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 12986 20300 13126
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20260 12368 20312 12374
rect 20074 12336 20130 12345
rect 20260 12310 20312 12316
rect 20074 12271 20130 12280
rect 20088 11801 20116 12271
rect 20272 11830 20300 12310
rect 20364 12102 20392 12582
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20260 11824 20312 11830
rect 20074 11792 20130 11801
rect 20260 11766 20312 11772
rect 20074 11727 20130 11736
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20180 11218 20208 11630
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19984 11008 20036 11014
rect 19982 10976 19984 10985
rect 20036 10976 20038 10985
rect 19982 10911 20038 10920
rect 20180 10742 20208 11154
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19904 10130 19932 10474
rect 19996 10266 20024 10542
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19904 9926 19932 10066
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 8566 19932 9862
rect 20088 9586 20116 10542
rect 20272 9654 20300 11562
rect 20350 10976 20406 10985
rect 20350 10911 20406 10920
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20272 9178 20300 9590
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8294 20024 8434
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19904 7018 19932 7890
rect 19996 7818 20024 8230
rect 20088 7954 20116 9114
rect 20364 9110 20392 10911
rect 20456 10198 20484 13330
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 11354 20576 13126
rect 20640 12306 20668 13738
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20640 11286 20668 12038
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20548 10198 20576 11086
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20180 8838 20208 9046
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 20088 7478 20116 7890
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 19904 7002 20024 7018
rect 19892 6996 20024 7002
rect 19944 6990 20024 6996
rect 19892 6938 19944 6944
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19536 6118 19564 6258
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19536 5234 19564 6054
rect 19904 5778 19932 6802
rect 19996 6390 20024 6990
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19996 5778 20024 6326
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19720 5370 19748 5510
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19996 5302 20024 5714
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19996 5166 20024 5238
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 20088 2961 20116 7414
rect 20180 7154 20208 8774
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20272 7274 20300 8434
rect 20364 8022 20392 8910
rect 20456 8906 20484 9998
rect 20548 9586 20576 10134
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20180 7126 20300 7154
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20074 2952 20130 2961
rect 20074 2887 20130 2896
rect 20180 2774 20208 6598
rect 20272 5574 20300 7126
rect 20364 6662 20392 7482
rect 20456 7206 20484 8842
rect 20548 8838 20576 9522
rect 20640 9042 20668 9522
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20456 5642 20484 7142
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20260 5568 20312 5574
rect 20548 5522 20576 8774
rect 20732 8634 20760 15943
rect 20916 14906 20944 17598
rect 20994 17232 21050 17241
rect 20994 17167 21050 17176
rect 20824 14878 20944 14906
rect 20824 14006 20852 14878
rect 20902 14376 20958 14385
rect 20902 14311 20958 14320
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20824 11898 20852 13194
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20824 11150 20852 11698
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20824 11014 20852 11086
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20824 9722 20852 9862
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20916 9450 20944 14311
rect 21008 11898 21036 17167
rect 21100 17066 21128 18566
rect 21192 17542 21220 19790
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21362 18320 21418 18329
rect 21362 18255 21418 18264
rect 21270 17640 21326 17649
rect 21270 17575 21326 17584
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21086 16552 21142 16561
rect 21086 16487 21142 16496
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10810 21036 10950
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20994 10704 21050 10713
rect 20994 10639 20996 10648
rect 21048 10639 21050 10648
rect 20996 10610 21048 10616
rect 21100 10266 21128 16487
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 14482 21220 14962
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21284 14074 21312 17575
rect 21376 17338 21404 18255
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21362 16824 21418 16833
rect 21362 16759 21418 16768
rect 21376 15162 21404 16759
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 22006 15600 22062 15609
rect 22062 15558 22140 15586
rect 22006 15535 22062 15544
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21454 15056 21510 15065
rect 21454 14991 21510 15000
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21362 13968 21418 13977
rect 21362 13903 21418 13912
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21178 13288 21234 13297
rect 21178 13223 21234 13232
rect 21192 12986 21220 13223
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21178 12880 21234 12889
rect 21178 12815 21234 12824
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21192 10146 21220 12815
rect 21284 12170 21312 13806
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21100 10118 21220 10146
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7274 20668 8230
rect 20824 7886 20852 8910
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20824 7478 20852 7822
rect 21100 7546 21128 10118
rect 21376 9450 21404 13903
rect 21468 12442 21496 14991
rect 21546 14784 21602 14793
rect 21546 14719 21602 14728
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21456 11008 21508 11014
rect 21454 10976 21456 10985
rect 21508 10976 21510 10985
rect 21454 10911 21510 10920
rect 21364 9444 21416 9450
rect 21364 9386 21416 9392
rect 21560 8090 21588 14719
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21638 13560 21694 13569
rect 21638 13495 21694 13504
rect 21652 8634 21680 13495
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 22112 8022 22140 15558
rect 22388 12374 22416 19110
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22376 12368 22428 12374
rect 22376 12310 22428 12316
rect 22480 10674 22508 17478
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20640 6458 20668 7210
rect 20732 7002 20760 7278
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 21100 6866 21128 7482
rect 21192 6934 21220 7822
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20260 5510 20312 5516
rect 20272 4593 20300 5510
rect 20364 5494 20576 5522
rect 20364 5030 20392 5494
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20548 5030 20576 5170
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20258 4584 20314 4593
rect 20258 4519 20314 4528
rect 20364 3777 20392 4966
rect 20548 4185 20576 4966
rect 20534 4176 20590 4185
rect 20534 4111 20590 4120
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20640 3505 20668 6394
rect 20626 3496 20682 3505
rect 20626 3431 20682 3440
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 20180 2746 20576 2774
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 20548 2553 20576 2746
rect 20534 2544 20590 2553
rect 20534 2479 20590 2488
rect 19062 1728 19118 1737
rect 19062 1663 19118 1672
rect 20640 800 20668 2790
rect 20916 2009 20944 6802
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5001 21220 5510
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21178 4992 21234 5001
rect 21178 4927 21234 4936
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 20902 2000 20958 2009
rect 20902 1935 20958 1944
rect 2226 0 2282 800
rect 6826 0 6882 800
rect 11426 0 11482 800
rect 16026 0 16082 800
rect 20626 0 20682 800
<< via2 >>
rect 1950 20848 2006 20904
rect 1582 20032 1638 20088
rect 1398 15544 1454 15600
rect 2778 21256 2834 21312
rect 2870 20440 2926 20496
rect 2778 19896 2834 19952
rect 2778 19624 2834 19680
rect 2686 18128 2742 18184
rect 1950 17992 2006 18048
rect 2410 18028 2412 18048
rect 2412 18028 2464 18048
rect 2464 18028 2466 18048
rect 2410 17992 2466 18028
rect 4434 20848 4490 20904
rect 3514 20440 3570 20496
rect 3146 20304 3202 20360
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 2962 19216 3018 19272
rect 2318 17176 2374 17232
rect 1858 15136 1914 15192
rect 2226 14864 2282 14920
rect 2318 14320 2374 14376
rect 2226 9560 2282 9616
rect 2778 17584 2834 17640
rect 2778 16768 2834 16824
rect 2502 12960 2558 13016
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3146 18808 3202 18864
rect 3238 18400 3294 18456
rect 3146 15952 3202 16008
rect 2870 14728 2926 14784
rect 2962 13776 3018 13832
rect 2870 10648 2926 10704
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3882 16360 3938 16416
rect 3054 11736 3110 11792
rect 3054 10648 3110 10704
rect 2962 9632 3018 9688
rect 2226 4936 2282 4992
rect 2134 4120 2190 4176
rect 2318 3732 2374 3768
rect 2318 3712 2320 3732
rect 2320 3712 2372 3732
rect 2372 3712 2374 3732
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3790 15036 3792 15056
rect 3792 15036 3844 15056
rect 3844 15036 3846 15056
rect 3790 15000 3846 15036
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3330 13504 3386 13560
rect 4250 19780 4306 19816
rect 4250 19760 4252 19780
rect 4252 19760 4304 19780
rect 4304 19760 4306 19780
rect 4342 18128 4398 18184
rect 4342 15000 4398 15056
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3422 11464 3478 11520
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3790 11056 3846 11112
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3882 9832 3938 9888
rect 3698 9596 3700 9616
rect 3700 9596 3752 9616
rect 3752 9596 3754 9616
rect 3698 9560 3754 9596
rect 3974 9424 4030 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3974 8608 4030 8664
rect 4434 12824 4490 12880
rect 4526 12280 4582 12336
rect 4434 11192 4490 11248
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3974 7792 4030 7848
rect 3238 6976 3294 7032
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4342 9016 4398 9072
rect 4618 8372 4620 8392
rect 4620 8372 4672 8392
rect 4672 8372 4674 8392
rect 4618 8336 4674 8372
rect 4066 7384 4122 7440
rect 4066 6568 4122 6624
rect 3974 6160 4030 6216
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4066 5752 4122 5808
rect 4066 5364 4122 5400
rect 4066 5344 4068 5364
rect 4068 5344 4120 5364
rect 4120 5344 4122 5364
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3238 4564 3240 4584
rect 3240 4564 3292 4584
rect 3292 4564 3294 4584
rect 3238 4528 3294 4564
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3054 3304 3110 3360
rect 5538 20052 5594 20088
rect 5538 20032 5540 20052
rect 5540 20032 5592 20052
rect 5592 20032 5594 20052
rect 5538 18808 5594 18864
rect 5722 17992 5778 18048
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6734 20576 6790 20632
rect 7470 20848 7526 20904
rect 6182 20440 6238 20496
rect 6918 20204 6920 20224
rect 6920 20204 6972 20224
rect 6972 20204 6974 20224
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6182 19352 6238 19408
rect 6918 20168 6974 20204
rect 6458 18672 6514 18728
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6734 19216 6790 19272
rect 6734 18672 6790 18728
rect 6550 17720 6606 17776
rect 7102 20440 7158 20496
rect 7654 20460 7710 20496
rect 7654 20440 7656 20460
rect 7656 20440 7708 20460
rect 7708 20440 7710 20460
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5906 17312 5962 17368
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6458 15428 6514 15464
rect 6458 15408 6460 15428
rect 6460 15408 6512 15428
rect 6512 15408 6514 15428
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6734 17604 6790 17640
rect 6734 17584 6736 17604
rect 6736 17584 6788 17604
rect 6788 17584 6790 17604
rect 6642 15000 6698 15056
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6366 13796 6422 13832
rect 6366 13776 6368 13796
rect 6368 13776 6420 13796
rect 6420 13776 6422 13796
rect 5078 11056 5134 11112
rect 5170 9560 5226 9616
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5538 11892 5594 11928
rect 5538 11872 5540 11892
rect 5540 11872 5592 11892
rect 5592 11872 5594 11892
rect 5354 9560 5410 9616
rect 3422 2932 3424 2952
rect 3424 2932 3476 2952
rect 3476 2932 3478 2952
rect 3422 2896 3478 2932
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 5354 8336 5410 8392
rect 5354 7792 5410 7848
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 7562 18536 7618 18592
rect 7470 18128 7526 18184
rect 6826 13096 6882 13152
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5262 3984 5318 4040
rect 5814 5208 5870 5264
rect 6550 9036 6606 9072
rect 6550 9016 6552 9036
rect 6552 9016 6604 9036
rect 6604 9016 6606 9036
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6458 8372 6460 8392
rect 6460 8372 6512 8392
rect 6512 8372 6514 8392
rect 6458 8336 6514 8372
rect 5998 7792 6054 7848
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 8206 20576 8262 20632
rect 8022 20032 8078 20088
rect 8206 20168 8262 20224
rect 8298 20032 8354 20088
rect 7746 17040 7802 17096
rect 7010 11600 7066 11656
rect 6734 7248 6790 7304
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6458 5208 6514 5264
rect 7470 10104 7526 10160
rect 7378 8916 7380 8936
rect 7380 8916 7432 8936
rect 7432 8916 7434 8936
rect 7378 8880 7434 8916
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 7286 5208 7342 5264
rect 6826 3984 6882 4040
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 4618 2488 4674 2544
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 4158 2080 4214 2136
rect 4066 1672 4122 1728
rect 8298 14320 8354 14376
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8758 19488 8814 19544
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9034 18572 9036 18592
rect 9036 18572 9088 18592
rect 9088 18572 9090 18592
rect 9034 18536 9090 18572
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9494 20168 9550 20224
rect 9862 20168 9918 20224
rect 9770 19760 9826 19816
rect 10046 19896 10102 19952
rect 9954 19760 10010 19816
rect 10230 17992 10286 18048
rect 9954 17176 10010 17232
rect 9586 15680 9642 15736
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8850 10512 8906 10568
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9678 14592 9734 14648
rect 9310 8336 9366 8392
rect 9126 8064 9182 8120
rect 10690 17604 10746 17640
rect 10690 17584 10692 17604
rect 10692 17584 10744 17604
rect 10744 17584 10746 17604
rect 11058 20304 11114 20360
rect 11150 20032 11206 20088
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11058 17584 11114 17640
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11242 18284 11298 18320
rect 11242 18264 11244 18284
rect 11244 18264 11296 18284
rect 11296 18264 11298 18284
rect 11150 17040 11206 17096
rect 10230 15952 10286 16008
rect 10414 14592 10470 14648
rect 10046 10240 10102 10296
rect 9678 9560 9734 9616
rect 9586 8472 9642 8528
rect 10782 14048 10838 14104
rect 11058 13368 11114 13424
rect 11058 11192 11114 11248
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11978 20204 11980 20224
rect 11980 20204 12032 20224
rect 12032 20204 12034 20224
rect 11978 20168 12034 20204
rect 11978 18400 12034 18456
rect 11886 17448 11942 17504
rect 11886 15272 11942 15328
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11058 9424 11114 9480
rect 11518 10240 11574 10296
rect 11334 9968 11390 10024
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 7746 5208 7802 5264
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 11978 12008 12034 12064
rect 11978 11600 12034 11656
rect 11886 11056 11942 11112
rect 12438 20460 12494 20496
rect 12438 20440 12440 20460
rect 12440 20440 12492 20460
rect 12492 20440 12494 20460
rect 12438 19660 12440 19680
rect 12440 19660 12492 19680
rect 12492 19660 12494 19680
rect 12438 19624 12494 19660
rect 12622 18128 12678 18184
rect 12714 17584 12770 17640
rect 13174 20304 13230 20360
rect 12990 18128 13046 18184
rect 13266 20204 13268 20224
rect 13268 20204 13320 20224
rect 13320 20204 13322 20224
rect 13266 20168 13322 20204
rect 13174 17448 13230 17504
rect 12990 17312 13046 17368
rect 12990 17040 13046 17096
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 14646 20168 14702 20224
rect 13818 19116 13820 19136
rect 13820 19116 13872 19136
rect 13872 19116 13874 19136
rect 13818 19080 13874 19116
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13542 17584 13598 17640
rect 12898 16496 12954 16552
rect 12530 16088 12586 16144
rect 12346 14456 12402 14512
rect 12530 14456 12586 14512
rect 11978 10512 12034 10568
rect 11978 7792 12034 7848
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 12438 12960 12494 13016
rect 12254 9968 12310 10024
rect 12898 11056 12954 11112
rect 12622 10512 12678 10568
rect 13450 17040 13506 17096
rect 13450 16632 13506 16688
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13818 17856 13874 17912
rect 13818 17584 13874 17640
rect 13910 17312 13966 17368
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13818 15700 13874 15736
rect 13818 15680 13820 15700
rect 13820 15680 13872 15700
rect 13872 15680 13874 15700
rect 13818 15428 13874 15464
rect 13818 15408 13820 15428
rect 13820 15408 13872 15428
rect 13872 15408 13874 15428
rect 14002 14864 14058 14920
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13818 13912 13874 13968
rect 13542 13776 13598 13832
rect 13450 12960 13506 13016
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13818 12960 13874 13016
rect 13450 12688 13506 12744
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14738 19896 14794 19952
rect 14646 17740 14702 17776
rect 14646 17720 14648 17740
rect 14648 17720 14700 17740
rect 14700 17720 14702 17740
rect 15198 19352 15254 19408
rect 14554 16904 14610 16960
rect 14462 14864 14518 14920
rect 14278 11756 14334 11792
rect 14278 11736 14280 11756
rect 14280 11736 14332 11756
rect 14332 11736 14334 11756
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13358 11056 13414 11112
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14094 8492 14150 8528
rect 14094 8472 14096 8492
rect 14096 8472 14148 8492
rect 14148 8472 14150 8492
rect 13818 8336 13874 8392
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13726 7384 13782 7440
rect 14646 15408 14702 15464
rect 14830 14592 14886 14648
rect 14830 13640 14886 13696
rect 14738 12436 14794 12472
rect 14738 12416 14740 12436
rect 14740 12416 14792 12436
rect 14792 12416 14794 12436
rect 15750 18828 15806 18864
rect 15750 18808 15752 18828
rect 15752 18808 15804 18828
rect 15804 18808 15806 18828
rect 15382 16496 15438 16552
rect 15106 15000 15162 15056
rect 15750 18164 15752 18184
rect 15752 18164 15804 18184
rect 15804 18164 15806 18184
rect 15750 18128 15806 18164
rect 15106 14592 15162 14648
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16670 20304 16726 20360
rect 16578 20204 16580 20224
rect 16580 20204 16632 20224
rect 16632 20204 16634 20224
rect 16578 20168 16634 20204
rect 16762 19896 16818 19952
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16118 18400 16174 18456
rect 16026 16496 16082 16552
rect 15934 16088 15990 16144
rect 15474 11600 15530 11656
rect 15106 9016 15162 9072
rect 16026 14320 16082 14376
rect 16394 18692 16450 18728
rect 16394 18672 16396 18692
rect 16396 18672 16448 18692
rect 16448 18672 16450 18692
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16394 17720 16450 17776
rect 16670 17620 16672 17640
rect 16672 17620 16724 17640
rect 16724 17620 16726 17640
rect 16670 17584 16726 17620
rect 16394 17448 16450 17504
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 17222 19252 17224 19272
rect 17224 19252 17276 19272
rect 17276 19252 17278 19272
rect 17222 19216 17278 19252
rect 17590 20440 17646 20496
rect 17222 17076 17224 17096
rect 17224 17076 17276 17096
rect 17276 17076 17278 17096
rect 17222 17040 17278 17076
rect 16210 15272 16266 15328
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 17222 16632 17278 16688
rect 16946 15544 17002 15600
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16118 12144 16174 12200
rect 16118 11736 16174 11792
rect 16118 9968 16174 10024
rect 15842 8880 15898 8936
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 17406 15544 17462 15600
rect 17406 14456 17462 14512
rect 17774 19760 17830 19816
rect 17774 15408 17830 15464
rect 17498 12824 17554 12880
rect 18234 16088 18290 16144
rect 17866 12824 17922 12880
rect 17314 11192 17370 11248
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16578 10548 16580 10568
rect 16580 10548 16632 10568
rect 16632 10548 16634 10568
rect 16578 10512 16634 10548
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 18142 15952 18198 16008
rect 18142 13640 18198 13696
rect 18142 12824 18198 12880
rect 17590 10512 17646 10568
rect 17590 10104 17646 10160
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16302 8472 16358 8528
rect 16854 7948 16910 7984
rect 16854 7928 16856 7948
rect 16856 7928 16908 7948
rect 16908 7928 16910 7948
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 17406 6724 17462 6760
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 18786 17176 18842 17232
rect 18694 16904 18750 16960
rect 18234 11600 18290 11656
rect 18418 11600 18474 11656
rect 18234 11192 18290 11248
rect 17682 9560 17738 9616
rect 17682 7928 17738 7984
rect 17682 7248 17738 7304
rect 17406 6704 17408 6724
rect 17408 6704 17460 6724
rect 17460 6704 17462 6724
rect 17958 10784 18014 10840
rect 17958 7928 18014 7984
rect 18326 9968 18382 10024
rect 18234 9424 18290 9480
rect 18326 7248 18382 7304
rect 18142 6704 18198 6760
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 17958 6160 18014 6216
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19798 18264 19854 18320
rect 19522 17720 19578 17776
rect 19246 17060 19302 17096
rect 19246 17040 19248 17060
rect 19248 17040 19300 17060
rect 19300 17040 19302 17060
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 18970 13812 18972 13832
rect 18972 13812 19024 13832
rect 19024 13812 19026 13832
rect 18970 13776 19026 13812
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19430 13932 19486 13968
rect 19430 13912 19432 13932
rect 19432 13912 19484 13932
rect 19484 13912 19486 13932
rect 20534 20032 20590 20088
rect 20442 19216 20498 19272
rect 20350 18944 20406 19000
rect 20350 18808 20406 18864
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19798 13388 19854 13424
rect 19798 13368 19800 13388
rect 19800 13368 19852 13388
rect 19852 13368 19854 13388
rect 18602 9424 18658 9480
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19430 12164 19486 12200
rect 19430 12144 19432 12164
rect 19432 12144 19484 12164
rect 19484 12144 19486 12164
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 18786 9424 18842 9480
rect 18694 9016 18750 9072
rect 19798 11772 19800 11792
rect 19800 11772 19852 11792
rect 19852 11772 19854 11792
rect 19798 11736 19854 11772
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19246 9560 19302 9616
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 18786 7828 18788 7848
rect 18788 7828 18840 7848
rect 18840 7828 18842 7848
rect 18786 7792 18842 7828
rect 18970 7792 19026 7848
rect 18694 7112 18750 7168
rect 18510 5752 18566 5808
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17958 5208 18014 5264
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 12254 3440 12310 3496
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19154 8336 19210 8392
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19522 8084 19578 8120
rect 19522 8064 19524 8084
rect 19524 8064 19576 8084
rect 19576 8064 19578 8084
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 20626 19760 20682 19816
rect 20994 21256 21050 21312
rect 21086 20848 21142 20904
rect 20534 17992 20590 18048
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21362 20440 21418 20496
rect 20810 16496 20866 16552
rect 20718 15952 20774 16008
rect 20074 12280 20130 12336
rect 20074 11736 20130 11792
rect 19982 10956 19984 10976
rect 19984 10956 20036 10976
rect 20036 10956 20038 10976
rect 19982 10920 20038 10956
rect 20350 10920 20406 10976
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 20074 2896 20130 2952
rect 20994 17176 21050 17232
rect 20902 14320 20958 14376
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21362 18264 21418 18320
rect 21270 17584 21326 17640
rect 21086 16496 21142 16552
rect 20994 10668 21050 10704
rect 20994 10648 20996 10668
rect 20996 10648 21048 10668
rect 21048 10648 21050 10668
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21362 16768 21418 16824
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 22006 15544 22062 15600
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21454 15000 21510 15056
rect 21362 13912 21418 13968
rect 21178 13232 21234 13288
rect 21178 12824 21234 12880
rect 21546 14728 21602 14784
rect 21454 10956 21456 10976
rect 21456 10956 21508 10976
rect 21508 10956 21510 10976
rect 21454 10920 21510 10956
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21638 13504 21694 13560
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 20258 4528 20314 4584
rect 20534 4120 20590 4176
rect 20350 3712 20406 3768
rect 20626 3440 20682 3496
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20534 2488 20590 2544
rect 19062 1672 19118 1728
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21178 4936 21234 4992
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 20902 1944 20958 2000
<< metal3 >>
rect 0 21314 800 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 800 21254
rect 2773 21251 2839 21254
rect 20989 21314 21055 21317
rect 22200 21314 23000 21344
rect 20989 21312 23000 21314
rect 20989 21256 20994 21312
rect 21050 21256 23000 21312
rect 20989 21254 23000 21256
rect 20989 21251 21055 21254
rect 22200 21224 23000 21254
rect 0 20906 800 20936
rect 1945 20906 2011 20909
rect 0 20904 2011 20906
rect 0 20848 1950 20904
rect 2006 20848 2011 20904
rect 0 20846 2011 20848
rect 0 20816 800 20846
rect 1945 20843 2011 20846
rect 4429 20906 4495 20909
rect 7465 20906 7531 20909
rect 4429 20904 7531 20906
rect 4429 20848 4434 20904
rect 4490 20848 7470 20904
rect 7526 20848 7531 20904
rect 4429 20846 7531 20848
rect 4429 20843 4495 20846
rect 7465 20843 7531 20846
rect 21081 20906 21147 20909
rect 22200 20906 23000 20936
rect 21081 20904 23000 20906
rect 21081 20848 21086 20904
rect 21142 20848 23000 20904
rect 21081 20846 23000 20848
rect 21081 20843 21147 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 6729 20634 6795 20637
rect 8201 20634 8267 20637
rect 6729 20632 8267 20634
rect 6729 20576 6734 20632
rect 6790 20576 8206 20632
rect 8262 20576 8267 20632
rect 6729 20574 8267 20576
rect 6729 20571 6795 20574
rect 8201 20571 8267 20574
rect 0 20498 800 20528
rect 2865 20498 2931 20501
rect 0 20496 2931 20498
rect 0 20440 2870 20496
rect 2926 20440 2931 20496
rect 0 20438 2931 20440
rect 0 20408 800 20438
rect 2865 20435 2931 20438
rect 3509 20498 3575 20501
rect 6177 20498 6243 20501
rect 7097 20498 7163 20501
rect 7649 20498 7715 20501
rect 12433 20498 12499 20501
rect 17585 20498 17651 20501
rect 3509 20496 17651 20498
rect 3509 20440 3514 20496
rect 3570 20440 6182 20496
rect 6238 20440 7102 20496
rect 7158 20440 7654 20496
rect 7710 20440 12438 20496
rect 12494 20440 17590 20496
rect 17646 20440 17651 20496
rect 3509 20438 17651 20440
rect 3509 20435 3575 20438
rect 6177 20435 6243 20438
rect 7097 20435 7163 20438
rect 7649 20435 7715 20438
rect 12433 20435 12499 20438
rect 17585 20435 17651 20438
rect 21357 20498 21423 20501
rect 22200 20498 23000 20528
rect 21357 20496 23000 20498
rect 21357 20440 21362 20496
rect 21418 20440 23000 20496
rect 21357 20438 23000 20440
rect 21357 20435 21423 20438
rect 22200 20408 23000 20438
rect 3141 20362 3207 20365
rect 11053 20362 11119 20365
rect 13169 20362 13235 20365
rect 16665 20362 16731 20365
rect 16982 20362 16988 20364
rect 3141 20360 13002 20362
rect 3141 20304 3146 20360
rect 3202 20304 11058 20360
rect 11114 20304 13002 20360
rect 3141 20302 13002 20304
rect 3141 20299 3207 20302
rect 11053 20299 11119 20302
rect 6913 20226 6979 20229
rect 8201 20226 8267 20229
rect 6913 20224 8267 20226
rect 6913 20168 6918 20224
rect 6974 20168 8206 20224
rect 8262 20168 8267 20224
rect 6913 20166 8267 20168
rect 6913 20163 6979 20166
rect 8201 20163 8267 20166
rect 9254 20164 9260 20228
rect 9324 20226 9330 20228
rect 9489 20226 9555 20229
rect 9324 20224 9555 20226
rect 9324 20168 9494 20224
rect 9550 20168 9555 20224
rect 9324 20166 9555 20168
rect 9324 20164 9330 20166
rect 9489 20163 9555 20166
rect 9857 20226 9923 20229
rect 11973 20226 12039 20229
rect 9857 20224 12039 20226
rect 9857 20168 9862 20224
rect 9918 20168 11978 20224
rect 12034 20168 12039 20224
rect 9857 20166 12039 20168
rect 12942 20226 13002 20302
rect 13169 20360 14658 20362
rect 13169 20304 13174 20360
rect 13230 20304 14658 20360
rect 13169 20302 14658 20304
rect 13169 20299 13235 20302
rect 14598 20229 14658 20302
rect 16665 20360 16988 20362
rect 16665 20304 16670 20360
rect 16726 20304 16988 20360
rect 16665 20302 16988 20304
rect 16665 20299 16731 20302
rect 16982 20300 16988 20302
rect 17052 20300 17058 20364
rect 13261 20226 13327 20229
rect 12942 20224 13327 20226
rect 12942 20168 13266 20224
rect 13322 20168 13327 20224
rect 12942 20166 13327 20168
rect 14598 20226 14707 20229
rect 16573 20226 16639 20229
rect 14598 20224 16639 20226
rect 14598 20168 14646 20224
rect 14702 20168 16578 20224
rect 16634 20168 16639 20224
rect 14598 20166 16639 20168
rect 9857 20163 9923 20166
rect 11973 20163 12039 20166
rect 13261 20163 13327 20166
rect 14641 20163 14707 20166
rect 16573 20163 16639 20166
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 5533 20090 5599 20093
rect 8017 20090 8083 20093
rect 8293 20090 8359 20093
rect 11145 20090 11211 20093
rect 5533 20088 8359 20090
rect 5533 20032 5538 20088
rect 5594 20032 8022 20088
rect 8078 20032 8298 20088
rect 8354 20032 8359 20088
rect 5533 20030 8359 20032
rect 5533 20027 5599 20030
rect 8017 20027 8083 20030
rect 8293 20027 8359 20030
rect 9446 20088 11211 20090
rect 9446 20032 11150 20088
rect 11206 20032 11211 20088
rect 9446 20030 11211 20032
rect 2773 19954 2839 19957
rect 9446 19954 9506 20030
rect 11145 20027 11211 20030
rect 20529 20090 20595 20093
rect 22200 20090 23000 20120
rect 20529 20088 23000 20090
rect 20529 20032 20534 20088
rect 20590 20032 23000 20088
rect 20529 20030 23000 20032
rect 20529 20027 20595 20030
rect 22200 20000 23000 20030
rect 2773 19952 9506 19954
rect 2773 19896 2778 19952
rect 2834 19896 9506 19952
rect 2773 19894 9506 19896
rect 10041 19954 10107 19957
rect 14733 19954 14799 19957
rect 10041 19952 14799 19954
rect 10041 19896 10046 19952
rect 10102 19896 14738 19952
rect 14794 19896 14799 19952
rect 10041 19894 14799 19896
rect 2773 19891 2839 19894
rect 10041 19891 10107 19894
rect 14733 19891 14799 19894
rect 16757 19954 16823 19957
rect 17902 19954 17908 19956
rect 16757 19952 17908 19954
rect 16757 19896 16762 19952
rect 16818 19896 17908 19952
rect 16757 19894 17908 19896
rect 16757 19891 16823 19894
rect 17902 19892 17908 19894
rect 17972 19892 17978 19956
rect 4245 19818 4311 19821
rect 9765 19818 9831 19821
rect 4245 19816 9831 19818
rect 4245 19760 4250 19816
rect 4306 19760 9770 19816
rect 9826 19760 9831 19816
rect 4245 19758 9831 19760
rect 4245 19755 4311 19758
rect 9765 19755 9831 19758
rect 9949 19818 10015 19821
rect 17769 19818 17835 19821
rect 9949 19816 17835 19818
rect 9949 19760 9954 19816
rect 10010 19760 17774 19816
rect 17830 19760 17835 19816
rect 9949 19758 17835 19760
rect 9949 19755 10015 19758
rect 17769 19755 17835 19758
rect 20621 19818 20687 19821
rect 20621 19816 22202 19818
rect 20621 19760 20626 19816
rect 20682 19760 22202 19816
rect 20621 19758 22202 19760
rect 20621 19755 20687 19758
rect 22142 19712 22202 19758
rect 0 19682 800 19712
rect 2773 19682 2839 19685
rect 12433 19682 12499 19685
rect 12566 19682 12572 19684
rect 0 19680 2839 19682
rect 0 19624 2778 19680
rect 2834 19624 2839 19680
rect 0 19622 2839 19624
rect 0 19592 800 19622
rect 2773 19619 2839 19622
rect 8526 19622 9874 19682
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 6177 19410 6243 19413
rect 6862 19410 6868 19412
rect 6177 19408 6868 19410
rect 6177 19352 6182 19408
rect 6238 19352 6868 19408
rect 6177 19350 6868 19352
rect 6177 19347 6243 19350
rect 6862 19348 6868 19350
rect 6932 19410 6938 19412
rect 8526 19410 8586 19622
rect 8753 19546 8819 19549
rect 9622 19546 9628 19548
rect 8753 19544 9628 19546
rect 8753 19488 8758 19544
rect 8814 19488 9628 19544
rect 8753 19486 9628 19488
rect 8753 19483 8819 19486
rect 9622 19484 9628 19486
rect 9692 19484 9698 19548
rect 6932 19350 8586 19410
rect 9814 19410 9874 19622
rect 12433 19680 12572 19682
rect 12433 19624 12438 19680
rect 12494 19624 12572 19680
rect 12433 19622 12572 19624
rect 12433 19619 12499 19622
rect 12566 19620 12572 19622
rect 12636 19620 12642 19684
rect 22142 19622 23000 19712
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 15193 19410 15259 19413
rect 9814 19408 15259 19410
rect 9814 19352 15198 19408
rect 15254 19352 15259 19408
rect 9814 19350 15259 19352
rect 6932 19348 6938 19350
rect 15193 19347 15259 19350
rect 0 19274 800 19304
rect 2957 19274 3023 19277
rect 0 19272 3023 19274
rect 0 19216 2962 19272
rect 3018 19216 3023 19272
rect 0 19214 3023 19216
rect 0 19184 800 19214
rect 2957 19211 3023 19214
rect 6729 19274 6795 19277
rect 17217 19274 17283 19277
rect 6729 19272 17283 19274
rect 6729 19216 6734 19272
rect 6790 19216 17222 19272
rect 17278 19216 17283 19272
rect 6729 19214 17283 19216
rect 6729 19211 6795 19214
rect 17217 19211 17283 19214
rect 20437 19274 20503 19277
rect 22200 19274 23000 19304
rect 20437 19272 23000 19274
rect 20437 19216 20442 19272
rect 20498 19216 23000 19272
rect 20437 19214 23000 19216
rect 20437 19211 20503 19214
rect 22200 19184 23000 19214
rect 12198 19076 12204 19140
rect 12268 19138 12274 19140
rect 13813 19138 13879 19141
rect 12268 19136 13879 19138
rect 12268 19080 13818 19136
rect 13874 19080 13879 19136
rect 12268 19078 13879 19080
rect 12268 19076 12274 19078
rect 13813 19075 13879 19078
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 19558 18940 19564 19004
rect 19628 19002 19634 19004
rect 20345 19002 20411 19005
rect 19628 19000 20411 19002
rect 19628 18944 20350 19000
rect 20406 18944 20411 19000
rect 19628 18942 20411 18944
rect 19628 18940 19634 18942
rect 20345 18939 20411 18942
rect 0 18866 800 18896
rect 3141 18866 3207 18869
rect 0 18864 3207 18866
rect 0 18808 3146 18864
rect 3202 18808 3207 18864
rect 0 18806 3207 18808
rect 0 18776 800 18806
rect 3141 18803 3207 18806
rect 5533 18866 5599 18869
rect 15745 18866 15811 18869
rect 5533 18864 15811 18866
rect 5533 18808 5538 18864
rect 5594 18808 15750 18864
rect 15806 18808 15811 18864
rect 5533 18806 15811 18808
rect 5533 18803 5599 18806
rect 15745 18803 15811 18806
rect 20345 18866 20411 18869
rect 22200 18866 23000 18896
rect 20345 18864 23000 18866
rect 20345 18808 20350 18864
rect 20406 18808 23000 18864
rect 20345 18806 23000 18808
rect 20345 18803 20411 18806
rect 22200 18776 23000 18806
rect 6453 18730 6519 18733
rect 6729 18730 6795 18733
rect 16389 18730 16455 18733
rect 6453 18728 6795 18730
rect 6453 18672 6458 18728
rect 6514 18672 6734 18728
rect 6790 18672 6795 18728
rect 6453 18670 6795 18672
rect 6453 18667 6519 18670
rect 6729 18667 6795 18670
rect 7238 18728 16455 18730
rect 7238 18672 16394 18728
rect 16450 18672 16455 18728
rect 7238 18670 16455 18672
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 3233 18458 3299 18461
rect 0 18456 3299 18458
rect 0 18400 3238 18456
rect 3294 18400 3299 18456
rect 0 18398 3299 18400
rect 0 18368 800 18398
rect 3233 18395 3299 18398
rect 2681 18186 2747 18189
rect 4337 18186 4403 18189
rect 7238 18186 7298 18670
rect 16389 18667 16455 18670
rect 7557 18594 7623 18597
rect 9029 18594 9095 18597
rect 7557 18592 9095 18594
rect 7557 18536 7562 18592
rect 7618 18536 9034 18592
rect 9090 18536 9095 18592
rect 7557 18534 9095 18536
rect 7557 18531 7623 18534
rect 9029 18531 9095 18534
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 11973 18458 12039 18461
rect 16113 18458 16179 18461
rect 22200 18458 23000 18488
rect 11973 18456 16179 18458
rect 11973 18400 11978 18456
rect 12034 18400 16118 18456
rect 16174 18400 16179 18456
rect 11973 18398 16179 18400
rect 11973 18395 12039 18398
rect 16113 18395 16179 18398
rect 22142 18368 23000 18458
rect 11237 18322 11303 18325
rect 19793 18322 19859 18325
rect 11237 18320 19859 18322
rect 11237 18264 11242 18320
rect 11298 18264 19798 18320
rect 19854 18264 19859 18320
rect 11237 18262 19859 18264
rect 11237 18259 11303 18262
rect 19793 18259 19859 18262
rect 21357 18322 21423 18325
rect 22142 18322 22202 18368
rect 21357 18320 22202 18322
rect 21357 18264 21362 18320
rect 21418 18264 22202 18320
rect 21357 18262 22202 18264
rect 21357 18259 21423 18262
rect 2681 18184 7298 18186
rect 2681 18128 2686 18184
rect 2742 18128 4342 18184
rect 4398 18128 7298 18184
rect 2681 18126 7298 18128
rect 7465 18186 7531 18189
rect 12617 18186 12683 18189
rect 7465 18184 12683 18186
rect 7465 18128 7470 18184
rect 7526 18128 12622 18184
rect 12678 18128 12683 18184
rect 7465 18126 12683 18128
rect 2681 18123 2747 18126
rect 4337 18123 4403 18126
rect 7465 18123 7531 18126
rect 12617 18123 12683 18126
rect 12750 18124 12756 18188
rect 12820 18186 12826 18188
rect 12985 18186 13051 18189
rect 15745 18186 15811 18189
rect 12820 18184 13051 18186
rect 12820 18128 12990 18184
rect 13046 18128 13051 18184
rect 12820 18126 13051 18128
rect 12820 18124 12826 18126
rect 12985 18123 13051 18126
rect 13816 18184 15811 18186
rect 13816 18128 15750 18184
rect 15806 18128 15811 18184
rect 13816 18126 15811 18128
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 2405 18050 2471 18053
rect 3366 18050 3372 18052
rect 2405 18048 3372 18050
rect 2405 17992 2410 18048
rect 2466 17992 3372 18048
rect 2405 17990 3372 17992
rect 2405 17987 2471 17990
rect 3366 17988 3372 17990
rect 3436 17988 3442 18052
rect 5717 18050 5783 18053
rect 5942 18050 5948 18052
rect 5717 18048 5948 18050
rect 5717 17992 5722 18048
rect 5778 17992 5948 18048
rect 5717 17990 5948 17992
rect 5717 17987 5783 17990
rect 5942 17988 5948 17990
rect 6012 17988 6018 18052
rect 10225 18050 10291 18053
rect 13816 18050 13876 18126
rect 15745 18123 15811 18126
rect 10225 18048 13876 18050
rect 10225 17992 10230 18048
rect 10286 17992 13876 18048
rect 10225 17990 13876 17992
rect 20529 18050 20595 18053
rect 22200 18050 23000 18080
rect 20529 18048 23000 18050
rect 20529 17992 20534 18048
rect 20590 17992 23000 18048
rect 20529 17990 23000 17992
rect 10225 17987 10291 17990
rect 20529 17987 20595 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 9622 17852 9628 17916
rect 9692 17914 9698 17916
rect 13813 17914 13879 17917
rect 9692 17912 13879 17914
rect 9692 17856 13818 17912
rect 13874 17856 13879 17912
rect 9692 17854 13879 17856
rect 9692 17852 9698 17854
rect 13813 17851 13879 17854
rect 6545 17778 6611 17781
rect 14641 17778 14707 17781
rect 6545 17776 14707 17778
rect 6545 17720 6550 17776
rect 6606 17720 14646 17776
rect 14702 17720 14707 17776
rect 6545 17718 14707 17720
rect 6545 17715 6611 17718
rect 14641 17715 14707 17718
rect 16389 17778 16455 17781
rect 19517 17778 19583 17781
rect 16389 17776 19583 17778
rect 16389 17720 16394 17776
rect 16450 17720 19522 17776
rect 19578 17720 19583 17776
rect 16389 17718 19583 17720
rect 16389 17715 16455 17718
rect 19517 17715 19583 17718
rect 0 17642 800 17672
rect 2773 17642 2839 17645
rect 0 17640 2839 17642
rect 0 17584 2778 17640
rect 2834 17584 2839 17640
rect 0 17582 2839 17584
rect 0 17552 800 17582
rect 2773 17579 2839 17582
rect 6729 17642 6795 17645
rect 10685 17642 10751 17645
rect 6729 17640 10751 17642
rect 6729 17584 6734 17640
rect 6790 17584 10690 17640
rect 10746 17584 10751 17640
rect 6729 17582 10751 17584
rect 6729 17579 6795 17582
rect 10685 17579 10751 17582
rect 11053 17642 11119 17645
rect 12709 17642 12775 17645
rect 13537 17642 13603 17645
rect 11053 17640 12775 17642
rect 11053 17584 11058 17640
rect 11114 17584 12714 17640
rect 12770 17584 12775 17640
rect 11053 17582 12775 17584
rect 11053 17579 11119 17582
rect 12709 17579 12775 17582
rect 12896 17640 13603 17642
rect 12896 17584 13542 17640
rect 13598 17584 13603 17640
rect 12896 17582 13603 17584
rect 11881 17506 11947 17509
rect 12896 17506 12956 17582
rect 13537 17579 13603 17582
rect 13813 17642 13879 17645
rect 16665 17642 16731 17645
rect 13813 17640 16731 17642
rect 13813 17584 13818 17640
rect 13874 17584 16670 17640
rect 16726 17584 16731 17640
rect 13813 17582 16731 17584
rect 13813 17579 13879 17582
rect 16665 17579 16731 17582
rect 21265 17642 21331 17645
rect 22200 17642 23000 17672
rect 21265 17640 23000 17642
rect 21265 17584 21270 17640
rect 21326 17584 23000 17640
rect 21265 17582 23000 17584
rect 21265 17579 21331 17582
rect 22200 17552 23000 17582
rect 11881 17504 12956 17506
rect 11881 17448 11886 17504
rect 11942 17448 12956 17504
rect 11881 17446 12956 17448
rect 13169 17506 13235 17509
rect 16389 17506 16455 17509
rect 13169 17504 16455 17506
rect 13169 17448 13174 17504
rect 13230 17448 16394 17504
rect 16450 17448 16455 17504
rect 13169 17446 16455 17448
rect 11881 17443 11947 17446
rect 13169 17443 13235 17446
rect 16389 17443 16455 17446
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 5390 17308 5396 17372
rect 5460 17370 5466 17372
rect 5901 17370 5967 17373
rect 5460 17368 5967 17370
rect 5460 17312 5906 17368
rect 5962 17312 5967 17368
rect 5460 17310 5967 17312
rect 5460 17308 5466 17310
rect 5901 17307 5967 17310
rect 12985 17370 13051 17373
rect 13905 17370 13971 17373
rect 12985 17368 13971 17370
rect 12985 17312 12990 17368
rect 13046 17312 13910 17368
rect 13966 17312 13971 17368
rect 12985 17310 13971 17312
rect 12985 17307 13051 17310
rect 13905 17307 13971 17310
rect 0 17234 800 17264
rect 2313 17234 2379 17237
rect 0 17232 2379 17234
rect 0 17176 2318 17232
rect 2374 17176 2379 17232
rect 0 17174 2379 17176
rect 0 17144 800 17174
rect 2313 17171 2379 17174
rect 9949 17234 10015 17237
rect 18781 17234 18847 17237
rect 9949 17232 18847 17234
rect 9949 17176 9954 17232
rect 10010 17176 18786 17232
rect 18842 17176 18847 17232
rect 9949 17174 18847 17176
rect 9949 17171 10015 17174
rect 18781 17171 18847 17174
rect 20989 17234 21055 17237
rect 22200 17234 23000 17264
rect 20989 17232 23000 17234
rect 20989 17176 20994 17232
rect 21050 17176 23000 17232
rect 20989 17174 23000 17176
rect 20989 17171 21055 17174
rect 22200 17144 23000 17174
rect 7741 17098 7807 17101
rect 11145 17098 11211 17101
rect 12985 17098 13051 17101
rect 7741 17096 9322 17098
rect 7741 17040 7746 17096
rect 7802 17040 9322 17096
rect 7741 17038 9322 17040
rect 7741 17035 7807 17038
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 2773 16826 2839 16829
rect 0 16824 2839 16826
rect 0 16768 2778 16824
rect 2834 16768 2839 16824
rect 0 16766 2839 16768
rect 9262 16826 9322 17038
rect 11145 17096 13051 17098
rect 11145 17040 11150 17096
rect 11206 17040 12990 17096
rect 13046 17040 13051 17096
rect 11145 17038 13051 17040
rect 11145 17035 11211 17038
rect 12985 17035 13051 17038
rect 13445 17098 13511 17101
rect 17217 17098 17283 17101
rect 18086 17098 18092 17100
rect 13445 17096 17050 17098
rect 13445 17040 13450 17096
rect 13506 17040 17050 17096
rect 13445 17038 17050 17040
rect 13445 17035 13511 17038
rect 14549 16964 14615 16965
rect 14549 16960 14596 16964
rect 14660 16962 14666 16964
rect 16990 16962 17050 17038
rect 17217 17096 18092 17098
rect 17217 17040 17222 17096
rect 17278 17040 18092 17096
rect 17217 17038 18092 17040
rect 17217 17035 17283 17038
rect 18086 17036 18092 17038
rect 18156 17098 18162 17100
rect 19241 17098 19307 17101
rect 18156 17096 19307 17098
rect 18156 17040 19246 17096
rect 19302 17040 19307 17096
rect 18156 17038 19307 17040
rect 18156 17036 18162 17038
rect 19241 17035 19307 17038
rect 18689 16964 18755 16965
rect 18638 16962 18644 16964
rect 14549 16904 14554 16960
rect 14549 16900 14596 16904
rect 14660 16902 14706 16962
rect 16990 16902 18644 16962
rect 18708 16960 18755 16964
rect 18750 16904 18755 16960
rect 14660 16900 14666 16902
rect 18638 16900 18644 16902
rect 18708 16900 18755 16904
rect 14549 16899 14615 16900
rect 18689 16899 18755 16900
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 21357 16826 21423 16829
rect 22200 16826 23000 16856
rect 9262 16766 13738 16826
rect 0 16736 800 16766
rect 2773 16763 2839 16766
rect 3366 16628 3372 16692
rect 3436 16690 3442 16692
rect 13445 16690 13511 16693
rect 3436 16688 13511 16690
rect 3436 16632 13450 16688
rect 13506 16632 13511 16688
rect 3436 16630 13511 16632
rect 13678 16690 13738 16766
rect 21357 16824 23000 16826
rect 21357 16768 21362 16824
rect 21418 16768 23000 16824
rect 21357 16766 23000 16768
rect 21357 16763 21423 16766
rect 22200 16736 23000 16766
rect 17217 16690 17283 16693
rect 13678 16688 17283 16690
rect 13678 16632 17222 16688
rect 17278 16632 17283 16688
rect 13678 16630 17283 16632
rect 3436 16628 3442 16630
rect 13445 16627 13511 16630
rect 17217 16627 17283 16630
rect 12893 16554 12959 16557
rect 15377 16554 15443 16557
rect 12893 16552 15443 16554
rect 12893 16496 12898 16552
rect 12954 16496 15382 16552
rect 15438 16496 15443 16552
rect 12893 16494 15443 16496
rect 12893 16491 12959 16494
rect 15377 16491 15443 16494
rect 16021 16554 16087 16557
rect 18270 16554 18276 16556
rect 16021 16552 18276 16554
rect 16021 16496 16026 16552
rect 16082 16496 18276 16552
rect 16021 16494 18276 16496
rect 16021 16491 16087 16494
rect 18270 16492 18276 16494
rect 18340 16554 18346 16556
rect 20805 16554 20871 16557
rect 18340 16552 20871 16554
rect 18340 16496 20810 16552
rect 20866 16496 20871 16552
rect 18340 16494 20871 16496
rect 18340 16492 18346 16494
rect 20805 16491 20871 16494
rect 21081 16554 21147 16557
rect 21081 16552 22202 16554
rect 21081 16496 21086 16552
rect 21142 16496 22202 16552
rect 21081 16494 22202 16496
rect 21081 16491 21147 16494
rect 22142 16448 22202 16494
rect 0 16418 800 16448
rect 3877 16418 3943 16421
rect 0 16416 3943 16418
rect 0 16360 3882 16416
rect 3938 16360 3943 16416
rect 0 16358 3943 16360
rect 22142 16358 23000 16448
rect 0 16328 800 16358
rect 3877 16355 3943 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 12525 16146 12591 16149
rect 15929 16146 15995 16149
rect 18229 16146 18295 16149
rect 12525 16144 18295 16146
rect 12525 16088 12530 16144
rect 12586 16088 15934 16144
rect 15990 16088 18234 16144
rect 18290 16088 18295 16144
rect 12525 16086 18295 16088
rect 12525 16083 12591 16086
rect 15929 16083 15995 16086
rect 18229 16083 18295 16086
rect 0 16010 800 16040
rect 3141 16010 3207 16013
rect 0 16008 3207 16010
rect 0 15952 3146 16008
rect 3202 15952 3207 16008
rect 0 15950 3207 15952
rect 0 15920 800 15950
rect 3141 15947 3207 15950
rect 10225 16010 10291 16013
rect 18137 16010 18203 16013
rect 10225 16008 18203 16010
rect 10225 15952 10230 16008
rect 10286 15952 18142 16008
rect 18198 15952 18203 16008
rect 10225 15950 18203 15952
rect 10225 15947 10291 15950
rect 18137 15947 18203 15950
rect 20713 16010 20779 16013
rect 22200 16010 23000 16040
rect 20713 16008 23000 16010
rect 20713 15952 20718 16008
rect 20774 15952 23000 16008
rect 20713 15950 23000 15952
rect 20713 15947 20779 15950
rect 22200 15920 23000 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 9581 15738 9647 15741
rect 13813 15738 13879 15741
rect 9581 15736 13879 15738
rect 9581 15680 9586 15736
rect 9642 15680 13818 15736
rect 13874 15680 13879 15736
rect 9581 15678 13879 15680
rect 9581 15675 9647 15678
rect 13813 15675 13879 15678
rect 0 15602 800 15632
rect 1393 15602 1459 15605
rect 0 15600 1459 15602
rect 0 15544 1398 15600
rect 1454 15544 1459 15600
rect 0 15542 1459 15544
rect 0 15512 800 15542
rect 1393 15539 1459 15542
rect 16941 15602 17007 15605
rect 17401 15602 17467 15605
rect 16941 15600 17467 15602
rect 16941 15544 16946 15600
rect 17002 15544 17406 15600
rect 17462 15544 17467 15600
rect 16941 15542 17467 15544
rect 16941 15539 17007 15542
rect 17401 15539 17467 15542
rect 22001 15602 22067 15605
rect 22200 15602 23000 15632
rect 22001 15600 23000 15602
rect 22001 15544 22006 15600
rect 22062 15544 23000 15600
rect 22001 15542 23000 15544
rect 22001 15539 22067 15542
rect 22200 15512 23000 15542
rect 6453 15466 6519 15469
rect 13813 15466 13879 15469
rect 6453 15464 13879 15466
rect 6453 15408 6458 15464
rect 6514 15408 13818 15464
rect 13874 15408 13879 15464
rect 6453 15406 13879 15408
rect 6453 15403 6519 15406
rect 13813 15403 13879 15406
rect 14641 15466 14707 15469
rect 17769 15466 17835 15469
rect 14641 15464 17835 15466
rect 14641 15408 14646 15464
rect 14702 15408 17774 15464
rect 17830 15408 17835 15464
rect 14641 15406 17835 15408
rect 14641 15403 14707 15406
rect 17769 15403 17835 15406
rect 11881 15330 11947 15333
rect 16205 15330 16271 15333
rect 11881 15328 16271 15330
rect 11881 15272 11886 15328
rect 11942 15272 16210 15328
rect 16266 15272 16271 15328
rect 11881 15270 16271 15272
rect 11881 15267 11947 15270
rect 16205 15267 16271 15270
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1853 15194 1919 15197
rect 22200 15194 23000 15224
rect 0 15192 1919 15194
rect 0 15136 1858 15192
rect 1914 15136 1919 15192
rect 0 15134 1919 15136
rect 0 15104 800 15134
rect 1853 15131 1919 15134
rect 22142 15104 23000 15194
rect 3785 15058 3851 15061
rect 4337 15058 4403 15061
rect 6637 15058 6703 15061
rect 15101 15058 15167 15061
rect 3785 15056 15167 15058
rect 3785 15000 3790 15056
rect 3846 15000 4342 15056
rect 4398 15000 6642 15056
rect 6698 15000 15106 15056
rect 15162 15000 15167 15056
rect 3785 14998 15167 15000
rect 3785 14995 3851 14998
rect 4337 14995 4403 14998
rect 6637 14995 6703 14998
rect 15101 14995 15167 14998
rect 21449 15058 21515 15061
rect 22142 15058 22202 15104
rect 21449 15056 22202 15058
rect 21449 15000 21454 15056
rect 21510 15000 22202 15056
rect 21449 14998 22202 15000
rect 21449 14995 21515 14998
rect 2221 14922 2287 14925
rect 13997 14922 14063 14925
rect 2221 14920 14063 14922
rect 2221 14864 2226 14920
rect 2282 14864 14002 14920
rect 14058 14864 14063 14920
rect 2221 14862 14063 14864
rect 2221 14859 2287 14862
rect 13997 14859 14063 14862
rect 14457 14922 14523 14925
rect 16982 14922 16988 14924
rect 14457 14920 16988 14922
rect 14457 14864 14462 14920
rect 14518 14864 16988 14920
rect 14457 14862 16988 14864
rect 14457 14859 14523 14862
rect 16982 14860 16988 14862
rect 17052 14860 17058 14924
rect 0 14786 800 14816
rect 2865 14786 2931 14789
rect 0 14784 2931 14786
rect 0 14728 2870 14784
rect 2926 14728 2931 14784
rect 0 14726 2931 14728
rect 0 14696 800 14726
rect 2865 14723 2931 14726
rect 21541 14786 21607 14789
rect 22200 14786 23000 14816
rect 21541 14784 23000 14786
rect 21541 14728 21546 14784
rect 21602 14728 23000 14784
rect 21541 14726 23000 14728
rect 21541 14723 21607 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 9673 14650 9739 14653
rect 10409 14650 10475 14653
rect 12198 14650 12204 14652
rect 9673 14648 12204 14650
rect 9673 14592 9678 14648
rect 9734 14592 10414 14648
rect 10470 14592 12204 14648
rect 9673 14590 12204 14592
rect 9673 14587 9739 14590
rect 10409 14587 10475 14590
rect 12198 14588 12204 14590
rect 12268 14650 12274 14652
rect 14825 14650 14891 14653
rect 15101 14650 15167 14653
rect 12268 14590 13738 14650
rect 12268 14588 12274 14590
rect 12341 14514 12407 14517
rect 12525 14514 12591 14517
rect 12341 14512 12591 14514
rect 12341 14456 12346 14512
rect 12402 14456 12530 14512
rect 12586 14456 12591 14512
rect 12341 14454 12591 14456
rect 13678 14514 13738 14590
rect 14825 14648 15167 14650
rect 14825 14592 14830 14648
rect 14886 14592 15106 14648
rect 15162 14592 15167 14648
rect 14825 14590 15167 14592
rect 14825 14587 14891 14590
rect 15101 14587 15167 14590
rect 17401 14514 17467 14517
rect 13678 14512 17467 14514
rect 13678 14456 17406 14512
rect 17462 14456 17467 14512
rect 13678 14454 17467 14456
rect 12341 14451 12407 14454
rect 12525 14451 12591 14454
rect 17401 14451 17467 14454
rect 0 14378 800 14408
rect 2313 14378 2379 14381
rect 0 14376 2379 14378
rect 0 14320 2318 14376
rect 2374 14320 2379 14376
rect 0 14318 2379 14320
rect 0 14288 800 14318
rect 2313 14315 2379 14318
rect 8293 14378 8359 14381
rect 16021 14378 16087 14381
rect 8293 14376 16087 14378
rect 8293 14320 8298 14376
rect 8354 14320 16026 14376
rect 16082 14320 16087 14376
rect 8293 14318 16087 14320
rect 8293 14315 8359 14318
rect 16021 14315 16087 14318
rect 20897 14378 20963 14381
rect 22200 14378 23000 14408
rect 20897 14376 23000 14378
rect 20897 14320 20902 14376
rect 20958 14320 23000 14376
rect 20897 14318 23000 14320
rect 20897 14315 20963 14318
rect 22200 14288 23000 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 10777 14106 10843 14109
rect 10777 14104 11162 14106
rect 10777 14048 10782 14104
rect 10838 14048 11162 14104
rect 10777 14046 11162 14048
rect 10777 14043 10843 14046
rect 0 13970 800 14000
rect 0 13910 2790 13970
rect 0 13880 800 13910
rect 2730 13834 2790 13910
rect 2957 13834 3023 13837
rect 2730 13832 3023 13834
rect 2730 13776 2962 13832
rect 3018 13776 3023 13832
rect 2730 13774 3023 13776
rect 2957 13771 3023 13774
rect 5758 13772 5764 13836
rect 5828 13834 5834 13836
rect 6361 13834 6427 13837
rect 5828 13832 6427 13834
rect 5828 13776 6366 13832
rect 6422 13776 6427 13832
rect 5828 13774 6427 13776
rect 11102 13834 11162 14046
rect 13813 13970 13879 13973
rect 19425 13970 19491 13973
rect 13813 13968 19491 13970
rect 13813 13912 13818 13968
rect 13874 13912 19430 13968
rect 19486 13912 19491 13968
rect 13813 13910 19491 13912
rect 13813 13907 13879 13910
rect 19425 13907 19491 13910
rect 21357 13970 21423 13973
rect 22200 13970 23000 14000
rect 21357 13968 23000 13970
rect 21357 13912 21362 13968
rect 21418 13912 23000 13968
rect 21357 13910 23000 13912
rect 21357 13907 21423 13910
rect 22200 13880 23000 13910
rect 13537 13834 13603 13837
rect 11102 13832 13603 13834
rect 11102 13776 13542 13832
rect 13598 13776 13603 13832
rect 11102 13774 13603 13776
rect 5828 13772 5834 13774
rect 6361 13771 6427 13774
rect 13537 13771 13603 13774
rect 15142 13772 15148 13836
rect 15212 13834 15218 13836
rect 18965 13834 19031 13837
rect 15212 13832 19031 13834
rect 15212 13776 18970 13832
rect 19026 13776 19031 13832
rect 15212 13774 19031 13776
rect 15212 13772 15218 13774
rect 18965 13771 19031 13774
rect 14825 13698 14891 13701
rect 18137 13698 18203 13701
rect 14825 13696 18203 13698
rect 14825 13640 14830 13696
rect 14886 13640 18142 13696
rect 18198 13640 18203 13696
rect 14825 13638 18203 13640
rect 14825 13635 14891 13638
rect 18137 13635 18203 13638
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 3325 13562 3391 13565
rect 0 13560 3391 13562
rect 0 13504 3330 13560
rect 3386 13504 3391 13560
rect 0 13502 3391 13504
rect 0 13472 800 13502
rect 3325 13499 3391 13502
rect 21633 13562 21699 13565
rect 22200 13562 23000 13592
rect 21633 13560 23000 13562
rect 21633 13504 21638 13560
rect 21694 13504 23000 13560
rect 21633 13502 23000 13504
rect 21633 13499 21699 13502
rect 22200 13472 23000 13502
rect 11053 13426 11119 13429
rect 19793 13426 19859 13429
rect 11053 13424 19859 13426
rect 11053 13368 11058 13424
rect 11114 13368 19798 13424
rect 19854 13368 19859 13424
rect 11053 13366 19859 13368
rect 11053 13363 11119 13366
rect 19793 13363 19859 13366
rect 12566 13290 12572 13292
rect 2638 13230 12572 13290
rect 0 13154 800 13184
rect 2638 13154 2698 13230
rect 12566 13228 12572 13230
rect 12636 13228 12642 13292
rect 21173 13290 21239 13293
rect 21173 13288 22202 13290
rect 21173 13232 21178 13288
rect 21234 13232 22202 13288
rect 21173 13230 22202 13232
rect 21173 13227 21239 13230
rect 22142 13184 22202 13230
rect 6821 13156 6887 13157
rect 6821 13154 6868 13156
rect 0 13094 2698 13154
rect 6776 13152 6868 13154
rect 6776 13096 6826 13152
rect 6776 13094 6868 13096
rect 0 13064 800 13094
rect 6821 13092 6868 13094
rect 6932 13092 6938 13156
rect 22142 13094 23000 13184
rect 6821 13091 6887 13092
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 2497 13018 2563 13021
rect 4654 13018 4660 13020
rect 2497 13016 4660 13018
rect 2497 12960 2502 13016
rect 2558 12960 4660 13016
rect 2497 12958 4660 12960
rect 2497 12955 2563 12958
rect 4654 12956 4660 12958
rect 4724 12956 4730 13020
rect 12433 13018 12499 13021
rect 12750 13018 12756 13020
rect 6686 12958 8034 13018
rect 4429 12882 4495 12885
rect 6686 12882 6746 12958
rect 4429 12880 6746 12882
rect 4429 12824 4434 12880
rect 4490 12824 6746 12880
rect 4429 12822 6746 12824
rect 7974 12882 8034 12958
rect 12433 13016 12756 13018
rect 12433 12960 12438 13016
rect 12494 12960 12756 13016
rect 12433 12958 12756 12960
rect 12433 12955 12499 12958
rect 12750 12956 12756 12958
rect 12820 12956 12826 13020
rect 13445 13018 13511 13021
rect 13813 13018 13879 13021
rect 13445 13016 13879 13018
rect 13445 12960 13450 13016
rect 13506 12960 13818 13016
rect 13874 12960 13879 13016
rect 13445 12958 13879 12960
rect 13445 12955 13511 12958
rect 13813 12955 13879 12958
rect 17493 12882 17559 12885
rect 17861 12882 17927 12885
rect 7974 12822 17418 12882
rect 4429 12819 4495 12822
rect 0 12746 800 12776
rect 13445 12746 13511 12749
rect 0 12744 13511 12746
rect 0 12688 13450 12744
rect 13506 12688 13511 12744
rect 0 12686 13511 12688
rect 17358 12746 17418 12822
rect 17493 12880 17927 12882
rect 17493 12824 17498 12880
rect 17554 12824 17866 12880
rect 17922 12824 17927 12880
rect 17493 12822 17927 12824
rect 17493 12819 17559 12822
rect 17861 12819 17927 12822
rect 18137 12882 18203 12885
rect 21173 12882 21239 12885
rect 18137 12880 21239 12882
rect 18137 12824 18142 12880
rect 18198 12824 21178 12880
rect 21234 12824 21239 12880
rect 18137 12822 21239 12824
rect 18137 12819 18203 12822
rect 21173 12819 21239 12822
rect 22200 12746 23000 12776
rect 17358 12686 23000 12746
rect 0 12656 800 12686
rect 13445 12683 13511 12686
rect 22200 12656 23000 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 14590 12412 14596 12476
rect 14660 12474 14666 12476
rect 14733 12474 14799 12477
rect 14660 12472 14799 12474
rect 14660 12416 14738 12472
rect 14794 12416 14799 12472
rect 14660 12414 14799 12416
rect 14660 12412 14666 12414
rect 14733 12411 14799 12414
rect 0 12338 800 12368
rect 4521 12338 4587 12341
rect 4654 12338 4660 12340
rect 0 12278 2790 12338
rect 0 12248 800 12278
rect 2730 12202 2790 12278
rect 4521 12336 4660 12338
rect 4521 12280 4526 12336
rect 4582 12280 4660 12336
rect 4521 12278 4660 12280
rect 4521 12275 4587 12278
rect 4654 12276 4660 12278
rect 4724 12338 4730 12340
rect 20069 12338 20135 12341
rect 22200 12338 23000 12368
rect 4724 12336 20135 12338
rect 4724 12280 20074 12336
rect 20130 12280 20135 12336
rect 4724 12278 20135 12280
rect 4724 12276 4730 12278
rect 20069 12275 20135 12278
rect 20302 12278 23000 12338
rect 16113 12202 16179 12205
rect 19425 12202 19491 12205
rect 2730 12200 16179 12202
rect 2730 12144 16118 12200
rect 16174 12144 16179 12200
rect 2730 12142 16179 12144
rect 16113 12139 16179 12142
rect 16254 12200 19491 12202
rect 16254 12144 19430 12200
rect 19486 12144 19491 12200
rect 16254 12142 19491 12144
rect 11973 12066 12039 12069
rect 16254 12066 16314 12142
rect 19425 12139 19491 12142
rect 11973 12064 16314 12066
rect 11973 12008 11978 12064
rect 12034 12008 16314 12064
rect 11973 12006 16314 12008
rect 11973 12003 12039 12006
rect 17902 12004 17908 12068
rect 17972 12066 17978 12068
rect 20302 12066 20362 12278
rect 22200 12248 23000 12278
rect 17972 12006 20362 12066
rect 17972 12004 17978 12006
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 5533 11930 5599 11933
rect 5758 11930 5764 11932
rect 0 11870 2790 11930
rect 0 11840 800 11870
rect 2730 11794 2790 11870
rect 5533 11928 5764 11930
rect 5533 11872 5538 11928
rect 5594 11872 5764 11928
rect 5533 11870 5764 11872
rect 5533 11867 5599 11870
rect 5758 11868 5764 11870
rect 5828 11868 5834 11932
rect 22200 11930 23000 11960
rect 22142 11840 23000 11930
rect 3049 11794 3115 11797
rect 2730 11792 3115 11794
rect 2730 11736 3054 11792
rect 3110 11736 3115 11792
rect 2730 11734 3115 11736
rect 3049 11731 3115 11734
rect 9254 11732 9260 11796
rect 9324 11794 9330 11796
rect 14273 11794 14339 11797
rect 9324 11792 14339 11794
rect 9324 11736 14278 11792
rect 14334 11736 14339 11792
rect 9324 11734 14339 11736
rect 9324 11732 9330 11734
rect 14273 11731 14339 11734
rect 16113 11794 16179 11797
rect 19793 11794 19859 11797
rect 16113 11792 19859 11794
rect 16113 11736 16118 11792
rect 16174 11736 19798 11792
rect 19854 11736 19859 11792
rect 16113 11734 19859 11736
rect 16113 11731 16179 11734
rect 19793 11731 19859 11734
rect 20069 11794 20135 11797
rect 22142 11794 22202 11840
rect 20069 11792 22202 11794
rect 20069 11736 20074 11792
rect 20130 11736 22202 11792
rect 20069 11734 22202 11736
rect 20069 11731 20135 11734
rect 7005 11658 7071 11661
rect 11973 11658 12039 11661
rect 15469 11658 15535 11661
rect 18229 11658 18295 11661
rect 7005 11656 12039 11658
rect 7005 11600 7010 11656
rect 7066 11600 11978 11656
rect 12034 11600 12039 11656
rect 7005 11598 12039 11600
rect 7005 11595 7071 11598
rect 11973 11595 12039 11598
rect 12390 11656 18295 11658
rect 12390 11600 15474 11656
rect 15530 11600 18234 11656
rect 18290 11600 18295 11656
rect 12390 11598 18295 11600
rect 0 11522 800 11552
rect 3417 11522 3483 11525
rect 0 11520 3483 11522
rect 0 11464 3422 11520
rect 3478 11464 3483 11520
rect 0 11462 3483 11464
rect 0 11432 800 11462
rect 3417 11459 3483 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 12390 11386 12450 11598
rect 15469 11595 15535 11598
rect 18229 11595 18295 11598
rect 18413 11658 18479 11661
rect 18413 11656 19626 11658
rect 18413 11600 18418 11656
rect 18474 11600 19626 11656
rect 18413 11598 19626 11600
rect 18413 11595 18479 11598
rect 19566 11522 19626 11598
rect 22200 11522 23000 11552
rect 19566 11462 23000 11522
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 11102 11326 12450 11386
rect 11102 11253 11162 11326
rect 3918 11188 3924 11252
rect 3988 11250 3994 11252
rect 4429 11250 4495 11253
rect 3988 11248 4495 11250
rect 3988 11192 4434 11248
rect 4490 11192 4495 11248
rect 3988 11190 4495 11192
rect 3988 11188 3994 11190
rect 4429 11187 4495 11190
rect 11053 11248 11162 11253
rect 17309 11250 17375 11253
rect 11053 11192 11058 11248
rect 11114 11192 11162 11248
rect 11053 11190 11162 11192
rect 11286 11248 17375 11250
rect 11286 11192 17314 11248
rect 17370 11192 17375 11248
rect 11286 11190 17375 11192
rect 11053 11187 11119 11190
rect 0 11114 800 11144
rect 3785 11114 3851 11117
rect 0 11112 3851 11114
rect 0 11056 3790 11112
rect 3846 11056 3851 11112
rect 0 11054 3851 11056
rect 0 11024 800 11054
rect 3785 11051 3851 11054
rect 5073 11114 5139 11117
rect 11286 11114 11346 11190
rect 17309 11187 17375 11190
rect 18229 11252 18295 11253
rect 18229 11248 18276 11252
rect 18340 11250 18346 11252
rect 18229 11192 18234 11248
rect 18229 11188 18276 11192
rect 18340 11190 18386 11250
rect 18340 11188 18346 11190
rect 18229 11187 18295 11188
rect 5073 11112 11346 11114
rect 5073 11056 5078 11112
rect 5134 11056 11346 11112
rect 5073 11054 11346 11056
rect 11881 11114 11947 11117
rect 12893 11114 12959 11117
rect 11881 11112 12959 11114
rect 11881 11056 11886 11112
rect 11942 11056 12898 11112
rect 12954 11056 12959 11112
rect 11881 11054 12959 11056
rect 5073 11051 5139 11054
rect 11881 11051 11947 11054
rect 12893 11051 12959 11054
rect 13353 11114 13419 11117
rect 17902 11114 17908 11116
rect 13353 11112 17908 11114
rect 13353 11056 13358 11112
rect 13414 11056 17908 11112
rect 13353 11054 17908 11056
rect 13353 11051 13419 11054
rect 17902 11052 17908 11054
rect 17972 11052 17978 11116
rect 18638 11052 18644 11116
rect 18708 11114 18714 11116
rect 22200 11114 23000 11144
rect 18708 11054 23000 11114
rect 18708 11052 18714 11054
rect 22200 11024 23000 11054
rect 19977 10978 20043 10981
rect 20345 10978 20411 10981
rect 21449 10978 21515 10981
rect 19977 10976 21515 10978
rect 19977 10920 19982 10976
rect 20038 10920 20350 10976
rect 20406 10920 21454 10976
rect 21510 10920 21515 10976
rect 19977 10918 21515 10920
rect 19977 10915 20043 10918
rect 20345 10915 20411 10918
rect 21449 10915 21515 10918
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 17953 10842 18019 10845
rect 17953 10840 21282 10842
rect 17953 10784 17958 10840
rect 18014 10784 21282 10840
rect 17953 10782 21282 10784
rect 17953 10779 18019 10782
rect 0 10706 800 10736
rect 2865 10706 2931 10709
rect 0 10704 2931 10706
rect 0 10648 2870 10704
rect 2926 10648 2931 10704
rect 0 10646 2931 10648
rect 0 10616 800 10646
rect 2865 10643 2931 10646
rect 3049 10706 3115 10709
rect 20989 10706 21055 10709
rect 3049 10704 21055 10706
rect 3049 10648 3054 10704
rect 3110 10648 20994 10704
rect 21050 10648 21055 10704
rect 3049 10646 21055 10648
rect 21222 10706 21282 10782
rect 22200 10706 23000 10736
rect 21222 10646 23000 10706
rect 3049 10643 3115 10646
rect 20989 10643 21055 10646
rect 22200 10616 23000 10646
rect 8845 10570 8911 10573
rect 11973 10570 12039 10573
rect 8845 10568 12039 10570
rect 8845 10512 8850 10568
rect 8906 10512 11978 10568
rect 12034 10512 12039 10568
rect 8845 10510 12039 10512
rect 8845 10507 8911 10510
rect 11973 10507 12039 10510
rect 12617 10570 12683 10573
rect 16573 10570 16639 10573
rect 12617 10568 16639 10570
rect 12617 10512 12622 10568
rect 12678 10512 16578 10568
rect 16634 10512 16639 10568
rect 12617 10510 16639 10512
rect 12617 10507 12683 10510
rect 16573 10507 16639 10510
rect 17585 10570 17651 10573
rect 17585 10568 19626 10570
rect 17585 10512 17590 10568
rect 17646 10512 19626 10568
rect 17585 10510 19626 10512
rect 17585 10507 17651 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 3366 10298 3372 10300
rect 0 10238 3372 10298
rect 0 10208 800 10238
rect 3366 10236 3372 10238
rect 3436 10236 3442 10300
rect 10041 10298 10107 10301
rect 11513 10298 11579 10301
rect 10041 10296 11579 10298
rect 10041 10240 10046 10296
rect 10102 10240 11518 10296
rect 11574 10240 11579 10296
rect 10041 10238 11579 10240
rect 19566 10298 19626 10510
rect 22200 10298 23000 10328
rect 19566 10238 23000 10298
rect 10041 10235 10107 10238
rect 11513 10235 11579 10238
rect 22200 10208 23000 10238
rect 7465 10162 7531 10165
rect 17585 10162 17651 10165
rect 7465 10160 17651 10162
rect 7465 10104 7470 10160
rect 7526 10104 17590 10160
rect 17646 10104 17651 10160
rect 7465 10102 17651 10104
rect 7465 10099 7531 10102
rect 17585 10099 17651 10102
rect 11329 10026 11395 10029
rect 12249 10026 12315 10029
rect 16113 10026 16179 10029
rect 11329 10024 16179 10026
rect 11329 9968 11334 10024
rect 11390 9968 12254 10024
rect 12310 9968 16118 10024
rect 16174 9968 16179 10024
rect 11329 9966 16179 9968
rect 11329 9963 11395 9966
rect 12249 9963 12315 9966
rect 16113 9963 16179 9966
rect 18321 10026 18387 10029
rect 18321 10024 22202 10026
rect 18321 9968 18326 10024
rect 18382 9968 22202 10024
rect 18321 9966 22202 9968
rect 18321 9963 18387 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 3877 9890 3943 9893
rect 0 9888 3943 9890
rect 0 9832 3882 9888
rect 3938 9832 3943 9888
rect 0 9830 3943 9832
rect 22142 9830 23000 9920
rect 0 9800 800 9830
rect 3877 9827 3943 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 2957 9690 3023 9693
rect 2638 9688 3023 9690
rect 2638 9632 2962 9688
rect 3018 9632 3023 9688
rect 2638 9630 3023 9632
rect 2221 9618 2287 9621
rect 2638 9618 2698 9630
rect 2957 9627 3023 9630
rect 2221 9616 2698 9618
rect 2221 9560 2226 9616
rect 2282 9560 2698 9616
rect 2221 9558 2698 9560
rect 3693 9618 3759 9621
rect 3918 9618 3924 9620
rect 3693 9616 3924 9618
rect 3693 9560 3698 9616
rect 3754 9560 3924 9616
rect 3693 9558 3924 9560
rect 2221 9555 2287 9558
rect 3693 9555 3759 9558
rect 3918 9556 3924 9558
rect 3988 9556 3994 9620
rect 5165 9618 5231 9621
rect 5349 9618 5415 9621
rect 5165 9616 5415 9618
rect 5165 9560 5170 9616
rect 5226 9560 5354 9616
rect 5410 9560 5415 9616
rect 5165 9558 5415 9560
rect 5165 9555 5231 9558
rect 5349 9555 5415 9558
rect 9673 9618 9739 9621
rect 17677 9618 17743 9621
rect 19241 9618 19307 9621
rect 9673 9616 17743 9618
rect 9673 9560 9678 9616
rect 9734 9560 17682 9616
rect 17738 9560 17743 9616
rect 9673 9558 17743 9560
rect 9673 9555 9739 9558
rect 17677 9555 17743 9558
rect 18646 9616 19307 9618
rect 18646 9560 19246 9616
rect 19302 9560 19307 9616
rect 18646 9558 19307 9560
rect 0 9482 800 9512
rect 18646 9485 18706 9558
rect 19241 9555 19307 9558
rect 3969 9482 4035 9485
rect 0 9480 4035 9482
rect 0 9424 3974 9480
rect 4030 9424 4035 9480
rect 0 9422 4035 9424
rect 0 9392 800 9422
rect 3969 9419 4035 9422
rect 11053 9482 11119 9485
rect 18229 9482 18295 9485
rect 18597 9482 18706 9485
rect 11053 9480 18706 9482
rect 11053 9424 11058 9480
rect 11114 9424 18234 9480
rect 18290 9424 18602 9480
rect 18658 9424 18706 9480
rect 11053 9422 18706 9424
rect 18781 9482 18847 9485
rect 22200 9482 23000 9512
rect 18781 9480 23000 9482
rect 18781 9424 18786 9480
rect 18842 9424 23000 9480
rect 18781 9422 23000 9424
rect 11053 9419 11119 9422
rect 18229 9419 18295 9422
rect 18597 9419 18663 9422
rect 18781 9419 18847 9422
rect 22200 9392 23000 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 4337 9074 4403 9077
rect 0 9072 4403 9074
rect 0 9016 4342 9072
rect 4398 9016 4403 9072
rect 0 9014 4403 9016
rect 0 8984 800 9014
rect 4337 9011 4403 9014
rect 6545 9074 6611 9077
rect 15101 9074 15167 9077
rect 6545 9072 15167 9074
rect 6545 9016 6550 9072
rect 6606 9016 15106 9072
rect 15162 9016 15167 9072
rect 6545 9014 15167 9016
rect 6545 9011 6611 9014
rect 15101 9011 15167 9014
rect 18689 9074 18755 9077
rect 22200 9074 23000 9104
rect 18689 9072 23000 9074
rect 18689 9016 18694 9072
rect 18750 9016 23000 9072
rect 18689 9014 23000 9016
rect 18689 9011 18755 9014
rect 22200 8984 23000 9014
rect 7373 8938 7439 8941
rect 15837 8938 15903 8941
rect 7373 8936 15903 8938
rect 7373 8880 7378 8936
rect 7434 8880 15842 8936
rect 15898 8880 15903 8936
rect 7373 8878 15903 8880
rect 7373 8875 7439 8878
rect 15837 8875 15903 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 3969 8666 4035 8669
rect 22200 8666 23000 8696
rect 0 8664 4035 8666
rect 0 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 3969 8603 4035 8606
rect 22142 8576 23000 8666
rect 9581 8530 9647 8533
rect 14089 8530 14155 8533
rect 9581 8528 14155 8530
rect 9581 8472 9586 8528
rect 9642 8472 14094 8528
rect 14150 8472 14155 8528
rect 9581 8470 14155 8472
rect 9581 8467 9647 8470
rect 14089 8467 14155 8470
rect 16297 8530 16363 8533
rect 22142 8530 22202 8576
rect 16297 8528 22202 8530
rect 16297 8472 16302 8528
rect 16358 8472 22202 8528
rect 16297 8470 22202 8472
rect 16297 8467 16363 8470
rect 4613 8394 4679 8397
rect 5349 8394 5415 8397
rect 6453 8394 6519 8397
rect 4613 8392 6519 8394
rect 4613 8336 4618 8392
rect 4674 8336 5354 8392
rect 5410 8336 6458 8392
rect 6514 8336 6519 8392
rect 4613 8334 6519 8336
rect 4613 8331 4679 8334
rect 5349 8331 5415 8334
rect 6453 8331 6519 8334
rect 9305 8394 9371 8397
rect 13813 8394 13879 8397
rect 9305 8392 13879 8394
rect 9305 8336 9310 8392
rect 9366 8336 13818 8392
rect 13874 8336 13879 8392
rect 9305 8334 13879 8336
rect 9305 8331 9371 8334
rect 13813 8331 13879 8334
rect 19149 8394 19215 8397
rect 19149 8392 19626 8394
rect 19149 8336 19154 8392
rect 19210 8336 19626 8392
rect 19149 8334 19626 8336
rect 19149 8331 19215 8334
rect 0 8258 800 8288
rect 19566 8258 19626 8334
rect 22200 8258 23000 8288
rect 0 8198 2790 8258
rect 19566 8198 23000 8258
rect 0 8168 800 8198
rect 2730 7986 2790 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 22200 8168 23000 8198
rect 19139 8127 19455 8128
rect 9121 8122 9187 8125
rect 19517 8124 19583 8125
rect 9121 8120 12450 8122
rect 9121 8064 9126 8120
rect 9182 8064 12450 8120
rect 9121 8062 12450 8064
rect 9121 8059 9187 8062
rect 12390 7986 12450 8062
rect 19517 8120 19564 8124
rect 19628 8122 19634 8124
rect 19517 8064 19522 8120
rect 19517 8060 19564 8064
rect 19628 8062 19674 8122
rect 19628 8060 19634 8062
rect 19517 8059 19583 8060
rect 16849 7986 16915 7989
rect 2730 7926 11898 7986
rect 12390 7984 16915 7986
rect 12390 7928 16854 7984
rect 16910 7928 16915 7984
rect 12390 7926 16915 7928
rect 0 7850 800 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 800 7790
rect 3969 7787 4035 7790
rect 5349 7850 5415 7853
rect 5993 7850 6059 7853
rect 5349 7848 6059 7850
rect 5349 7792 5354 7848
rect 5410 7792 5998 7848
rect 6054 7792 6059 7848
rect 5349 7790 6059 7792
rect 5349 7787 5415 7790
rect 5993 7787 6059 7790
rect 11838 7714 11898 7926
rect 16849 7923 16915 7926
rect 17677 7986 17743 7989
rect 17953 7986 18019 7989
rect 17677 7984 18019 7986
rect 17677 7928 17682 7984
rect 17738 7928 17958 7984
rect 18014 7928 18019 7984
rect 17677 7926 18019 7928
rect 17677 7923 17743 7926
rect 17953 7923 18019 7926
rect 11973 7850 12039 7853
rect 18086 7850 18092 7852
rect 11973 7848 18092 7850
rect 11973 7792 11978 7848
rect 12034 7792 18092 7848
rect 11973 7790 18092 7792
rect 11973 7787 12039 7790
rect 18086 7788 18092 7790
rect 18156 7850 18162 7852
rect 18781 7850 18847 7853
rect 18156 7848 18847 7850
rect 18156 7792 18786 7848
rect 18842 7792 18847 7848
rect 18156 7790 18847 7792
rect 18156 7788 18162 7790
rect 18781 7787 18847 7790
rect 18965 7850 19031 7853
rect 22200 7850 23000 7880
rect 18965 7848 23000 7850
rect 18965 7792 18970 7848
rect 19026 7792 23000 7848
rect 18965 7790 23000 7792
rect 18965 7787 19031 7790
rect 22200 7760 23000 7790
rect 11838 7654 12450 7714
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 12390 7578 12450 7654
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 15142 7578 15148 7580
rect 12390 7518 15148 7578
rect 15142 7516 15148 7518
rect 15212 7516 15218 7580
rect 0 7442 800 7472
rect 4061 7442 4127 7445
rect 0 7440 4127 7442
rect 0 7384 4066 7440
rect 4122 7384 4127 7440
rect 0 7382 4127 7384
rect 0 7352 800 7382
rect 4061 7379 4127 7382
rect 13721 7442 13787 7445
rect 22200 7442 23000 7472
rect 13721 7440 23000 7442
rect 13721 7384 13726 7440
rect 13782 7384 23000 7440
rect 13721 7382 23000 7384
rect 13721 7379 13787 7382
rect 22200 7352 23000 7382
rect 6729 7306 6795 7309
rect 17677 7306 17743 7309
rect 6729 7304 17743 7306
rect 6729 7248 6734 7304
rect 6790 7248 17682 7304
rect 17738 7248 17743 7304
rect 6729 7246 17743 7248
rect 6729 7243 6795 7246
rect 17677 7243 17743 7246
rect 18321 7306 18387 7309
rect 18321 7304 19626 7306
rect 18321 7248 18326 7304
rect 18382 7248 19626 7304
rect 18321 7246 19626 7248
rect 18321 7243 18387 7246
rect 18689 7172 18755 7173
rect 18638 7170 18644 7172
rect 18598 7110 18644 7170
rect 18708 7168 18755 7172
rect 18750 7112 18755 7168
rect 18638 7108 18644 7110
rect 18708 7108 18755 7112
rect 18689 7107 18755 7108
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 3233 7034 3299 7037
rect 0 7032 3299 7034
rect 0 6976 3238 7032
rect 3294 6976 3299 7032
rect 0 6974 3299 6976
rect 19566 7034 19626 7246
rect 22200 7034 23000 7064
rect 19566 6974 23000 7034
rect 0 6944 800 6974
rect 3233 6971 3299 6974
rect 22200 6944 23000 6974
rect 3366 6700 3372 6764
rect 3436 6762 3442 6764
rect 17401 6762 17467 6765
rect 3436 6760 17467 6762
rect 3436 6704 17406 6760
rect 17462 6704 17467 6760
rect 3436 6702 17467 6704
rect 3436 6700 3442 6702
rect 17401 6699 17467 6702
rect 18137 6762 18203 6765
rect 18137 6760 22202 6762
rect 18137 6704 18142 6760
rect 18198 6704 22202 6760
rect 18137 6702 22202 6704
rect 18137 6699 18203 6702
rect 22142 6656 22202 6702
rect 0 6626 800 6656
rect 4061 6626 4127 6629
rect 0 6624 4127 6626
rect 0 6568 4066 6624
rect 4122 6568 4127 6624
rect 0 6566 4127 6568
rect 22142 6566 23000 6656
rect 0 6536 800 6566
rect 4061 6563 4127 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 0 6218 800 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 800 6158
rect 3969 6155 4035 6158
rect 17953 6218 18019 6221
rect 22200 6218 23000 6248
rect 17953 6216 23000 6218
rect 17953 6160 17958 6216
rect 18014 6160 23000 6216
rect 17953 6158 23000 6160
rect 17953 6155 18019 6158
rect 22200 6128 23000 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 18505 5810 18571 5813
rect 22200 5810 23000 5840
rect 18505 5808 23000 5810
rect 18505 5752 18510 5808
rect 18566 5752 23000 5808
rect 18505 5750 23000 5752
rect 18505 5747 18571 5750
rect 22200 5720 23000 5750
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 4061 5402 4127 5405
rect 22200 5402 23000 5432
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 800 5342
rect 4061 5339 4127 5342
rect 22142 5312 23000 5402
rect 5809 5266 5875 5269
rect 6453 5266 6519 5269
rect 7281 5266 7347 5269
rect 7741 5266 7807 5269
rect 5809 5264 7807 5266
rect 5809 5208 5814 5264
rect 5870 5208 6458 5264
rect 6514 5208 7286 5264
rect 7342 5208 7746 5264
rect 7802 5208 7807 5264
rect 5809 5206 7807 5208
rect 5809 5203 5875 5206
rect 6453 5203 6519 5206
rect 7281 5203 7347 5206
rect 7741 5203 7807 5206
rect 17953 5266 18019 5269
rect 22142 5266 22202 5312
rect 17953 5264 22202 5266
rect 17953 5208 17958 5264
rect 18014 5208 22202 5264
rect 17953 5206 22202 5208
rect 17953 5203 18019 5206
rect 0 4994 800 5024
rect 2221 4994 2287 4997
rect 0 4992 2287 4994
rect 0 4936 2226 4992
rect 2282 4936 2287 4992
rect 0 4934 2287 4936
rect 0 4904 800 4934
rect 2221 4931 2287 4934
rect 21173 4994 21239 4997
rect 22200 4994 23000 5024
rect 21173 4992 23000 4994
rect 21173 4936 21178 4992
rect 21234 4936 23000 4992
rect 21173 4934 23000 4936
rect 21173 4931 21239 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 0 4586 800 4616
rect 3233 4586 3299 4589
rect 0 4584 3299 4586
rect 0 4528 3238 4584
rect 3294 4528 3299 4584
rect 0 4526 3299 4528
rect 0 4496 800 4526
rect 3233 4523 3299 4526
rect 20253 4586 20319 4589
rect 22200 4586 23000 4616
rect 20253 4584 23000 4586
rect 20253 4528 20258 4584
rect 20314 4528 23000 4584
rect 20253 4526 23000 4528
rect 20253 4523 20319 4526
rect 22200 4496 23000 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4178 800 4208
rect 2129 4178 2195 4181
rect 0 4176 2195 4178
rect 0 4120 2134 4176
rect 2190 4120 2195 4176
rect 0 4118 2195 4120
rect 0 4088 800 4118
rect 2129 4115 2195 4118
rect 20529 4178 20595 4181
rect 22200 4178 23000 4208
rect 20529 4176 23000 4178
rect 20529 4120 20534 4176
rect 20590 4120 23000 4176
rect 20529 4118 23000 4120
rect 20529 4115 20595 4118
rect 22200 4088 23000 4118
rect 5257 4042 5323 4045
rect 5390 4042 5396 4044
rect 5257 4040 5396 4042
rect 5257 3984 5262 4040
rect 5318 3984 5396 4040
rect 5257 3982 5396 3984
rect 5257 3979 5323 3982
rect 5390 3980 5396 3982
rect 5460 3980 5466 4044
rect 5758 3980 5764 4044
rect 5828 4042 5834 4044
rect 6821 4042 6887 4045
rect 5828 4040 6887 4042
rect 5828 3984 6826 4040
rect 6882 3984 6887 4040
rect 5828 3982 6887 3984
rect 5828 3980 5834 3982
rect 6821 3979 6887 3982
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 2313 3770 2379 3773
rect 0 3768 2379 3770
rect 0 3712 2318 3768
rect 2374 3712 2379 3768
rect 0 3710 2379 3712
rect 0 3680 800 3710
rect 2313 3707 2379 3710
rect 20345 3770 20411 3773
rect 22200 3770 23000 3800
rect 20345 3768 23000 3770
rect 20345 3712 20350 3768
rect 20406 3712 23000 3768
rect 20345 3710 23000 3712
rect 20345 3707 20411 3710
rect 22200 3680 23000 3710
rect 5942 3436 5948 3500
rect 6012 3498 6018 3500
rect 12249 3498 12315 3501
rect 6012 3496 12315 3498
rect 6012 3440 12254 3496
rect 12310 3440 12315 3496
rect 6012 3438 12315 3440
rect 6012 3436 6018 3438
rect 12249 3435 12315 3438
rect 20621 3498 20687 3501
rect 20621 3496 22202 3498
rect 20621 3440 20626 3496
rect 20682 3440 22202 3496
rect 20621 3438 22202 3440
rect 20621 3435 20687 3438
rect 22142 3392 22202 3438
rect 0 3362 800 3392
rect 3049 3362 3115 3365
rect 0 3360 3115 3362
rect 0 3304 3054 3360
rect 3110 3304 3115 3360
rect 0 3302 3115 3304
rect 22142 3302 23000 3392
rect 0 3272 800 3302
rect 3049 3299 3115 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 0 2954 800 2984
rect 3417 2954 3483 2957
rect 0 2952 3483 2954
rect 0 2896 3422 2952
rect 3478 2896 3483 2952
rect 0 2894 3483 2896
rect 0 2864 800 2894
rect 3417 2891 3483 2894
rect 20069 2954 20135 2957
rect 22200 2954 23000 2984
rect 20069 2952 23000 2954
rect 20069 2896 20074 2952
rect 20130 2896 23000 2952
rect 20069 2894 23000 2896
rect 20069 2891 20135 2894
rect 22200 2864 23000 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 0 2546 800 2576
rect 4613 2546 4679 2549
rect 0 2544 4679 2546
rect 0 2488 4618 2544
rect 4674 2488 4679 2544
rect 0 2486 4679 2488
rect 0 2456 800 2486
rect 4613 2483 4679 2486
rect 20529 2546 20595 2549
rect 22200 2546 23000 2576
rect 20529 2544 23000 2546
rect 20529 2488 20534 2544
rect 20590 2488 23000 2544
rect 20529 2486 23000 2488
rect 20529 2483 20595 2486
rect 22200 2456 23000 2486
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 4153 2138 4219 2141
rect 22200 2138 23000 2168
rect 0 2136 4219 2138
rect 0 2080 4158 2136
rect 4214 2080 4219 2136
rect 0 2078 4219 2080
rect 0 2048 800 2078
rect 4153 2075 4219 2078
rect 22142 2048 23000 2138
rect 20897 2002 20963 2005
rect 22142 2002 22202 2048
rect 20897 2000 22202 2002
rect 20897 1944 20902 2000
rect 20958 1944 22202 2000
rect 20897 1942 22202 1944
rect 20897 1939 20963 1942
rect 0 1730 800 1760
rect 4061 1730 4127 1733
rect 0 1728 4127 1730
rect 0 1672 4066 1728
rect 4122 1672 4127 1728
rect 0 1670 4127 1672
rect 0 1640 800 1670
rect 4061 1667 4127 1670
rect 19057 1730 19123 1733
rect 22200 1730 23000 1760
rect 19057 1728 23000 1730
rect 19057 1672 19062 1728
rect 19118 1672 23000 1728
rect 19057 1670 23000 1672
rect 19057 1667 19123 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 9260 20164 9324 20228
rect 16988 20300 17052 20364
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 17908 19892 17972 19956
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 6868 19348 6932 19412
rect 9628 19484 9692 19548
rect 12572 19620 12636 19684
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 12204 19076 12268 19140
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 19564 18940 19628 19004
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 12756 18124 12820 18188
rect 3372 17988 3436 18052
rect 5948 17988 6012 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 9628 17852 9692 17916
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 5396 17308 5460 17372
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 14596 16960 14660 16964
rect 18092 17036 18156 17100
rect 14596 16904 14610 16960
rect 14610 16904 14660 16960
rect 14596 16900 14660 16904
rect 18644 16960 18708 16964
rect 18644 16904 18694 16960
rect 18694 16904 18708 16960
rect 18644 16900 18708 16904
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 3372 16628 3436 16692
rect 18276 16492 18340 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 16988 14860 17052 14924
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 12204 14588 12268 14652
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 5764 13772 5828 13836
rect 15148 13772 15212 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 12572 13228 12636 13292
rect 6868 13152 6932 13156
rect 6868 13096 6882 13152
rect 6882 13096 6932 13152
rect 6868 13092 6932 13096
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 4660 12956 4724 13020
rect 12756 12956 12820 13020
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 14596 12412 14660 12476
rect 4660 12276 4724 12340
rect 17908 12004 17972 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 5764 11868 5828 11932
rect 9260 11732 9324 11796
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 3924 11188 3988 11252
rect 18276 11248 18340 11252
rect 18276 11192 18290 11248
rect 18290 11192 18340 11248
rect 18276 11188 18340 11192
rect 17908 11052 17972 11116
rect 18644 11052 18708 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 3372 10236 3436 10300
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3924 9556 3988 9620
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 19564 8120 19628 8124
rect 19564 8064 19578 8120
rect 19578 8064 19628 8120
rect 19564 8060 19628 8064
rect 18092 7788 18156 7852
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 15148 7516 15212 7580
rect 18644 7168 18708 7172
rect 18644 7112 18694 7168
rect 18694 7112 18708 7168
rect 18644 7108 18708 7112
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 3372 6700 3436 6764
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 5396 3980 5460 4044
rect 5764 3980 5828 4044
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 5948 3436 6012 3500
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3371 18052 3437 18053
rect 3371 17988 3372 18052
rect 3436 17988 3437 18052
rect 3371 17987 3437 17988
rect 3374 16693 3434 17987
rect 3543 17984 3863 19008
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 8741 20160 9061 20720
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 9259 20228 9325 20229
rect 9259 20164 9260 20228
rect 9324 20164 9325 20228
rect 9259 20163 9325 20164
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 6867 19412 6933 19413
rect 6867 19348 6868 19412
rect 6932 19348 6933 19412
rect 6867 19347 6933 19348
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5947 18052 6013 18053
rect 5947 17988 5948 18052
rect 6012 17988 6013 18052
rect 5947 17987 6013 17988
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 5395 17372 5461 17373
rect 5395 17308 5396 17372
rect 5460 17308 5461 17372
rect 5395 17307 5461 17308
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3371 16692 3437 16693
rect 3371 16628 3372 16692
rect 3436 16628 3437 16692
rect 3371 16627 3437 16628
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 4659 13020 4725 13021
rect 4659 12956 4660 13020
rect 4724 12956 4725 13020
rect 4659 12955 4725 12956
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 4662 12341 4722 12955
rect 4659 12340 4725 12341
rect 4659 12276 4660 12340
rect 4724 12276 4725 12340
rect 4659 12275 4725 12276
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3923 11252 3989 11253
rect 3923 11188 3924 11252
rect 3988 11188 3989 11252
rect 3923 11187 3989 11188
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3371 10300 3437 10301
rect 3371 10236 3372 10300
rect 3436 10236 3437 10300
rect 3371 10235 3437 10236
rect 3374 6765 3434 10235
rect 3543 9280 3863 10304
rect 3926 9621 3986 11187
rect 3923 9620 3989 9621
rect 3923 9556 3924 9620
rect 3988 9556 3989 9620
rect 3923 9555 3989 9556
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3371 6764 3437 6765
rect 3371 6700 3372 6764
rect 3436 6700 3437 6764
rect 3371 6699 3437 6700
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 5398 4045 5458 17307
rect 5763 13836 5829 13837
rect 5763 13772 5764 13836
rect 5828 13772 5829 13836
rect 5763 13771 5829 13772
rect 5766 11933 5826 13771
rect 5763 11932 5829 11933
rect 5763 11868 5764 11932
rect 5828 11868 5829 11932
rect 5763 11867 5829 11868
rect 5766 4045 5826 11867
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 5763 4044 5829 4045
rect 5763 3980 5764 4044
rect 5828 3980 5829 4044
rect 5763 3979 5829 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 5950 3501 6010 17987
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6870 13157 6930 19347
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 6867 13156 6933 13157
rect 6867 13092 6868 13156
rect 6932 13092 6933 13156
rect 6867 13091 6933 13092
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 3500 6013 3501
rect 5947 3436 5948 3500
rect 6012 3436 6013 3500
rect 5947 3435 6013 3436
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 9262 11797 9322 20163
rect 11340 19616 11660 20640
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 12571 19684 12637 19685
rect 12571 19620 12572 19684
rect 12636 19620 12637 19684
rect 12571 19619 12637 19620
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 9627 19548 9693 19549
rect 9627 19484 9628 19548
rect 9692 19484 9693 19548
rect 9627 19483 9693 19484
rect 9630 17917 9690 19483
rect 11340 18528 11660 19552
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9627 17916 9693 17917
rect 9627 17852 9628 17916
rect 9692 17852 9693 17916
rect 9627 17851 9693 17852
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 12206 14653 12266 19075
rect 12203 14652 12269 14653
rect 12203 14588 12204 14652
rect 12268 14588 12269 14652
rect 12203 14587 12269 14588
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 12574 13293 12634 19619
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 12755 18188 12821 18189
rect 12755 18124 12756 18188
rect 12820 18124 12821 18188
rect 12755 18123 12821 18124
rect 12571 13292 12637 13293
rect 12571 13228 12572 13292
rect 12636 13228 12637 13292
rect 12571 13227 12637 13228
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 12758 13021 12818 18123
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16987 20364 17053 20365
rect 16987 20300 16988 20364
rect 17052 20300 17053 20364
rect 16987 20299 17053 20300
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 14595 16964 14661 16965
rect 14595 16900 14596 16964
rect 14660 16900 14661 16964
rect 14595 16899 14661 16900
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 12755 13020 12821 13021
rect 12755 12956 12756 13020
rect 12820 12956 12821 13020
rect 12755 12955 12821 12956
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 9259 11796 9325 11797
rect 9259 11732 9260 11796
rect 9324 11732 9325 11796
rect 9259 11731 9325 11732
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 14598 12477 14658 16899
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16990 14925 17050 20299
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 17907 19956 17973 19957
rect 17907 19892 17908 19956
rect 17972 19892 17973 19956
rect 17907 19891 17973 19892
rect 16987 14924 17053 14925
rect 16987 14860 16988 14924
rect 17052 14860 17053 14924
rect 16987 14859 17053 14860
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 15147 13836 15213 13837
rect 15147 13772 15148 13836
rect 15212 13772 15213 13836
rect 15147 13771 15213 13772
rect 14595 12476 14661 12477
rect 14595 12412 14596 12476
rect 14660 12412 14661 12476
rect 14595 12411 14661 12412
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 15150 7581 15210 13771
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 17910 12069 17970 19891
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 19563 19004 19629 19005
rect 19563 18940 19564 19004
rect 19628 18940 19629 19004
rect 19563 18939 19629 18940
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 18091 17100 18157 17101
rect 18091 17036 18092 17100
rect 18156 17036 18157 17100
rect 18091 17035 18157 17036
rect 17907 12068 17973 12069
rect 17907 12004 17908 12068
rect 17972 12004 17973 12068
rect 17907 12003 17973 12004
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 17910 11117 17970 12003
rect 17907 11116 17973 11117
rect 17907 11052 17908 11116
rect 17972 11052 17973 11116
rect 17907 11051 17973 11052
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 18094 7853 18154 17035
rect 18643 16964 18709 16965
rect 18643 16900 18644 16964
rect 18708 16900 18709 16964
rect 18643 16899 18709 16900
rect 18275 16556 18341 16557
rect 18275 16492 18276 16556
rect 18340 16492 18341 16556
rect 18275 16491 18341 16492
rect 18278 11253 18338 16491
rect 18275 11252 18341 11253
rect 18275 11188 18276 11252
rect 18340 11188 18341 11252
rect 18275 11187 18341 11188
rect 18646 11117 18706 16899
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 18643 11116 18709 11117
rect 18643 11052 18644 11116
rect 18708 11052 18709 11116
rect 18643 11051 18709 11052
rect 18091 7852 18157 7853
rect 18091 7788 18092 7852
rect 18156 7788 18157 7852
rect 18091 7787 18157 7788
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 6560 16858 7584
rect 18646 7173 18706 11051
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 18643 7172 18709 7173
rect 18643 7108 18644 7172
rect 18708 7108 18709 7172
rect 18643 7107 18709 7108
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 7104 19457 8128
rect 19566 8125 19626 18939
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 19563 8124 19629 8125
rect 19563 8060 19564 8124
rect 19628 8060 19629 8124
rect 19563 8059 19629 8060
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1649977179
transform -1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform -1 0 2944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform 1 0 2944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 1840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform -1 0 2392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 2944 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform -1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 21620 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform -1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform 1 0 20608 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform -1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 20608 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform -1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 19596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 19136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5980 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 4232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 4692 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9844 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 7912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 13248 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 12420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 18952 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 17940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1649977179
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 16008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 19872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 19688 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 9200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17204 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17572 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 3312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_40
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_127
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_139
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_151
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_95
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_78
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_90
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_102
timestamp 1649977179
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_212
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_25
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1649977179
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_136
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_203
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_222
timestamp 1649977179
transform 1 0 21528 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_40
timestamp 1649977179
transform 1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_117
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_220
timestamp 1649977179
transform 1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1649977179
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_46
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_70
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1649977179
transform 1 0 21528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_39
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_62
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_99
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_111
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1649977179
transform 1 0 21528 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_14
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1649977179
transform 1 0 21528 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_44
timestamp 1649977179
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1649977179
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_172
timestamp 1649977179
transform 1 0 16928 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_180
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_190
timestamp 1649977179
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_79
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_87
timestamp 1649977179
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_135
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_152
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_178
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1649977179
transform 1 0 21528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp 1649977179
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_150
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_188
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1649977179
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_70
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_100
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_160
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_197
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_9
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1649977179
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_101
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_127
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_164
timestamp 1649977179
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_152
timestamp 1649977179
transform 1 0 15088 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1649977179
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_53
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_91
timestamp 1649977179
transform 1 0 9476 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_155
timestamp 1649977179
transform 1 0 15364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_182
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_186
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1649977179
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_127
timestamp 1649977179
transform 1 0 12788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1649977179
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_156
timestamp 1649977179
transform 1 0 15456 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_159
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1649977179
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_204
timestamp 1649977179
transform 1 0 19872 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1649977179
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_24
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_91
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_103
timestamp 1649977179
transform 1 0 10580 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1649977179
transform 1 0 15640 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_137
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1649977179
transform 1 0 16100 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_172
timestamp 1649977179
transform 1 0 16928 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1649977179
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_214
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_35
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1649977179
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_141
timestamp 1649977179
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_154
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_178
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_194
timestamp 1649977179
transform 1 0 18952 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_216
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_12
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1649977179
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1649977179
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1649977179
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1649977179
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_193
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_199
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_211
timestamp 1649977179
transform 1 0 20516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_63
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_91
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_151
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1649977179
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_35
timestamp 1649977179
transform 1 0 4324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_87
timestamp 1649977179
transform 1 0 9108 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_113
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_137
timestamp 1649977179
transform 1 0 13708 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_159
timestamp 1649977179
transform 1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_184
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_210
timestamp 1649977179
transform 1 0 20424 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_222
timestamp 1649977179
transform 1 0 21528 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_92
timestamp 1649977179
transform 1 0 9568 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1649977179
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1649977179
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_183
timestamp 1649977179
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_197
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_213
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1649977179
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1649977179
transform 1 0 21528 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_124
timestamp 1649977179
transform 1 0 12512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_149
timestamp 1649977179
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1649977179
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1649977179
transform 1 0 13156 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_195
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1649977179
transform 1 0 21528 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1649977179
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_150
timestamp 1649977179
transform 1 0 14904 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_184
timestamp 1649977179
transform 1 0 18032 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_214
timestamp 1649977179
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1649977179
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1649977179
transform -1 0 16468 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform 1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform -1 0 18032 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform -1 0 15640 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform -1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform -1 0 18032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform -1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform -1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform -1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1649977179
transform -1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1649977179
transform -1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1649977179
transform -1 0 2576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1649977179
transform -1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1649977179
transform -1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform -1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform -1 0 1840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform -1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform -1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform 1 0 20976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform 1 0 20884 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform -1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 18400 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1649977179
transform 1 0 19320 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5612 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 4784 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10120 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4140 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6072 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4692 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6256 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5520 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12788 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12696 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9568 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10580 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4232 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8832 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8372 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3864 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6992 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4692 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5888 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12788 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9476 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12512 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8188 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4324 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3864 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3312 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3404 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5796 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5796 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5796 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform -1 0 3312 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4784 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5520 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12604 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3036 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15824 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18584 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16468 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20240 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13984 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16928 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19320 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15272 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 19412 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17204 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 20240 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18768 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform -1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17848 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18860 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19320 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 19044 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20240 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19320 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18584 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4876 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 9292 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10212 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13984 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10580 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7360 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14628 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13892 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16192 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17296 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17112 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19412 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18308 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15732 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14720 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15272 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17940 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16560 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16560 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17756 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17204 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17112 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18216 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16652 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15180 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15916 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 5612 0 -1 3264
box -38 -48 590 592
<< labels >>
flabel metal2 s 1674 22200 1730 23000 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 21178 22200 21234 23000 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 1 nsew signal tristate
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 Test_en_N_out
port 2 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 3 nsew signal input
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 ccff_head
port 6 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 ccff_tail
port 7 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 8 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 9 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 10 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 11 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 12 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 13 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 14 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 15 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 16 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 17 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 18 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 19 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 20 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 21 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 22 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 23 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 24 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 25 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 26 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 27 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 28 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 29 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 30 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 31 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 32 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 33 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 34 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 35 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 36 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 37 nsew signal tristate
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 38 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 39 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 40 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 41 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 42 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 43 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 44 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 45 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 46 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 47 nsew signal tristate
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 48 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 49 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 50 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 51 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 52 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 53 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 54 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 55 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 56 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 57 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 58 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 59 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 60 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 61 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 62 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 63 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 64 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 65 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 66 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 67 nsew signal input
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 68 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 69 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 70 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 71 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 72 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 73 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 74 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 75 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 76 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 77 nsew signal tristate
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 78 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 79 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 80 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 81 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 82 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 83 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 84 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 85 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 86 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 87 nsew signal tristate
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal2 s 10138 22200 10194 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal2 s 10506 22200 10562 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 11610 22200 11666 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal2 s 12346 22200 12402 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 12714 22200 12770 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 13450 22200 13506 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 98 nsew signal input
flabel metal2 s 6826 22200 6882 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 99 nsew signal input
flabel metal2 s 7194 22200 7250 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 100 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 101 nsew signal input
flabel metal2 s 7930 22200 7986 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 102 nsew signal input
flabel metal2 s 8298 22200 8354 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 103 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 104 nsew signal input
flabel metal2 s 9034 22200 9090 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 105 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 106 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 107 nsew signal input
flabel metal2 s 13818 22200 13874 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 108 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 109 nsew signal tristate
flabel metal2 s 17866 22200 17922 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 110 nsew signal tristate
flabel metal2 s 18234 22200 18290 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 111 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 112 nsew signal tristate
flabel metal2 s 18970 22200 19026 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 113 nsew signal tristate
flabel metal2 s 19338 22200 19394 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 114 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 115 nsew signal tristate
flabel metal2 s 20074 22200 20130 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 116 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 117 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 118 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 119 nsew signal tristate
flabel metal2 s 14554 22200 14610 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 120 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 121 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 122 nsew signal tristate
flabel metal2 s 15658 22200 15714 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 123 nsew signal tristate
flabel metal2 s 16026 22200 16082 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 124 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 125 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 126 nsew signal tristate
flabel metal2 s 17130 22200 17186 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 127 nsew signal tristate
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 clk_3_N_out
port 128 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 clk_3_S_in
port 129 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_11_
port 130 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_13_
port 131 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_15_
port 132 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 left_bottom_grid_pin_17_
port 133 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_1_
port 134 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_3_
port 135 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_5_
port 136 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_7_
port 137 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_9_
port 138 nsew signal input
flabel metal2 s 4986 22200 5042 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 139 nsew signal input
flabel metal2 s 6090 22200 6146 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 140 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 prog_clk_3_S_in
port 141 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_11_
port 142 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_13_
port 143 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_15_
port 144 nsew signal input
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 right_bottom_grid_pin_17_
port 145 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_1_
port 146 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_3_
port 147 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_5_
port 148 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_7_
port 149 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_9_
port 150 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 151 nsew signal input
flabel metal2 s 2410 22200 2466 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 152 nsew signal input
flabel metal2 s 2778 22200 2834 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 153 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 154 nsew signal input
flabel metal2 s 3514 22200 3570 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 155 nsew signal input
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 156 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 157 nsew signal input
flabel metal2 s 4618 22200 4674 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 158 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
