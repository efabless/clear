VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tile
  CLASS BLOCK ;
  FOREIGN tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 255.000 BY 285.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.720 10.640 91.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.720 10.640 141.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 10.640 191.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.720 10.640 241.320 272.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.720 10.640 16.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 10.640 116.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.720 10.640 166.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.720 10.640 216.320 272.240 ;
    END
  END VPWR
  PIN bottom_width_0_height_0_subtile_0__pin_cout_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_cout_0_
  PIN bottom_width_0_height_0_subtile_0__pin_reg_out_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_reg_out_0_
  PIN ccff_head_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END ccff_head_1
  PIN ccff_head_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 237.450 281.000 237.730 285.000 ;
    END
  END ccff_head_2
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 21.120 255.000 21.720 ;
    END
  END ccff_tail
  PIN ccff_tail_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 16.650 281.000 16.930 285.000 ;
    END
  END ccff_tail_0
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END chanx_left_in[29]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END chanx_left_out[29]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 126.520 255.000 127.120 ;
    END
  END chanx_right_in_0[0]
  PIN chanx_right_in_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 160.520 255.000 161.120 ;
    END
  END chanx_right_in_0[10]
  PIN chanx_right_in_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 163.920 255.000 164.520 ;
    END
  END chanx_right_in_0[11]
  PIN chanx_right_in_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 167.320 255.000 167.920 ;
    END
  END chanx_right_in_0[12]
  PIN chanx_right_in_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 170.720 255.000 171.320 ;
    END
  END chanx_right_in_0[13]
  PIN chanx_right_in_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 174.120 255.000 174.720 ;
    END
  END chanx_right_in_0[14]
  PIN chanx_right_in_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 177.520 255.000 178.120 ;
    END
  END chanx_right_in_0[15]
  PIN chanx_right_in_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 180.920 255.000 181.520 ;
    END
  END chanx_right_in_0[16]
  PIN chanx_right_in_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 184.320 255.000 184.920 ;
    END
  END chanx_right_in_0[17]
  PIN chanx_right_in_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 187.720 255.000 188.320 ;
    END
  END chanx_right_in_0[18]
  PIN chanx_right_in_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 191.120 255.000 191.720 ;
    END
  END chanx_right_in_0[19]
  PIN chanx_right_in_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 129.920 255.000 130.520 ;
    END
  END chanx_right_in_0[1]
  PIN chanx_right_in_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 194.520 255.000 195.120 ;
    END
  END chanx_right_in_0[20]
  PIN chanx_right_in_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 197.920 255.000 198.520 ;
    END
  END chanx_right_in_0[21]
  PIN chanx_right_in_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 201.320 255.000 201.920 ;
    END
  END chanx_right_in_0[22]
  PIN chanx_right_in_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 204.720 255.000 205.320 ;
    END
  END chanx_right_in_0[23]
  PIN chanx_right_in_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 208.120 255.000 208.720 ;
    END
  END chanx_right_in_0[24]
  PIN chanx_right_in_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 211.520 255.000 212.120 ;
    END
  END chanx_right_in_0[25]
  PIN chanx_right_in_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 214.920 255.000 215.520 ;
    END
  END chanx_right_in_0[26]
  PIN chanx_right_in_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 218.320 255.000 218.920 ;
    END
  END chanx_right_in_0[27]
  PIN chanx_right_in_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 221.720 255.000 222.320 ;
    END
  END chanx_right_in_0[28]
  PIN chanx_right_in_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 225.120 255.000 225.720 ;
    END
  END chanx_right_in_0[29]
  PIN chanx_right_in_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 133.320 255.000 133.920 ;
    END
  END chanx_right_in_0[2]
  PIN chanx_right_in_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 136.720 255.000 137.320 ;
    END
  END chanx_right_in_0[3]
  PIN chanx_right_in_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 140.120 255.000 140.720 ;
    END
  END chanx_right_in_0[4]
  PIN chanx_right_in_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 143.520 255.000 144.120 ;
    END
  END chanx_right_in_0[5]
  PIN chanx_right_in_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 146.920 255.000 147.520 ;
    END
  END chanx_right_in_0[6]
  PIN chanx_right_in_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 150.320 255.000 150.920 ;
    END
  END chanx_right_in_0[7]
  PIN chanx_right_in_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 153.720 255.000 154.320 ;
    END
  END chanx_right_in_0[8]
  PIN chanx_right_in_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 157.120 255.000 157.720 ;
    END
  END chanx_right_in_0[9]
  PIN chanx_right_out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 24.520 255.000 25.120 ;
    END
  END chanx_right_out_0[0]
  PIN chanx_right_out_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 58.520 255.000 59.120 ;
    END
  END chanx_right_out_0[10]
  PIN chanx_right_out_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 61.920 255.000 62.520 ;
    END
  END chanx_right_out_0[11]
  PIN chanx_right_out_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 65.320 255.000 65.920 ;
    END
  END chanx_right_out_0[12]
  PIN chanx_right_out_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 68.720 255.000 69.320 ;
    END
  END chanx_right_out_0[13]
  PIN chanx_right_out_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 72.120 255.000 72.720 ;
    END
  END chanx_right_out_0[14]
  PIN chanx_right_out_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 75.520 255.000 76.120 ;
    END
  END chanx_right_out_0[15]
  PIN chanx_right_out_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 78.920 255.000 79.520 ;
    END
  END chanx_right_out_0[16]
  PIN chanx_right_out_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 82.320 255.000 82.920 ;
    END
  END chanx_right_out_0[17]
  PIN chanx_right_out_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 85.720 255.000 86.320 ;
    END
  END chanx_right_out_0[18]
  PIN chanx_right_out_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 89.120 255.000 89.720 ;
    END
  END chanx_right_out_0[19]
  PIN chanx_right_out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 27.920 255.000 28.520 ;
    END
  END chanx_right_out_0[1]
  PIN chanx_right_out_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 92.520 255.000 93.120 ;
    END
  END chanx_right_out_0[20]
  PIN chanx_right_out_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 95.920 255.000 96.520 ;
    END
  END chanx_right_out_0[21]
  PIN chanx_right_out_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 99.320 255.000 99.920 ;
    END
  END chanx_right_out_0[22]
  PIN chanx_right_out_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 102.720 255.000 103.320 ;
    END
  END chanx_right_out_0[23]
  PIN chanx_right_out_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 106.120 255.000 106.720 ;
    END
  END chanx_right_out_0[24]
  PIN chanx_right_out_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 109.520 255.000 110.120 ;
    END
  END chanx_right_out_0[25]
  PIN chanx_right_out_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 112.920 255.000 113.520 ;
    END
  END chanx_right_out_0[26]
  PIN chanx_right_out_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 116.320 255.000 116.920 ;
    END
  END chanx_right_out_0[27]
  PIN chanx_right_out_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 119.720 255.000 120.320 ;
    END
  END chanx_right_out_0[28]
  PIN chanx_right_out_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 123.120 255.000 123.720 ;
    END
  END chanx_right_out_0[29]
  PIN chanx_right_out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 31.320 255.000 31.920 ;
    END
  END chanx_right_out_0[2]
  PIN chanx_right_out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 34.720 255.000 35.320 ;
    END
  END chanx_right_out_0[3]
  PIN chanx_right_out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 38.120 255.000 38.720 ;
    END
  END chanx_right_out_0[4]
  PIN chanx_right_out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 41.520 255.000 42.120 ;
    END
  END chanx_right_out_0[5]
  PIN chanx_right_out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 44.920 255.000 45.520 ;
    END
  END chanx_right_out_0[6]
  PIN chanx_right_out_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 48.320 255.000 48.920 ;
    END
  END chanx_right_out_0[7]
  PIN chanx_right_out_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 51.720 255.000 52.320 ;
    END
  END chanx_right_out_0[8]
  PIN chanx_right_out_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 55.120 255.000 55.720 ;
    END
  END chanx_right_out_0[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END chany_bottom_in[29]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END chany_bottom_out[29]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 281.000 102.490 285.000 ;
    END
  END chany_top_in_0[0]
  PIN chany_top_in_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 281.000 130.090 285.000 ;
    END
  END chany_top_in_0[10]
  PIN chany_top_in_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 132.570 281.000 132.850 285.000 ;
    END
  END chany_top_in_0[11]
  PIN chany_top_in_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 281.000 135.610 285.000 ;
    END
  END chany_top_in_0[12]
  PIN chany_top_in_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 281.000 138.370 285.000 ;
    END
  END chany_top_in_0[13]
  PIN chany_top_in_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 281.000 141.130 285.000 ;
    END
  END chany_top_in_0[14]
  PIN chany_top_in_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 143.610 281.000 143.890 285.000 ;
    END
  END chany_top_in_0[15]
  PIN chany_top_in_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 146.370 281.000 146.650 285.000 ;
    END
  END chany_top_in_0[16]
  PIN chany_top_in_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 149.130 281.000 149.410 285.000 ;
    END
  END chany_top_in_0[17]
  PIN chany_top_in_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 281.000 152.170 285.000 ;
    END
  END chany_top_in_0[18]
  PIN chany_top_in_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 281.000 154.930 285.000 ;
    END
  END chany_top_in_0[19]
  PIN chany_top_in_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 104.970 281.000 105.250 285.000 ;
    END
  END chany_top_in_0[1]
  PIN chany_top_in_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 281.000 157.690 285.000 ;
    END
  END chany_top_in_0[20]
  PIN chany_top_in_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 160.170 281.000 160.450 285.000 ;
    END
  END chany_top_in_0[21]
  PIN chany_top_in_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 162.930 281.000 163.210 285.000 ;
    END
  END chany_top_in_0[22]
  PIN chany_top_in_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 165.690 281.000 165.970 285.000 ;
    END
  END chany_top_in_0[23]
  PIN chany_top_in_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 281.000 168.730 285.000 ;
    END
  END chany_top_in_0[24]
  PIN chany_top_in_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 281.000 171.490 285.000 ;
    END
  END chany_top_in_0[25]
  PIN chany_top_in_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 281.000 174.250 285.000 ;
    END
  END chany_top_in_0[26]
  PIN chany_top_in_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 176.730 281.000 177.010 285.000 ;
    END
  END chany_top_in_0[27]
  PIN chany_top_in_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 179.490 281.000 179.770 285.000 ;
    END
  END chany_top_in_0[28]
  PIN chany_top_in_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 182.250 281.000 182.530 285.000 ;
    END
  END chany_top_in_0[29]
  PIN chany_top_in_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 281.000 108.010 285.000 ;
    END
  END chany_top_in_0[2]
  PIN chany_top_in_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 281.000 110.770 285.000 ;
    END
  END chany_top_in_0[3]
  PIN chany_top_in_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 113.250 281.000 113.530 285.000 ;
    END
  END chany_top_in_0[4]
  PIN chany_top_in_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 281.000 116.290 285.000 ;
    END
  END chany_top_in_0[5]
  PIN chany_top_in_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 281.000 119.050 285.000 ;
    END
  END chany_top_in_0[6]
  PIN chany_top_in_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 281.000 121.810 285.000 ;
    END
  END chany_top_in_0[7]
  PIN chany_top_in_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 124.290 281.000 124.570 285.000 ;
    END
  END chany_top_in_0[8]
  PIN chany_top_in_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 127.050 281.000 127.330 285.000 ;
    END
  END chany_top_in_0[9]
  PIN chany_top_out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 19.410 281.000 19.690 285.000 ;
    END
  END chany_top_out_0[0]
  PIN chany_top_out_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 47.010 281.000 47.290 285.000 ;
    END
  END chany_top_out_0[10]
  PIN chany_top_out_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 49.770 281.000 50.050 285.000 ;
    END
  END chany_top_out_0[11]
  PIN chany_top_out_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 52.530 281.000 52.810 285.000 ;
    END
  END chany_top_out_0[12]
  PIN chany_top_out_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 55.290 281.000 55.570 285.000 ;
    END
  END chany_top_out_0[13]
  PIN chany_top_out_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 281.000 58.330 285.000 ;
    END
  END chany_top_out_0[14]
  PIN chany_top_out_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 60.810 281.000 61.090 285.000 ;
    END
  END chany_top_out_0[15]
  PIN chany_top_out_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 63.570 281.000 63.850 285.000 ;
    END
  END chany_top_out_0[16]
  PIN chany_top_out_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 66.330 281.000 66.610 285.000 ;
    END
  END chany_top_out_0[17]
  PIN chany_top_out_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 69.090 281.000 69.370 285.000 ;
    END
  END chany_top_out_0[18]
  PIN chany_top_out_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 71.850 281.000 72.130 285.000 ;
    END
  END chany_top_out_0[19]
  PIN chany_top_out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 22.170 281.000 22.450 285.000 ;
    END
  END chany_top_out_0[1]
  PIN chany_top_out_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 74.610 281.000 74.890 285.000 ;
    END
  END chany_top_out_0[20]
  PIN chany_top_out_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 77.370 281.000 77.650 285.000 ;
    END
  END chany_top_out_0[21]
  PIN chany_top_out_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 80.130 281.000 80.410 285.000 ;
    END
  END chany_top_out_0[22]
  PIN chany_top_out_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 82.890 281.000 83.170 285.000 ;
    END
  END chany_top_out_0[23]
  PIN chany_top_out_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 85.650 281.000 85.930 285.000 ;
    END
  END chany_top_out_0[24]
  PIN chany_top_out_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 88.410 281.000 88.690 285.000 ;
    END
  END chany_top_out_0[25]
  PIN chany_top_out_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 91.170 281.000 91.450 285.000 ;
    END
  END chany_top_out_0[26]
  PIN chany_top_out_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 93.930 281.000 94.210 285.000 ;
    END
  END chany_top_out_0[27]
  PIN chany_top_out_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 96.690 281.000 96.970 285.000 ;
    END
  END chany_top_out_0[28]
  PIN chany_top_out_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 99.450 281.000 99.730 285.000 ;
    END
  END chany_top_out_0[29]
  PIN chany_top_out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 24.930 281.000 25.210 285.000 ;
    END
  END chany_top_out_0[2]
  PIN chany_top_out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 27.690 281.000 27.970 285.000 ;
    END
  END chany_top_out_0[3]
  PIN chany_top_out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 30.450 281.000 30.730 285.000 ;
    END
  END chany_top_out_0[4]
  PIN chany_top_out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 33.210 281.000 33.490 285.000 ;
    END
  END chany_top_out_0[5]
  PIN chany_top_out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 35.970 281.000 36.250 285.000 ;
    END
  END chany_top_out_0[6]
  PIN chany_top_out_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 38.730 281.000 39.010 285.000 ;
    END
  END chany_top_out_0[7]
  PIN chany_top_out_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 41.490 281.000 41.770 285.000 ;
    END
  END chany_top_out_0[8]
  PIN chany_top_out_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 44.250 281.000 44.530 285.000 ;
    END
  END chany_top_out_0[9]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END clk0
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END prog_clk
  PIN prog_reset_bottom_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END prog_reset_bottom_in
  PIN prog_reset_bottom_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END prog_reset_bottom_out
  PIN prog_reset_left_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END prog_reset_left_in
  PIN prog_reset_right_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 228.520 255.000 229.120 ;
    END
  END prog_reset_right_out
  PIN prog_reset_top_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 281.000 193.570 285.000 ;
    END
  END prog_reset_top_in
  PIN prog_reset_top_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 190.530 281.000 190.810 285.000 ;
    END
  END prog_reset_top_out
  PIN reset_bottom_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END reset_bottom_in
  PIN reset_bottom_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END reset_bottom_out
  PIN reset_left_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END reset_left_out
  PIN reset_right_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 231.920 255.000 232.520 ;
    END
  END reset_right_in
  PIN reset_top_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 198.810 281.000 199.090 285.000 ;
    END
  END reset_top_in
  PIN reset_top_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 196.050 281.000 196.330 285.000 ;
    END
  END reset_top_out
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 235.320 255.000 235.920 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 238.720 255.000 239.320 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 242.120 255.000 242.720 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 245.520 255.000 246.120 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 248.920 255.000 249.520 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 252.320 255.000 252.920 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 255.720 255.000 256.320 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 259.120 255.000 259.720 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN right_width_0_height_0_subtile_0__pin_O_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_10_
  PIN right_width_0_height_0_subtile_0__pin_O_11_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_11_
  PIN right_width_0_height_0_subtile_0__pin_O_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_12_
  PIN right_width_0_height_0_subtile_0__pin_O_13_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_13_
  PIN right_width_0_height_0_subtile_0__pin_O_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_14_
  PIN right_width_0_height_0_subtile_0__pin_O_15_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_15_
  PIN right_width_0_height_0_subtile_0__pin_O_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_8_
  PIN right_width_0_height_0_subtile_0__pin_O_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_9_
  PIN sc_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 234.690 281.000 234.970 285.000 ;
    END
  END sc_in
  PIN sc_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END sc_out
  PIN test_enable_bottom_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END test_enable_bottom_in
  PIN test_enable_bottom_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END test_enable_bottom_out
  PIN test_enable_left_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END test_enable_left_out
  PIN test_enable_right_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 262.520 255.000 263.120 ;
    END
  END test_enable_right_in
  PIN test_enable_top_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 204.330 281.000 204.610 285.000 ;
    END
  END test_enable_top_in
  PIN test_enable_top_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 201.570 281.000 201.850 285.000 ;
    END
  END test_enable_top_out
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 281.000 212.890 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 215.370 281.000 215.650 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 218.130 281.000 218.410 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 220.890 281.000 221.170 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 223.650 281.000 223.930 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 226.410 281.000 226.690 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 281.000 207.370 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 281.000 210.130 285.000 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
  PIN top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_0_
  PIN top_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_1_
  PIN top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_2_
  PIN top_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_3_
  PIN top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_4_
  PIN top_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_5_
  PIN top_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_6_
  PIN top_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_7_
  PIN top_width_0_height_0_subtile_0__pin_cin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 281.000 229.450 285.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_cin_0_
  PIN top_width_0_height_0_subtile_0__pin_reg_in_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 281.000 232.210 285.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_reg_in_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 249.320 272.085 ;
      LAYER met1 ;
        RECT 5.520 8.540 249.320 273.320 ;
      LAYER met2 ;
        RECT 5.610 280.720 16.370 281.250 ;
        RECT 17.210 280.720 19.130 281.250 ;
        RECT 19.970 280.720 21.890 281.250 ;
        RECT 22.730 280.720 24.650 281.250 ;
        RECT 25.490 280.720 27.410 281.250 ;
        RECT 28.250 280.720 30.170 281.250 ;
        RECT 31.010 280.720 32.930 281.250 ;
        RECT 33.770 280.720 35.690 281.250 ;
        RECT 36.530 280.720 38.450 281.250 ;
        RECT 39.290 280.720 41.210 281.250 ;
        RECT 42.050 280.720 43.970 281.250 ;
        RECT 44.810 280.720 46.730 281.250 ;
        RECT 47.570 280.720 49.490 281.250 ;
        RECT 50.330 280.720 52.250 281.250 ;
        RECT 53.090 280.720 55.010 281.250 ;
        RECT 55.850 280.720 57.770 281.250 ;
        RECT 58.610 280.720 60.530 281.250 ;
        RECT 61.370 280.720 63.290 281.250 ;
        RECT 64.130 280.720 66.050 281.250 ;
        RECT 66.890 280.720 68.810 281.250 ;
        RECT 69.650 280.720 71.570 281.250 ;
        RECT 72.410 280.720 74.330 281.250 ;
        RECT 75.170 280.720 77.090 281.250 ;
        RECT 77.930 280.720 79.850 281.250 ;
        RECT 80.690 280.720 82.610 281.250 ;
        RECT 83.450 280.720 85.370 281.250 ;
        RECT 86.210 280.720 88.130 281.250 ;
        RECT 88.970 280.720 90.890 281.250 ;
        RECT 91.730 280.720 93.650 281.250 ;
        RECT 94.490 280.720 96.410 281.250 ;
        RECT 97.250 280.720 99.170 281.250 ;
        RECT 100.010 280.720 101.930 281.250 ;
        RECT 102.770 280.720 104.690 281.250 ;
        RECT 105.530 280.720 107.450 281.250 ;
        RECT 108.290 280.720 110.210 281.250 ;
        RECT 111.050 280.720 112.970 281.250 ;
        RECT 113.810 280.720 115.730 281.250 ;
        RECT 116.570 280.720 118.490 281.250 ;
        RECT 119.330 280.720 121.250 281.250 ;
        RECT 122.090 280.720 124.010 281.250 ;
        RECT 124.850 280.720 126.770 281.250 ;
        RECT 127.610 280.720 129.530 281.250 ;
        RECT 130.370 280.720 132.290 281.250 ;
        RECT 133.130 280.720 135.050 281.250 ;
        RECT 135.890 280.720 137.810 281.250 ;
        RECT 138.650 280.720 140.570 281.250 ;
        RECT 141.410 280.720 143.330 281.250 ;
        RECT 144.170 280.720 146.090 281.250 ;
        RECT 146.930 280.720 148.850 281.250 ;
        RECT 149.690 280.720 151.610 281.250 ;
        RECT 152.450 280.720 154.370 281.250 ;
        RECT 155.210 280.720 157.130 281.250 ;
        RECT 157.970 280.720 159.890 281.250 ;
        RECT 160.730 280.720 162.650 281.250 ;
        RECT 163.490 280.720 165.410 281.250 ;
        RECT 166.250 280.720 168.170 281.250 ;
        RECT 169.010 280.720 170.930 281.250 ;
        RECT 171.770 280.720 173.690 281.250 ;
        RECT 174.530 280.720 176.450 281.250 ;
        RECT 177.290 280.720 179.210 281.250 ;
        RECT 180.050 280.720 181.970 281.250 ;
        RECT 182.810 280.720 190.250 281.250 ;
        RECT 191.090 280.720 193.010 281.250 ;
        RECT 193.850 280.720 195.770 281.250 ;
        RECT 196.610 280.720 198.530 281.250 ;
        RECT 199.370 280.720 201.290 281.250 ;
        RECT 202.130 280.720 204.050 281.250 ;
        RECT 204.890 280.720 206.810 281.250 ;
        RECT 207.650 280.720 209.570 281.250 ;
        RECT 210.410 280.720 212.330 281.250 ;
        RECT 213.170 280.720 215.090 281.250 ;
        RECT 215.930 280.720 217.850 281.250 ;
        RECT 218.690 280.720 220.610 281.250 ;
        RECT 221.450 280.720 223.370 281.250 ;
        RECT 224.210 280.720 226.130 281.250 ;
        RECT 226.970 280.720 228.890 281.250 ;
        RECT 229.730 280.720 231.650 281.250 ;
        RECT 232.490 280.720 234.410 281.250 ;
        RECT 235.250 280.720 237.170 281.250 ;
        RECT 238.010 280.720 248.310 281.250 ;
        RECT 5.610 4.280 248.310 280.720 ;
        RECT 5.610 3.670 16.370 4.280 ;
        RECT 17.210 3.670 19.130 4.280 ;
        RECT 19.970 3.670 21.890 4.280 ;
        RECT 22.730 3.670 24.650 4.280 ;
        RECT 25.490 3.670 27.410 4.280 ;
        RECT 28.250 3.670 30.170 4.280 ;
        RECT 31.010 3.670 32.930 4.280 ;
        RECT 33.770 3.670 35.690 4.280 ;
        RECT 36.530 3.670 38.450 4.280 ;
        RECT 39.290 3.670 41.210 4.280 ;
        RECT 42.050 3.670 43.970 4.280 ;
        RECT 44.810 3.670 46.730 4.280 ;
        RECT 47.570 3.670 49.490 4.280 ;
        RECT 50.330 3.670 52.250 4.280 ;
        RECT 53.090 3.670 55.010 4.280 ;
        RECT 55.850 3.670 57.770 4.280 ;
        RECT 58.610 3.670 60.530 4.280 ;
        RECT 61.370 3.670 63.290 4.280 ;
        RECT 64.130 3.670 66.050 4.280 ;
        RECT 66.890 3.670 68.810 4.280 ;
        RECT 69.650 3.670 71.570 4.280 ;
        RECT 72.410 3.670 74.330 4.280 ;
        RECT 75.170 3.670 77.090 4.280 ;
        RECT 77.930 3.670 79.850 4.280 ;
        RECT 80.690 3.670 82.610 4.280 ;
        RECT 83.450 3.670 85.370 4.280 ;
        RECT 86.210 3.670 88.130 4.280 ;
        RECT 88.970 3.670 90.890 4.280 ;
        RECT 91.730 3.670 93.650 4.280 ;
        RECT 94.490 3.670 96.410 4.280 ;
        RECT 97.250 3.670 99.170 4.280 ;
        RECT 100.010 3.670 101.930 4.280 ;
        RECT 102.770 3.670 104.690 4.280 ;
        RECT 105.530 3.670 107.450 4.280 ;
        RECT 108.290 3.670 110.210 4.280 ;
        RECT 111.050 3.670 112.970 4.280 ;
        RECT 113.810 3.670 115.730 4.280 ;
        RECT 116.570 3.670 118.490 4.280 ;
        RECT 119.330 3.670 121.250 4.280 ;
        RECT 122.090 3.670 124.010 4.280 ;
        RECT 124.850 3.670 126.770 4.280 ;
        RECT 127.610 3.670 129.530 4.280 ;
        RECT 130.370 3.670 132.290 4.280 ;
        RECT 133.130 3.670 135.050 4.280 ;
        RECT 135.890 3.670 137.810 4.280 ;
        RECT 138.650 3.670 140.570 4.280 ;
        RECT 141.410 3.670 143.330 4.280 ;
        RECT 144.170 3.670 146.090 4.280 ;
        RECT 146.930 3.670 148.850 4.280 ;
        RECT 149.690 3.670 151.610 4.280 ;
        RECT 152.450 3.670 154.370 4.280 ;
        RECT 155.210 3.670 157.130 4.280 ;
        RECT 157.970 3.670 159.890 4.280 ;
        RECT 160.730 3.670 162.650 4.280 ;
        RECT 163.490 3.670 165.410 4.280 ;
        RECT 166.250 3.670 168.170 4.280 ;
        RECT 169.010 3.670 170.930 4.280 ;
        RECT 171.770 3.670 173.690 4.280 ;
        RECT 174.530 3.670 176.450 4.280 ;
        RECT 177.290 3.670 179.210 4.280 ;
        RECT 180.050 3.670 181.970 4.280 ;
        RECT 182.810 3.670 184.730 4.280 ;
        RECT 185.570 3.670 187.490 4.280 ;
        RECT 188.330 3.670 190.250 4.280 ;
        RECT 191.090 3.670 193.010 4.280 ;
        RECT 193.850 3.670 195.770 4.280 ;
        RECT 196.610 3.670 198.530 4.280 ;
        RECT 199.370 3.670 201.290 4.280 ;
        RECT 202.130 3.670 204.050 4.280 ;
        RECT 204.890 3.670 206.810 4.280 ;
        RECT 207.650 3.670 209.570 4.280 ;
        RECT 210.410 3.670 212.330 4.280 ;
        RECT 213.170 3.670 215.090 4.280 ;
        RECT 215.930 3.670 217.850 4.280 ;
        RECT 218.690 3.670 220.610 4.280 ;
        RECT 221.450 3.670 223.370 4.280 ;
        RECT 224.210 3.670 226.130 4.280 ;
        RECT 226.970 3.670 228.890 4.280 ;
        RECT 229.730 3.670 231.650 4.280 ;
        RECT 232.490 3.670 234.410 4.280 ;
        RECT 235.250 3.670 248.310 4.280 ;
      LAYER met3 ;
        RECT 4.000 263.520 251.000 272.165 ;
        RECT 4.400 262.120 250.600 263.520 ;
        RECT 4.000 260.120 251.000 262.120 ;
        RECT 4.400 258.720 250.600 260.120 ;
        RECT 4.000 256.720 251.000 258.720 ;
        RECT 4.400 255.320 250.600 256.720 ;
        RECT 4.000 253.320 251.000 255.320 ;
        RECT 4.400 251.920 250.600 253.320 ;
        RECT 4.000 249.920 251.000 251.920 ;
        RECT 4.400 248.520 250.600 249.920 ;
        RECT 4.000 246.520 251.000 248.520 ;
        RECT 4.400 245.120 250.600 246.520 ;
        RECT 4.000 243.120 251.000 245.120 ;
        RECT 4.400 241.720 250.600 243.120 ;
        RECT 4.000 239.720 251.000 241.720 ;
        RECT 4.400 238.320 250.600 239.720 ;
        RECT 4.000 236.320 251.000 238.320 ;
        RECT 4.400 234.920 250.600 236.320 ;
        RECT 4.000 232.920 251.000 234.920 ;
        RECT 4.400 231.520 250.600 232.920 ;
        RECT 4.000 229.520 251.000 231.520 ;
        RECT 4.400 228.120 250.600 229.520 ;
        RECT 4.000 226.120 251.000 228.120 ;
        RECT 4.400 224.720 250.600 226.120 ;
        RECT 4.000 222.720 251.000 224.720 ;
        RECT 4.400 221.320 250.600 222.720 ;
        RECT 4.000 219.320 251.000 221.320 ;
        RECT 4.400 217.920 250.600 219.320 ;
        RECT 4.000 215.920 251.000 217.920 ;
        RECT 4.400 214.520 250.600 215.920 ;
        RECT 4.000 212.520 251.000 214.520 ;
        RECT 4.400 211.120 250.600 212.520 ;
        RECT 4.000 209.120 251.000 211.120 ;
        RECT 4.400 207.720 250.600 209.120 ;
        RECT 4.000 205.720 251.000 207.720 ;
        RECT 4.400 204.320 250.600 205.720 ;
        RECT 4.000 202.320 251.000 204.320 ;
        RECT 4.400 200.920 250.600 202.320 ;
        RECT 4.000 198.920 251.000 200.920 ;
        RECT 4.400 197.520 250.600 198.920 ;
        RECT 4.000 195.520 251.000 197.520 ;
        RECT 4.400 194.120 250.600 195.520 ;
        RECT 4.000 192.120 251.000 194.120 ;
        RECT 4.400 190.720 250.600 192.120 ;
        RECT 4.000 188.720 251.000 190.720 ;
        RECT 4.400 187.320 250.600 188.720 ;
        RECT 4.000 185.320 251.000 187.320 ;
        RECT 4.400 183.920 250.600 185.320 ;
        RECT 4.000 181.920 251.000 183.920 ;
        RECT 4.400 180.520 250.600 181.920 ;
        RECT 4.000 178.520 251.000 180.520 ;
        RECT 4.400 177.120 250.600 178.520 ;
        RECT 4.000 175.120 251.000 177.120 ;
        RECT 4.400 173.720 250.600 175.120 ;
        RECT 4.000 171.720 251.000 173.720 ;
        RECT 4.400 170.320 250.600 171.720 ;
        RECT 4.000 168.320 251.000 170.320 ;
        RECT 4.400 166.920 250.600 168.320 ;
        RECT 4.000 164.920 251.000 166.920 ;
        RECT 4.400 163.520 250.600 164.920 ;
        RECT 4.000 161.520 251.000 163.520 ;
        RECT 4.400 160.120 250.600 161.520 ;
        RECT 4.000 158.120 251.000 160.120 ;
        RECT 4.400 156.720 250.600 158.120 ;
        RECT 4.000 154.720 251.000 156.720 ;
        RECT 4.400 153.320 250.600 154.720 ;
        RECT 4.000 151.320 251.000 153.320 ;
        RECT 4.400 149.920 250.600 151.320 ;
        RECT 4.000 147.920 251.000 149.920 ;
        RECT 4.400 146.520 250.600 147.920 ;
        RECT 4.000 144.520 251.000 146.520 ;
        RECT 4.400 143.120 250.600 144.520 ;
        RECT 4.000 141.120 251.000 143.120 ;
        RECT 4.400 139.720 250.600 141.120 ;
        RECT 4.000 137.720 251.000 139.720 ;
        RECT 4.400 136.320 250.600 137.720 ;
        RECT 4.000 134.320 251.000 136.320 ;
        RECT 4.400 132.920 250.600 134.320 ;
        RECT 4.000 130.920 251.000 132.920 ;
        RECT 4.400 129.520 250.600 130.920 ;
        RECT 4.000 127.520 251.000 129.520 ;
        RECT 4.400 126.120 250.600 127.520 ;
        RECT 4.000 124.120 251.000 126.120 ;
        RECT 4.400 122.720 250.600 124.120 ;
        RECT 4.000 120.720 251.000 122.720 ;
        RECT 4.400 119.320 250.600 120.720 ;
        RECT 4.000 117.320 251.000 119.320 ;
        RECT 4.400 115.920 250.600 117.320 ;
        RECT 4.000 113.920 251.000 115.920 ;
        RECT 4.400 112.520 250.600 113.920 ;
        RECT 4.000 110.520 251.000 112.520 ;
        RECT 4.400 109.120 250.600 110.520 ;
        RECT 4.000 107.120 251.000 109.120 ;
        RECT 4.400 105.720 250.600 107.120 ;
        RECT 4.000 103.720 251.000 105.720 ;
        RECT 4.400 102.320 250.600 103.720 ;
        RECT 4.000 100.320 251.000 102.320 ;
        RECT 4.400 98.920 250.600 100.320 ;
        RECT 4.000 96.920 251.000 98.920 ;
        RECT 4.400 95.520 250.600 96.920 ;
        RECT 4.000 93.520 251.000 95.520 ;
        RECT 4.400 92.120 250.600 93.520 ;
        RECT 4.000 90.120 251.000 92.120 ;
        RECT 4.400 88.720 250.600 90.120 ;
        RECT 4.000 86.720 251.000 88.720 ;
        RECT 4.400 85.320 250.600 86.720 ;
        RECT 4.000 83.320 251.000 85.320 ;
        RECT 4.400 81.920 250.600 83.320 ;
        RECT 4.000 79.920 251.000 81.920 ;
        RECT 4.400 78.520 250.600 79.920 ;
        RECT 4.000 76.520 251.000 78.520 ;
        RECT 4.400 75.120 250.600 76.520 ;
        RECT 4.000 73.120 251.000 75.120 ;
        RECT 4.400 71.720 250.600 73.120 ;
        RECT 4.000 69.720 251.000 71.720 ;
        RECT 4.400 68.320 250.600 69.720 ;
        RECT 4.000 66.320 251.000 68.320 ;
        RECT 4.400 64.920 250.600 66.320 ;
        RECT 4.000 62.920 251.000 64.920 ;
        RECT 4.400 61.520 250.600 62.920 ;
        RECT 4.000 59.520 251.000 61.520 ;
        RECT 4.400 58.120 250.600 59.520 ;
        RECT 4.000 56.120 251.000 58.120 ;
        RECT 4.400 54.720 250.600 56.120 ;
        RECT 4.000 52.720 251.000 54.720 ;
        RECT 4.400 51.320 250.600 52.720 ;
        RECT 4.000 49.320 251.000 51.320 ;
        RECT 4.400 47.920 250.600 49.320 ;
        RECT 4.000 45.920 251.000 47.920 ;
        RECT 4.400 44.520 250.600 45.920 ;
        RECT 4.000 42.520 251.000 44.520 ;
        RECT 4.400 41.120 250.600 42.520 ;
        RECT 4.000 39.120 251.000 41.120 ;
        RECT 4.400 37.720 250.600 39.120 ;
        RECT 4.000 35.720 251.000 37.720 ;
        RECT 4.400 34.320 250.600 35.720 ;
        RECT 4.000 32.320 251.000 34.320 ;
        RECT 4.400 30.920 250.600 32.320 ;
        RECT 4.000 28.920 251.000 30.920 ;
        RECT 4.400 27.520 250.600 28.920 ;
        RECT 4.000 25.520 251.000 27.520 ;
        RECT 4.400 24.120 250.600 25.520 ;
        RECT 4.000 22.120 251.000 24.120 ;
        RECT 4.000 20.720 250.600 22.120 ;
        RECT 4.000 10.715 251.000 20.720 ;
      LAYER met4 ;
        RECT 50.895 19.895 64.320 269.785 ;
        RECT 66.720 19.895 89.320 269.785 ;
        RECT 91.720 19.895 114.320 269.785 ;
        RECT 116.720 19.895 139.320 269.785 ;
        RECT 141.720 19.895 164.320 269.785 ;
        RECT 166.720 19.895 189.320 269.785 ;
        RECT 191.720 19.895 214.320 269.785 ;
        RECT 216.720 19.895 221.425 269.785 ;
  END
END tile
END LIBRARY

