magic
tech sky130A
magscale 1 2
timestamp 1625785369
<< locali >>
rect 3709 17731 3743 17833
rect 8309 12223 8343 12325
rect 10333 9911 10367 10081
rect 6929 8823 6963 8925
rect 8493 8279 8527 8381
rect 5273 7735 5307 7905
rect 6469 7259 6503 7497
rect 12909 6647 12943 6817
rect 2973 6171 3007 6341
rect 12449 4471 12483 4573
rect 8125 3927 8159 4097
rect 8953 3383 8987 3485
rect 2973 2839 3007 3077
rect 3065 2907 3099 3145
rect 5181 2975 5215 3077
rect 8585 2839 8619 3077
rect 12357 2431 12391 2601
rect 13921 1887 13955 1989
<< viali >>
rect 2697 20485 2731 20519
rect 3249 20485 3283 20519
rect 4077 20485 4111 20519
rect 1685 20349 1719 20383
rect 1869 20349 1903 20383
rect 2145 20281 2179 20315
rect 2329 20281 2363 20315
rect 2881 20281 2915 20315
rect 3433 20281 3467 20315
rect 4261 20281 4295 20315
rect 2237 20009 2271 20043
rect 2881 20009 2915 20043
rect 3157 20009 3191 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 2697 19873 2731 19907
rect 1593 19805 1627 19839
rect 2329 19465 2363 19499
rect 2605 19465 2639 19499
rect 3249 19465 3283 19499
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 2789 19261 2823 19295
rect 3065 19261 3099 19295
rect 3709 19261 3743 19295
rect 1777 19193 1811 19227
rect 3525 19125 3559 19159
rect 2145 18921 2179 18955
rect 2605 18921 2639 18955
rect 3065 18921 3099 18955
rect 4537 18921 4571 18955
rect 10609 18921 10643 18955
rect 1593 18853 1627 18887
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2789 18785 2823 18819
rect 3249 18785 3283 18819
rect 4261 18785 4295 18819
rect 4721 18785 4755 18819
rect 10793 18785 10827 18819
rect 4077 18649 4111 18683
rect 2237 18377 2271 18411
rect 3157 18377 3191 18411
rect 9597 18377 9631 18411
rect 2697 18309 2731 18343
rect 10241 18241 10275 18275
rect 2881 18173 2915 18207
rect 3341 18173 3375 18207
rect 1777 18105 1811 18139
rect 2329 18105 2363 18139
rect 9965 18105 9999 18139
rect 1685 18037 1719 18071
rect 6101 18037 6135 18071
rect 10057 18037 10091 18071
rect 2145 17833 2179 17867
rect 2789 17833 2823 17867
rect 3065 17833 3099 17867
rect 3709 17833 3743 17867
rect 7297 17833 7331 17867
rect 7941 17833 7975 17867
rect 10977 17833 11011 17867
rect 11253 17833 11287 17867
rect 9842 17765 9876 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2605 17697 2639 17731
rect 3249 17697 3283 17731
rect 3709 17697 3743 17731
rect 5540 17697 5574 17731
rect 8309 17697 8343 17731
rect 9597 17697 9631 17731
rect 11437 17697 11471 17731
rect 5273 17629 5307 17663
rect 7389 17629 7423 17663
rect 7481 17629 7515 17663
rect 8401 17629 8435 17663
rect 8585 17629 8619 17663
rect 6929 17561 6963 17595
rect 1685 17493 1719 17527
rect 6653 17493 6687 17527
rect 2145 17289 2179 17323
rect 2605 17289 2639 17323
rect 5733 17289 5767 17323
rect 7389 17289 7423 17323
rect 11897 17289 11931 17323
rect 3525 17221 3559 17255
rect 6745 17153 6779 17187
rect 11069 17153 11103 17187
rect 12541 17153 12575 17187
rect 21373 17153 21407 17187
rect 2329 17085 2363 17119
rect 2789 17085 2823 17119
rect 3249 17085 3283 17119
rect 3709 17085 3743 17119
rect 4353 17085 4387 17119
rect 9137 17085 9171 17119
rect 9413 17085 9447 17119
rect 9669 17085 9703 17119
rect 21189 17085 21223 17119
rect 1593 17017 1627 17051
rect 1777 17017 1811 17051
rect 4598 17017 4632 17051
rect 6929 17017 6963 17051
rect 8892 17017 8926 17051
rect 12265 17017 12299 17051
rect 3065 16949 3099 16983
rect 6101 16949 6135 16983
rect 7021 16949 7055 16983
rect 7757 16949 7791 16983
rect 10793 16949 10827 16983
rect 12357 16949 12391 16983
rect 2329 16745 2363 16779
rect 2789 16745 2823 16779
rect 4077 16745 4111 16779
rect 8401 16745 8435 16779
rect 10333 16745 10367 16779
rect 13645 16745 13679 16779
rect 3157 16677 3191 16711
rect 6276 16677 6310 16711
rect 9873 16677 9907 16711
rect 10876 16677 10910 16711
rect 1593 16609 1627 16643
rect 1777 16609 1811 16643
rect 2513 16609 2547 16643
rect 3249 16609 3283 16643
rect 5190 16609 5224 16643
rect 5457 16609 5491 16643
rect 6009 16609 6043 16643
rect 9229 16609 9263 16643
rect 9965 16609 9999 16643
rect 12521 16609 12555 16643
rect 3433 16541 3467 16575
rect 9781 16541 9815 16575
rect 10609 16541 10643 16575
rect 12265 16541 12299 16575
rect 7389 16405 7423 16439
rect 11989 16405 12023 16439
rect 2145 16201 2179 16235
rect 4353 16201 4387 16235
rect 5089 16201 5123 16235
rect 8401 16201 8435 16235
rect 1593 16133 1627 16167
rect 6653 16133 6687 16167
rect 4629 16065 4663 16099
rect 7205 16065 7239 16099
rect 8953 16065 8987 16099
rect 12081 16065 12115 16099
rect 2329 15997 2363 16031
rect 2973 15997 3007 16031
rect 5273 15997 5307 16031
rect 1777 15929 1811 15963
rect 3240 15929 3274 15963
rect 5549 15929 5583 15963
rect 7021 15929 7055 15963
rect 7665 15929 7699 15963
rect 2697 15861 2731 15895
rect 7113 15861 7147 15895
rect 8769 15861 8803 15895
rect 8861 15861 8895 15895
rect 2145 15657 2179 15691
rect 2605 15657 2639 15691
rect 3065 15657 3099 15691
rect 4169 15657 4203 15691
rect 4537 15657 4571 15691
rect 6193 15657 6227 15691
rect 8309 15657 8343 15691
rect 9321 15657 9355 15691
rect 12173 15657 12207 15691
rect 1593 15589 1627 15623
rect 5549 15589 5583 15623
rect 7674 15589 7708 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 2789 15521 2823 15555
rect 3249 15521 3283 15555
rect 5641 15521 5675 15555
rect 10434 15521 10468 15555
rect 10701 15521 10735 15555
rect 11805 15521 11839 15555
rect 4629 15453 4663 15487
rect 4721 15453 4755 15487
rect 5825 15453 5859 15487
rect 7941 15453 7975 15487
rect 11621 15453 11655 15487
rect 11713 15453 11747 15487
rect 5181 15317 5215 15351
rect 6561 15317 6595 15351
rect 11069 15317 11103 15351
rect 1685 15113 1719 15147
rect 2145 15113 2179 15147
rect 2881 15113 2915 15147
rect 7205 15113 7239 15147
rect 8769 15113 8803 15147
rect 4721 15045 4755 15079
rect 3479 14977 3513 15011
rect 6101 14977 6135 15011
rect 7757 14977 7791 15011
rect 9413 14977 9447 15011
rect 10425 14977 10459 15011
rect 2329 14909 2363 14943
rect 3341 14909 3375 14943
rect 5834 14909 5868 14943
rect 1777 14841 1811 14875
rect 3249 14841 3283 14875
rect 3893 14841 3927 14875
rect 10241 14841 10275 14875
rect 4445 14773 4479 14807
rect 6929 14773 6963 14807
rect 7573 14773 7607 14807
rect 7665 14773 7699 14807
rect 9137 14773 9171 14807
rect 9229 14773 9263 14807
rect 9781 14773 9815 14807
rect 10149 14773 10183 14807
rect 10793 14773 10827 14807
rect 2237 14569 2271 14603
rect 2697 14569 2731 14603
rect 3157 14569 3191 14603
rect 5733 14569 5767 14603
rect 9505 14569 9539 14603
rect 9965 14569 9999 14603
rect 1777 14501 1811 14535
rect 8042 14501 8076 14535
rect 11078 14501 11112 14535
rect 2329 14433 2363 14467
rect 2881 14433 2915 14467
rect 3341 14433 3375 14467
rect 4609 14433 4643 14467
rect 11345 14433 11379 14467
rect 4353 14365 4387 14399
rect 8309 14365 8343 14399
rect 6009 14297 6043 14331
rect 1685 14229 1719 14263
rect 3985 14229 4019 14263
rect 6929 14229 6963 14263
rect 2145 14025 2179 14059
rect 2973 14025 3007 14059
rect 3985 14025 4019 14059
rect 7021 14025 7055 14059
rect 8585 14025 8619 14059
rect 10977 14025 11011 14059
rect 8309 13957 8343 13991
rect 2605 13889 2639 13923
rect 3617 13889 3651 13923
rect 5365 13889 5399 13923
rect 7665 13889 7699 13923
rect 9229 13889 9263 13923
rect 1593 13821 1627 13855
rect 2329 13821 2363 13855
rect 3433 13821 3467 13855
rect 6469 13821 6503 13855
rect 8125 13821 8159 13855
rect 9597 13821 9631 13855
rect 9853 13821 9887 13855
rect 1777 13753 1811 13787
rect 5098 13753 5132 13787
rect 3341 13685 3375 13719
rect 5733 13685 5767 13719
rect 6009 13685 6043 13719
rect 7389 13685 7423 13719
rect 7481 13685 7515 13719
rect 8953 13685 8987 13719
rect 9045 13685 9079 13719
rect 2145 13481 2179 13515
rect 2605 13481 2639 13515
rect 3065 13481 3099 13515
rect 4537 13481 4571 13515
rect 4997 13481 5031 13515
rect 5457 13481 5491 13515
rect 8309 13481 8343 13515
rect 9413 13481 9447 13515
rect 9873 13481 9907 13515
rect 7174 13413 7208 13447
rect 1777 13345 1811 13379
rect 2329 13345 2363 13379
rect 2789 13345 2823 13379
rect 3249 13345 3283 13379
rect 4261 13345 4295 13379
rect 5365 13345 5399 13379
rect 6009 13345 6043 13379
rect 6653 13345 6687 13379
rect 10986 13345 11020 13379
rect 11253 13345 11287 13379
rect 5549 13277 5583 13311
rect 6929 13277 6963 13311
rect 8585 13277 8619 13311
rect 1593 13209 1627 13243
rect 4077 13209 4111 13243
rect 6469 13209 6503 13243
rect 6193 13141 6227 13175
rect 1777 12937 1811 12971
rect 3709 12937 3743 12971
rect 4169 12937 4203 12971
rect 7481 12937 7515 12971
rect 7757 12937 7791 12971
rect 9597 12937 9631 12971
rect 2973 12869 3007 12903
rect 6009 12869 6043 12903
rect 2329 12801 2363 12835
rect 2513 12801 2547 12835
rect 5549 12801 5583 12835
rect 6929 12801 6963 12835
rect 8309 12801 8343 12835
rect 9229 12801 9263 12835
rect 10241 12801 10275 12835
rect 1961 12733 1995 12767
rect 3433 12733 3467 12767
rect 3893 12733 3927 12767
rect 5825 12733 5859 12767
rect 7113 12733 7147 12767
rect 9965 12733 9999 12767
rect 5282 12665 5316 12699
rect 8125 12665 8159 12699
rect 8217 12665 8251 12699
rect 1409 12597 1443 12631
rect 2605 12597 2639 12631
rect 3249 12597 3283 12631
rect 7021 12597 7055 12631
rect 8769 12597 8803 12631
rect 10057 12597 10091 12631
rect 4077 12393 4111 12427
rect 4997 12393 5031 12427
rect 9873 12393 9907 12427
rect 2982 12325 3016 12359
rect 7012 12325 7046 12359
rect 8309 12325 8343 12359
rect 1409 12257 1443 12291
rect 4261 12257 4295 12291
rect 6110 12257 6144 12291
rect 8585 12257 8619 12291
rect 10986 12257 11020 12291
rect 11253 12257 11287 12291
rect 19809 12257 19843 12291
rect 3249 12189 3283 12223
rect 4721 12189 4755 12223
rect 6377 12189 6411 12223
rect 6745 12189 6779 12223
rect 8309 12189 8343 12223
rect 9137 12189 9171 12223
rect 1593 12053 1627 12087
rect 1869 12053 1903 12087
rect 8125 12053 8159 12087
rect 8401 12053 8435 12087
rect 19993 12053 20027 12087
rect 2697 11849 2731 11883
rect 4629 11849 4663 11883
rect 7021 11849 7055 11883
rect 9965 11849 9999 11883
rect 12081 11849 12115 11883
rect 2145 11713 2179 11747
rect 2980 11713 3014 11747
rect 5181 11713 5215 11747
rect 7665 11713 7699 11747
rect 10609 11713 10643 11747
rect 1501 11645 1535 11679
rect 5641 11645 5675 11679
rect 8309 11645 8343 11679
rect 8565 11645 8599 11679
rect 11897 11645 11931 11679
rect 19165 11645 19199 11679
rect 3218 11577 3252 11611
rect 4997 11577 5031 11611
rect 6469 11577 6503 11611
rect 10333 11577 10367 11611
rect 10977 11577 11011 11611
rect 1685 11509 1719 11543
rect 2237 11509 2271 11543
rect 2329 11509 2363 11543
rect 4353 11509 4387 11543
rect 5089 11509 5123 11543
rect 6009 11509 6043 11543
rect 7389 11509 7423 11543
rect 7481 11509 7515 11543
rect 9689 11509 9723 11543
rect 10425 11509 10459 11543
rect 19349 11509 19383 11543
rect 1593 11305 1627 11339
rect 2237 11305 2271 11339
rect 2697 11305 2731 11339
rect 3157 11305 3191 11339
rect 4261 11305 4295 11339
rect 6009 11305 6043 11339
rect 6837 11305 6871 11339
rect 8493 11305 8527 11339
rect 10885 11305 10919 11339
rect 6285 11237 6319 11271
rect 7380 11237 7414 11271
rect 1409 11169 1443 11203
rect 3065 11169 3099 11203
rect 4077 11169 4111 11203
rect 4896 11169 4930 11203
rect 7113 11169 7147 11203
rect 9505 11169 9539 11203
rect 9772 11169 9806 11203
rect 18705 11169 18739 11203
rect 3249 11101 3283 11135
rect 4629 11101 4663 11135
rect 1869 11033 1903 11067
rect 9137 11033 9171 11067
rect 11161 11033 11195 11067
rect 18889 11033 18923 11067
rect 3065 10761 3099 10795
rect 3341 10761 3375 10795
rect 6837 10761 6871 10795
rect 7389 10761 7423 10795
rect 10057 10761 10091 10795
rect 8033 10625 8067 10659
rect 9597 10625 9631 10659
rect 10609 10625 10643 10659
rect 1685 10557 1719 10591
rect 3525 10557 3559 10591
rect 4077 10557 4111 10591
rect 4344 10557 4378 10591
rect 7021 10557 7055 10591
rect 8769 10557 8803 10591
rect 11897 10557 11931 10591
rect 18245 10557 18279 10591
rect 18705 10557 18739 10591
rect 1952 10489 1986 10523
rect 6469 10489 6503 10523
rect 7757 10489 7791 10523
rect 7849 10489 7883 10523
rect 10517 10489 10551 10523
rect 13645 10489 13679 10523
rect 5457 10421 5491 10455
rect 5733 10421 5767 10455
rect 8585 10421 8619 10455
rect 9045 10421 9079 10455
rect 9413 10421 9447 10455
rect 9505 10421 9539 10455
rect 10425 10421 10459 10455
rect 11069 10421 11103 10455
rect 18429 10421 18463 10455
rect 2053 10217 2087 10251
rect 7021 10217 7055 10251
rect 7481 10217 7515 10251
rect 9413 10217 9447 10251
rect 9781 10217 9815 10251
rect 4997 10149 5031 10183
rect 5089 10149 5123 10183
rect 6009 10149 6043 10183
rect 9873 10149 9907 10183
rect 1409 10081 1443 10115
rect 1869 10081 1903 10115
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 6101 10081 6135 10115
rect 7389 10081 7423 10115
rect 8401 10081 8435 10115
rect 8493 10081 8527 10115
rect 10333 10081 10367 10115
rect 10793 10081 10827 10115
rect 12837 10081 12871 10115
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 4353 10013 4387 10047
rect 5273 10013 5307 10047
rect 6193 10013 6227 10047
rect 7573 10013 7607 10047
rect 8677 10013 8711 10047
rect 9965 10013 9999 10047
rect 1593 9945 1627 9979
rect 5641 9945 5675 9979
rect 13093 10013 13127 10047
rect 11713 9945 11747 9979
rect 3065 9877 3099 9911
rect 3525 9877 3559 9911
rect 4629 9877 4663 9911
rect 6653 9877 6687 9911
rect 8033 9877 8067 9911
rect 10333 9877 10367 9911
rect 10425 9877 10459 9911
rect 11161 9877 11195 9911
rect 13553 9673 13587 9707
rect 3985 9605 4019 9639
rect 4261 9605 4295 9639
rect 6837 9605 6871 9639
rect 9321 9605 9355 9639
rect 10977 9605 11011 9639
rect 2973 9537 3007 9571
rect 3341 9537 3375 9571
rect 4721 9537 4755 9571
rect 4905 9537 4939 9571
rect 8493 9537 8527 9571
rect 8953 9537 8987 9571
rect 3617 9469 3651 9503
rect 4629 9469 4663 9503
rect 6101 9469 6135 9503
rect 8217 9469 8251 9503
rect 10701 9469 10735 9503
rect 11161 9469 11195 9503
rect 11897 9469 11931 9503
rect 2706 9401 2740 9435
rect 6469 9401 6503 9435
rect 7972 9401 8006 9435
rect 10456 9401 10490 9435
rect 12142 9401 12176 9435
rect 1593 9333 1627 9367
rect 3525 9333 3559 9367
rect 5457 9333 5491 9367
rect 5917 9333 5951 9367
rect 13277 9333 13311 9367
rect 2145 9129 2179 9163
rect 3157 9129 3191 9163
rect 3893 9129 3927 9163
rect 4813 9129 4847 9163
rect 7941 9129 7975 9163
rect 8309 9129 8343 9163
rect 8401 9129 8435 9163
rect 9689 9129 9723 9163
rect 11437 9129 11471 9163
rect 11805 9129 11839 9163
rect 12357 9129 12391 9163
rect 13553 9129 13587 9163
rect 14565 9129 14599 9163
rect 3433 9061 3467 9095
rect 10149 9061 10183 9095
rect 1409 8993 1443 9027
rect 2789 8993 2823 9027
rect 6570 8993 6604 9027
rect 7297 8993 7331 9027
rect 10057 8993 10091 9027
rect 12449 8993 12483 9027
rect 13093 8993 13127 9027
rect 15678 8993 15712 9027
rect 2605 8925 2639 8959
rect 2697 8925 2731 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 6837 8925 6871 8959
rect 6929 8925 6963 8959
rect 8585 8925 8619 8959
rect 10241 8925 10275 8959
rect 11253 8925 11287 8959
rect 11345 8925 11379 8959
rect 12265 8925 12299 8959
rect 15945 8925 15979 8959
rect 7573 8857 7607 8891
rect 1593 8789 1627 8823
rect 4445 8789 4479 8823
rect 5457 8789 5491 8823
rect 6929 8789 6963 8823
rect 7113 8789 7147 8823
rect 9137 8789 9171 8823
rect 10701 8789 10735 8823
rect 12817 8789 12851 8823
rect 14013 8789 14047 8823
rect 1593 8585 1627 8619
rect 3801 8585 3835 8619
rect 8677 8585 8711 8619
rect 9137 8585 9171 8619
rect 10609 8585 10643 8619
rect 13093 8585 13127 8619
rect 3341 8517 3375 8551
rect 5733 8517 5767 8551
rect 12633 8517 12667 8551
rect 14841 8517 14875 8551
rect 17325 8517 17359 8551
rect 10241 8449 10275 8483
rect 11069 8449 11103 8483
rect 11989 8449 12023 8483
rect 13461 8449 13495 8483
rect 15301 8449 15335 8483
rect 1409 8381 1443 8415
rect 1961 8381 1995 8415
rect 3617 8381 3651 8415
rect 4353 8381 4387 8415
rect 4620 8381 4654 8415
rect 8134 8381 8168 8415
rect 8401 8381 8435 8415
rect 8493 8381 8527 8415
rect 8861 8381 8895 8415
rect 9321 8381 9355 8415
rect 9965 8381 9999 8415
rect 12909 8381 12943 8415
rect 17141 8381 17175 8415
rect 2228 8313 2262 8347
rect 6009 8313 6043 8347
rect 6469 8313 6503 8347
rect 12173 8313 12207 8347
rect 13728 8313 13762 8347
rect 15485 8313 15519 8347
rect 16129 8313 16163 8347
rect 7021 8245 7055 8279
rect 8493 8245 8527 8279
rect 9781 8245 9815 8279
rect 12265 8245 12299 8279
rect 15393 8245 15427 8279
rect 15853 8245 15887 8279
rect 1409 8041 1443 8075
rect 2789 8041 2823 8075
rect 4353 8041 4387 8075
rect 4721 8041 4755 8075
rect 5733 8041 5767 8075
rect 6561 8041 6595 8075
rect 7665 8041 7699 8075
rect 8033 8041 8067 8075
rect 9597 8041 9631 8075
rect 11897 8041 11931 8075
rect 13921 8041 13955 8075
rect 14841 8041 14875 8075
rect 15301 8041 15335 8075
rect 3157 7973 3191 8007
rect 13286 7973 13320 8007
rect 14933 7973 14967 8007
rect 2053 7905 2087 7939
rect 2145 7905 2179 7939
rect 5273 7905 5307 7939
rect 6377 7905 6411 7939
rect 7021 7905 7055 7939
rect 8493 7905 8527 7939
rect 9689 7905 9723 7939
rect 10517 7905 10551 7939
rect 10784 7905 10818 7939
rect 13553 7905 13587 7939
rect 15761 7905 15795 7939
rect 17334 7905 17368 7939
rect 1961 7837 1995 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 2513 7769 2547 7803
rect 5825 7837 5859 7871
rect 6009 7837 6043 7871
rect 7481 7837 7515 7871
rect 7573 7837 7607 7871
rect 9413 7837 9447 7871
rect 14749 7837 14783 7871
rect 17601 7837 17635 7871
rect 8309 7769 8343 7803
rect 12173 7769 12207 7803
rect 16221 7769 16255 7803
rect 3985 7701 4019 7735
rect 5273 7701 5307 7735
rect 5365 7701 5399 7735
rect 6837 7701 6871 7735
rect 10057 7701 10091 7735
rect 15945 7701 15979 7735
rect 3157 7497 3191 7531
rect 5181 7497 5215 7531
rect 6469 7497 6503 7531
rect 6653 7497 6687 7531
rect 12633 7497 12667 7531
rect 15025 7497 15059 7531
rect 3617 7429 3651 7463
rect 5641 7361 5675 7395
rect 5733 7361 5767 7395
rect 1777 7293 1811 7327
rect 3433 7293 3467 7327
rect 3893 7293 3927 7327
rect 4353 7293 4387 7327
rect 4813 7293 4847 7327
rect 9045 7429 9079 7463
rect 7205 7361 7239 7395
rect 11345 7361 11379 7395
rect 11989 7361 12023 7395
rect 13369 7361 13403 7395
rect 7665 7293 7699 7327
rect 7932 7293 7966 7327
rect 9321 7293 9355 7327
rect 9577 7293 9611 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 12909 7293 12943 7327
rect 16405 7293 16439 7327
rect 2022 7225 2056 7259
rect 5549 7225 5583 7259
rect 6469 7225 6503 7259
rect 7021 7225 7055 7259
rect 13614 7225 13648 7259
rect 16138 7225 16172 7259
rect 16957 7225 16991 7259
rect 1409 7157 1443 7191
rect 4077 7157 4111 7191
rect 4537 7157 4571 7191
rect 7113 7157 7147 7191
rect 10701 7157 10735 7191
rect 14749 7157 14783 7191
rect 3157 6953 3191 6987
rect 2145 6885 2179 6919
rect 1501 6817 1535 6851
rect 5190 6817 5224 6851
rect 5917 6817 5951 6851
rect 6377 6817 6411 6851
rect 7021 6817 7055 6851
rect 7113 6817 7147 6851
rect 7757 6817 7791 6851
rect 8401 6817 8435 6851
rect 9505 6817 9539 6851
rect 9965 6817 9999 6851
rect 10865 6817 10899 6851
rect 12449 6817 12483 6851
rect 12909 6817 12943 6851
rect 13093 6817 13127 6851
rect 13553 6817 13587 6851
rect 14933 6817 14967 6851
rect 15577 6817 15611 6851
rect 17242 6817 17276 6851
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 5457 6749 5491 6783
rect 6929 6749 6963 6783
rect 8677 6749 8711 6783
rect 10609 6749 10643 6783
rect 2789 6681 2823 6715
rect 4077 6681 4111 6715
rect 6193 6681 6227 6715
rect 7481 6681 7515 6715
rect 9781 6681 9815 6715
rect 15025 6749 15059 6783
rect 15117 6749 15151 6783
rect 17509 6749 17543 6783
rect 15761 6681 15795 6715
rect 1777 6613 1811 6647
rect 5733 6613 5767 6647
rect 8217 6613 8251 6647
rect 10241 6613 10275 6647
rect 11989 6613 12023 6647
rect 12265 6613 12299 6647
rect 12725 6613 12759 6647
rect 12909 6613 12943 6647
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 14565 6613 14599 6647
rect 16129 6613 16163 6647
rect 1409 6409 1443 6443
rect 13553 6409 13587 6443
rect 14565 6409 14599 6443
rect 16589 6409 16623 6443
rect 2973 6341 3007 6375
rect 4629 6341 4663 6375
rect 9873 6341 9907 6375
rect 2789 6205 2823 6239
rect 3065 6273 3099 6307
rect 4169 6273 4203 6307
rect 6009 6273 6043 6307
rect 6837 6273 6871 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 13921 6273 13955 6307
rect 15025 6273 15059 6307
rect 16037 6273 16071 6307
rect 17693 6273 17727 6307
rect 3985 6205 4019 6239
rect 6561 6205 6595 6239
rect 7093 6205 7127 6239
rect 8493 6205 8527 6239
rect 10517 6205 10551 6239
rect 11345 6205 11379 6239
rect 12173 6205 12207 6239
rect 12429 6205 12463 6239
rect 15393 6205 15427 6239
rect 17601 6205 17635 6239
rect 18153 6205 18187 6239
rect 2544 6137 2578 6171
rect 2973 6137 3007 6171
rect 5742 6137 5776 6171
rect 8738 6137 8772 6171
rect 14197 6137 14231 6171
rect 16221 6137 16255 6171
rect 3617 6069 3651 6103
rect 4077 6069 4111 6103
rect 8217 6069 8251 6103
rect 10885 6069 10919 6103
rect 11161 6069 11195 6103
rect 11713 6069 11747 6103
rect 14105 6069 14139 6103
rect 15577 6069 15611 6103
rect 16129 6069 16163 6103
rect 17141 6069 17175 6103
rect 17509 6069 17543 6103
rect 2145 5865 2179 5899
rect 2513 5865 2547 5899
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 7389 5865 7423 5899
rect 12357 5865 12391 5899
rect 15393 5865 15427 5899
rect 16405 5865 16439 5899
rect 17601 5865 17635 5899
rect 3157 5797 3191 5831
rect 8033 5797 8067 5831
rect 9680 5797 9714 5831
rect 13553 5797 13587 5831
rect 16773 5797 16807 5831
rect 5089 5729 5123 5763
rect 5733 5729 5767 5763
rect 6276 5729 6310 5763
rect 9413 5729 9447 5763
rect 11713 5729 11747 5763
rect 12449 5729 12483 5763
rect 13093 5729 13127 5763
rect 14565 5729 14599 5763
rect 17969 5729 18003 5763
rect 20913 5729 20947 5763
rect 21373 5729 21407 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 3433 5661 3467 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 6009 5661 6043 5695
rect 7757 5661 7791 5695
rect 7941 5661 7975 5695
rect 11069 5661 11103 5695
rect 12173 5661 12207 5695
rect 13921 5661 13955 5695
rect 15025 5661 15059 5695
rect 16865 5661 16899 5695
rect 17049 5661 17083 5695
rect 2789 5593 2823 5627
rect 5273 5593 5307 5627
rect 8677 5593 8711 5627
rect 11529 5593 11563 5627
rect 18245 5593 18279 5627
rect 1501 5525 1535 5559
rect 5549 5525 5583 5559
rect 8401 5525 8435 5559
rect 10793 5525 10827 5559
rect 12817 5525 12851 5559
rect 14749 5525 14783 5559
rect 15761 5525 15795 5559
rect 21189 5525 21223 5559
rect 5917 5321 5951 5355
rect 7757 5321 7791 5355
rect 8769 5321 8803 5355
rect 11897 5321 11931 5355
rect 12357 5321 12391 5355
rect 17141 5321 17175 5355
rect 1869 5253 1903 5287
rect 4537 5253 4571 5287
rect 11069 5253 11103 5287
rect 14105 5253 14139 5287
rect 16221 5253 16255 5287
rect 2605 5185 2639 5219
rect 3433 5185 3467 5219
rect 6469 5185 6503 5219
rect 7113 5185 7147 5219
rect 8217 5185 8251 5219
rect 8309 5185 8343 5219
rect 9505 5185 9539 5219
rect 10517 5185 10551 5219
rect 15669 5185 15703 5219
rect 1685 5117 1719 5151
rect 3893 5117 3927 5151
rect 4353 5117 4387 5151
rect 4813 5117 4847 5151
rect 5273 5117 5307 5151
rect 5733 5117 5767 5151
rect 7389 5117 7423 5151
rect 9597 5117 9631 5151
rect 10701 5117 10735 5151
rect 12081 5117 12115 5151
rect 12541 5117 12575 5151
rect 12909 5117 12943 5151
rect 14473 5117 14507 5151
rect 14933 5117 14967 5151
rect 15853 5117 15887 5151
rect 18521 5117 18555 5151
rect 2789 5049 2823 5083
rect 8401 5049 8435 5083
rect 9689 5049 9723 5083
rect 15761 5049 15795 5083
rect 18254 5049 18288 5083
rect 2697 4981 2731 5015
rect 3157 4981 3191 5015
rect 4077 4981 4111 5015
rect 4997 4981 5031 5015
rect 5457 4981 5491 5015
rect 7297 4981 7331 5015
rect 10057 4981 10091 5015
rect 10609 4981 10643 5015
rect 13093 4981 13127 5015
rect 13369 4981 13403 5015
rect 13737 4981 13771 5015
rect 14657 4981 14691 5015
rect 15117 4981 15151 5015
rect 16589 4981 16623 5015
rect 1777 4777 1811 4811
rect 2145 4777 2179 4811
rect 2421 4777 2455 4811
rect 7849 4777 7883 4811
rect 8585 4777 8619 4811
rect 9597 4777 9631 4811
rect 10057 4777 10091 4811
rect 12173 4777 12207 4811
rect 17233 4777 17267 4811
rect 2881 4709 2915 4743
rect 7481 4709 7515 4743
rect 10784 4709 10818 4743
rect 16098 4709 16132 4743
rect 18705 4709 18739 4743
rect 21128 4709 21162 4743
rect 1685 4641 1719 4675
rect 2789 4641 2823 4675
rect 4077 4641 4111 4675
rect 4721 4641 4755 4675
rect 5549 4641 5583 4675
rect 6193 4641 6227 4675
rect 6837 4641 6871 4675
rect 7389 4641 7423 4675
rect 8309 4641 8343 4675
rect 8769 4641 8803 4675
rect 9413 4641 9447 4675
rect 9873 4641 9907 4675
rect 12357 4641 12391 4675
rect 12817 4641 12851 4675
rect 13277 4641 13311 4675
rect 13645 4641 13679 4675
rect 14565 4641 14599 4675
rect 15393 4641 15427 4675
rect 15853 4641 15887 4675
rect 21373 4641 21407 4675
rect 1593 4573 1627 4607
rect 2973 4573 3007 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 7205 4573 7239 4607
rect 10517 4573 10551 4607
rect 12449 4573 12483 4607
rect 15025 4573 15059 4607
rect 17509 4573 17543 4607
rect 8125 4505 8159 4539
rect 13093 4505 13127 4539
rect 13829 4505 13863 4539
rect 19993 4505 20027 4539
rect 3433 4437 3467 4471
rect 4261 4437 4295 4471
rect 4537 4437 4571 4471
rect 5917 4437 5951 4471
rect 6377 4437 6411 4471
rect 6653 4437 6687 4471
rect 11897 4437 11931 4471
rect 12449 4437 12483 4471
rect 12633 4437 12667 4471
rect 14749 4437 14783 4471
rect 15577 4437 15611 4471
rect 18061 4437 18095 4471
rect 18337 4437 18371 4471
rect 1593 4233 1627 4267
rect 3341 4233 3375 4267
rect 8033 4233 8067 4267
rect 16405 4233 16439 4267
rect 4997 4165 5031 4199
rect 17877 4165 17911 4199
rect 5917 4097 5951 4131
rect 6653 4097 6687 4131
rect 8125 4097 8159 4131
rect 10793 4097 10827 4131
rect 13737 4097 13771 4131
rect 17325 4097 17359 4131
rect 17417 4097 17451 4131
rect 1501 4029 1535 4063
rect 1961 4029 1995 4063
rect 2228 4029 2262 4063
rect 3617 4029 3651 4063
rect 3862 3961 3896 3995
rect 6920 3961 6954 3995
rect 9689 4029 9723 4063
rect 10885 4029 10919 4063
rect 10977 4029 11011 4063
rect 11897 4029 11931 4063
rect 12153 4029 12187 4063
rect 14565 4029 14599 4063
rect 15025 4029 15059 4063
rect 17509 4029 17543 4063
rect 18153 4029 18187 4063
rect 18613 4029 18647 4063
rect 20177 4029 20211 4063
rect 20453 4029 20487 4063
rect 21097 4029 21131 4063
rect 9444 3961 9478 3995
rect 13921 3961 13955 3995
rect 15292 3961 15326 3995
rect 20913 3961 20947 3995
rect 5273 3893 5307 3927
rect 5641 3893 5675 3927
rect 5733 3893 5767 3927
rect 8125 3893 8159 3927
rect 8309 3893 8343 3927
rect 9965 3893 9999 3927
rect 11345 3893 11379 3927
rect 13277 3893 13311 3927
rect 13829 3893 13863 3927
rect 14289 3893 14323 3927
rect 14749 3893 14783 3927
rect 18337 3893 18371 3927
rect 18797 3893 18831 3927
rect 19073 3893 19107 3927
rect 19809 3893 19843 3927
rect 20637 3893 20671 3927
rect 1501 3689 1535 3723
rect 5917 3689 5951 3723
rect 8401 3689 8435 3723
rect 9137 3689 9171 3723
rect 10057 3689 10091 3723
rect 10701 3689 10735 3723
rect 14013 3689 14047 3723
rect 15945 3689 15979 3723
rect 19073 3689 19107 3723
rect 21189 3689 21223 3723
rect 2636 3621 2670 3655
rect 6438 3621 6472 3655
rect 12900 3621 12934 3655
rect 14810 3621 14844 3655
rect 16405 3621 16439 3655
rect 20269 3621 20303 3655
rect 20821 3621 20855 3655
rect 3341 3553 3375 3587
rect 4069 3553 4103 3587
rect 4537 3553 4571 3587
rect 4804 3553 4838 3587
rect 10149 3553 10183 3587
rect 10885 3553 10919 3587
rect 11161 3553 11195 3587
rect 11713 3553 11747 3587
rect 14565 3553 14599 3587
rect 17417 3553 17451 3587
rect 17693 3553 17727 3587
rect 18153 3553 18187 3587
rect 18797 3553 18831 3587
rect 19257 3553 19291 3587
rect 21373 3553 21407 3587
rect 2881 3485 2915 3519
rect 6193 3485 6227 3519
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 8953 3485 8987 3519
rect 10241 3485 10275 3519
rect 12357 3485 12391 3519
rect 12633 3485 12667 3519
rect 16773 3485 16807 3519
rect 16221 3417 16255 3451
rect 18337 3417 18371 3451
rect 20085 3417 20119 3451
rect 20637 3417 20671 3451
rect 3249 3349 3283 3383
rect 4261 3349 4295 3383
rect 7573 3349 7607 3383
rect 8033 3349 8067 3383
rect 8953 3349 8987 3383
rect 9689 3349 9723 3383
rect 11345 3349 11379 3383
rect 11897 3349 11931 3383
rect 17233 3349 17267 3383
rect 17877 3349 17911 3383
rect 18613 3349 18647 3383
rect 19809 3349 19843 3383
rect 1777 3145 1811 3179
rect 2881 3145 2915 3179
rect 3065 3145 3099 3179
rect 13277 3145 13311 3179
rect 15853 3145 15887 3179
rect 2973 3077 3007 3111
rect 2329 3009 2363 3043
rect 1685 2941 1719 2975
rect 2421 2873 2455 2907
rect 5181 3077 5215 3111
rect 5089 3009 5123 3043
rect 8585 3077 8619 3111
rect 5549 3009 5583 3043
rect 7297 3009 7331 3043
rect 7757 3009 7791 3043
rect 7941 3009 7975 3043
rect 4281 2941 4315 2975
rect 4537 2941 4571 2975
rect 5181 2941 5215 2975
rect 5733 2941 5767 2975
rect 7113 2941 7147 2975
rect 8033 2941 8067 2975
rect 3065 2873 3099 2907
rect 5641 2873 5675 2907
rect 7021 2873 7055 2907
rect 10057 3009 10091 3043
rect 10977 3009 11011 3043
rect 12725 3009 12759 3043
rect 15301 3009 15335 3043
rect 20545 3009 20579 3043
rect 10793 2941 10827 2975
rect 11897 2941 11931 2975
rect 12909 2941 12943 2975
rect 13553 2941 13587 2975
rect 14013 2941 14047 2975
rect 14657 2941 14691 2975
rect 15393 2941 15427 2975
rect 15485 2941 15519 2975
rect 17325 2941 17359 2975
rect 17877 2941 17911 2975
rect 18337 2941 18371 2975
rect 18797 2941 18831 2975
rect 19349 2941 19383 2975
rect 19901 2941 19935 2975
rect 21189 2941 21223 2975
rect 9812 2873 9846 2907
rect 14841 2873 14875 2907
rect 16129 2873 16163 2907
rect 16313 2873 16347 2907
rect 17141 2873 17175 2907
rect 19165 2873 19199 2907
rect 19717 2873 19751 2907
rect 2513 2805 2547 2839
rect 2973 2805 3007 2839
rect 3157 2805 3191 2839
rect 6101 2805 6135 2839
rect 6653 2805 6687 2839
rect 8401 2805 8435 2839
rect 8585 2805 8619 2839
rect 8677 2805 8711 2839
rect 10333 2805 10367 2839
rect 10701 2805 10735 2839
rect 12081 2805 12115 2839
rect 12817 2805 12851 2839
rect 13737 2805 13771 2839
rect 14197 2805 14231 2839
rect 17693 2805 17727 2839
rect 18153 2805 18187 2839
rect 18613 2805 18647 2839
rect 2697 2601 2731 2635
rect 3065 2601 3099 2635
rect 4721 2601 4755 2635
rect 5825 2601 5859 2635
rect 6745 2601 6779 2635
rect 7205 2601 7239 2635
rect 8493 2601 8527 2635
rect 8861 2601 8895 2635
rect 9873 2601 9907 2635
rect 9965 2601 9999 2635
rect 12265 2601 12299 2635
rect 12357 2601 12391 2635
rect 20269 2601 20303 2635
rect 1685 2533 1719 2567
rect 2421 2533 2455 2567
rect 5733 2533 5767 2567
rect 7113 2533 7147 2567
rect 2237 2465 2271 2499
rect 3157 2465 3191 2499
rect 4261 2465 4295 2499
rect 4813 2465 4847 2499
rect 7757 2465 7791 2499
rect 10701 2465 10735 2499
rect 10977 2465 11011 2499
rect 11345 2465 11379 2499
rect 12081 2465 12115 2499
rect 12725 2533 12759 2567
rect 13829 2533 13863 2567
rect 14933 2533 14967 2567
rect 15485 2533 15519 2567
rect 16037 2533 16071 2567
rect 17601 2533 17635 2567
rect 18153 2533 18187 2567
rect 18705 2533 18739 2567
rect 19257 2533 19291 2567
rect 20637 2533 20671 2567
rect 13277 2465 13311 2499
rect 16681 2465 16715 2499
rect 20085 2465 20119 2499
rect 21281 2465 21315 2499
rect 3249 2397 3283 2431
rect 5641 2397 5675 2431
rect 7297 2397 7331 2431
rect 8309 2397 8343 2431
rect 8401 2397 8435 2431
rect 10057 2397 10091 2431
rect 12357 2397 12391 2431
rect 16865 2397 16899 2431
rect 19073 2397 19107 2431
rect 1869 2329 1903 2363
rect 9505 2329 9539 2363
rect 11529 2329 11563 2363
rect 12541 2329 12575 2363
rect 13093 2329 13127 2363
rect 13645 2329 13679 2363
rect 14749 2329 14783 2363
rect 15853 2329 15887 2363
rect 17417 2329 17451 2363
rect 17969 2329 18003 2363
rect 20821 2329 20855 2363
rect 4169 2261 4203 2295
rect 6193 2261 6227 2295
rect 10517 2261 10551 2295
rect 15393 2261 15427 2295
rect 18613 2261 18647 2295
rect 21189 2261 21223 2295
rect 13921 1989 13955 2023
rect 13921 1853 13955 1887
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 2685 20519 2743 20525
rect 2685 20485 2697 20519
rect 2731 20516 2743 20519
rect 2774 20516 2780 20528
rect 2731 20488 2780 20516
rect 2731 20485 2743 20488
rect 2685 20479 2743 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 3234 20516 3240 20528
rect 3195 20488 3240 20516
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 4062 20516 4068 20528
rect 4023 20488 4068 20516
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 2866 20448 2872 20460
rect 1688 20420 2872 20448
rect 1688 20389 1716 20420
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20349 1731 20383
rect 1673 20343 1731 20349
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 1903 20352 2452 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 2130 20312 2136 20324
rect 2091 20284 2136 20312
rect 2130 20272 2136 20284
rect 2188 20272 2194 20324
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 2424 20244 2452 20352
rect 2866 20312 2872 20324
rect 2827 20284 2872 20312
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 3418 20312 3424 20324
rect 3379 20284 3424 20312
rect 3418 20272 3424 20284
rect 3476 20272 3482 20324
rect 4249 20315 4307 20321
rect 4249 20281 4261 20315
rect 4295 20312 4307 20315
rect 10594 20312 10600 20324
rect 4295 20284 10600 20312
rect 4295 20281 4307 20284
rect 4249 20275 4307 20281
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 2774 20244 2780 20256
rect 2424 20216 2780 20244
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2222 20040 2228 20052
rect 2183 20012 2228 20040
rect 2222 20000 2228 20012
rect 2280 20000 2286 20052
rect 2866 20040 2872 20052
rect 2827 20012 2872 20040
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 2958 20000 2964 20052
rect 3016 20040 3022 20052
rect 3145 20043 3203 20049
rect 3145 20040 3157 20043
rect 3016 20012 3157 20040
rect 3016 20000 3022 20012
rect 3145 20009 3157 20012
rect 3191 20009 3203 20043
rect 3145 20003 3203 20009
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2222 19904 2228 19916
rect 1811 19876 2228 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19904 2375 19907
rect 2590 19904 2596 19916
rect 2363 19876 2596 19904
rect 2363 19873 2375 19876
rect 2317 19867 2375 19873
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19904 2743 19907
rect 4062 19904 4068 19916
rect 2731 19876 4068 19904
rect 2731 19873 2743 19876
rect 2685 19867 2743 19873
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 2590 19496 2596 19508
rect 2551 19468 2596 19496
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 3237 19499 3295 19505
rect 3237 19465 3249 19499
rect 3283 19496 3295 19499
rect 3418 19496 3424 19508
rect 3283 19468 3424 19496
rect 3283 19465 3295 19468
rect 3237 19459 3295 19465
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19261 2191 19295
rect 2133 19255 2191 19261
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2958 19292 2964 19304
rect 2823 19264 2964 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 1762 19224 1768 19236
rect 1723 19196 1768 19224
rect 1762 19184 1768 19196
rect 1820 19184 1826 19236
rect 2148 19224 2176 19255
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 3602 19292 3608 19304
rect 3099 19264 3608 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3602 19252 3608 19264
rect 3660 19252 3666 19304
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 8570 19292 8576 19304
rect 3743 19264 8576 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 2148 19196 3556 19224
rect 3528 19165 3556 19196
rect 3513 19159 3571 19165
rect 3513 19125 3525 19159
rect 3559 19125 3571 19159
rect 3513 19119 3571 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1762 18912 1768 18964
rect 1820 18952 1826 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1820 18924 2145 18952
rect 1820 18912 1826 18924
rect 2133 18921 2145 18924
rect 2179 18921 2191 18955
rect 2133 18915 2191 18921
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2593 18955 2651 18961
rect 2593 18952 2605 18955
rect 2280 18924 2605 18952
rect 2280 18912 2286 18924
rect 2593 18921 2605 18924
rect 2639 18921 2651 18955
rect 2593 18915 2651 18921
rect 2958 18912 2964 18964
rect 3016 18952 3022 18964
rect 3053 18955 3111 18961
rect 3053 18952 3065 18955
rect 3016 18924 3065 18952
rect 3016 18912 3022 18924
rect 3053 18921 3065 18924
rect 3099 18921 3111 18955
rect 3053 18915 3111 18921
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 3660 18924 4537 18952
rect 3660 18912 3666 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 10594 18952 10600 18964
rect 10555 18924 10600 18952
rect 4525 18915 4583 18921
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 1578 18884 1584 18896
rect 1539 18856 1584 18884
rect 1578 18844 1584 18856
rect 1636 18844 1642 18896
rect 8662 18884 8668 18896
rect 3252 18856 8668 18884
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 2777 18819 2835 18825
rect 2777 18785 2789 18819
rect 2823 18816 2835 18819
rect 3142 18816 3148 18828
rect 2823 18788 3148 18816
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 2332 18748 2360 18779
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 3252 18825 3280 18856
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18785 3295 18819
rect 3237 18779 3295 18785
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 9582 18816 9588 18828
rect 4755 18788 9588 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 3050 18748 3056 18760
rect 2332 18720 3056 18748
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 4264 18748 4292 18779
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 11238 18816 11244 18828
rect 10827 18788 11244 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 11238 18776 11244 18788
rect 11296 18776 11302 18828
rect 6822 18748 6828 18760
rect 4264 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 4062 18680 4068 18692
rect 4023 18652 4068 18680
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 3142 18408 3148 18420
rect 3103 18380 3148 18408
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 9582 18408 9588 18420
rect 9543 18380 9588 18408
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 1762 18300 1768 18352
rect 1820 18340 1826 18352
rect 2685 18343 2743 18349
rect 2685 18340 2697 18343
rect 1820 18312 2697 18340
rect 1820 18300 1826 18312
rect 2685 18309 2697 18312
rect 2731 18309 2743 18343
rect 2685 18303 2743 18309
rect 10226 18272 10232 18284
rect 10187 18244 10232 18272
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 2866 18204 2872 18216
rect 2827 18176 2872 18204
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18204 3387 18207
rect 9858 18204 9864 18216
rect 3375 18176 9864 18204
rect 3375 18173 3387 18176
rect 3329 18167 3387 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 1762 18136 1768 18148
rect 1723 18108 1768 18136
rect 1762 18096 1768 18108
rect 1820 18096 1826 18148
rect 2314 18136 2320 18148
rect 2275 18108 2320 18136
rect 2314 18096 2320 18108
rect 2372 18096 2378 18148
rect 9953 18139 10011 18145
rect 9953 18105 9965 18139
rect 9999 18136 10011 18139
rect 11054 18136 11060 18148
rect 9999 18108 11060 18136
rect 9999 18105 10011 18108
rect 9953 18099 10011 18105
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 6089 18071 6147 18077
rect 6089 18037 6101 18071
rect 6135 18068 6147 18071
rect 7282 18068 7288 18080
rect 6135 18040 7288 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10100 18040 10145 18068
rect 10100 18028 10106 18040
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1820 17836 2145 17864
rect 1820 17824 1826 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 2866 17864 2872 17876
rect 2823 17836 2872 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3050 17864 3056 17876
rect 3011 17836 3056 17864
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3697 17867 3755 17873
rect 3697 17833 3709 17867
rect 3743 17864 3755 17867
rect 6914 17864 6920 17876
rect 3743 17836 6920 17864
rect 3743 17833 3755 17836
rect 3697 17827 3755 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7282 17864 7288 17876
rect 7243 17836 7288 17864
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17833 7987 17867
rect 7929 17827 7987 17833
rect 2746 17768 6776 17796
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2498 17728 2504 17740
rect 2363 17700 2504 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2498 17688 2504 17700
rect 2556 17688 2562 17740
rect 2593 17731 2651 17737
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 2746 17728 2774 17768
rect 5534 17737 5540 17740
rect 2639 17700 2774 17728
rect 3237 17731 3295 17737
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 3237 17697 3249 17731
rect 3283 17728 3295 17731
rect 3697 17731 3755 17737
rect 3697 17728 3709 17731
rect 3283 17700 3709 17728
rect 3283 17697 3295 17700
rect 3237 17691 3295 17697
rect 3697 17697 3709 17700
rect 3743 17697 3755 17731
rect 3697 17691 3755 17697
rect 5528 17691 5540 17737
rect 5592 17728 5598 17740
rect 6748 17728 6776 17768
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 7944 17796 7972 17827
rect 10226 17824 10232 17876
rect 10284 17864 10290 17876
rect 10870 17864 10876 17876
rect 10284 17836 10876 17864
rect 10284 17824 10290 17836
rect 10870 17824 10876 17836
rect 10928 17864 10934 17876
rect 10965 17867 11023 17873
rect 10965 17864 10977 17867
rect 10928 17836 10977 17864
rect 10928 17824 10934 17836
rect 10965 17833 10977 17836
rect 11011 17833 11023 17867
rect 11238 17864 11244 17876
rect 11199 17836 11244 17864
rect 10965 17827 11023 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 6880 17768 7972 17796
rect 6880 17756 6886 17768
rect 9766 17756 9772 17808
rect 9824 17805 9830 17808
rect 9824 17799 9888 17805
rect 9824 17765 9842 17799
rect 9876 17765 9888 17799
rect 9824 17759 9888 17765
rect 9824 17756 9830 17759
rect 7006 17728 7012 17740
rect 5592 17700 5628 17728
rect 6748 17700 7012 17728
rect 5534 17688 5540 17691
rect 5592 17688 5598 17700
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 8294 17728 8300 17740
rect 8255 17700 8300 17728
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9585 17731 9643 17737
rect 9585 17728 9597 17731
rect 9180 17700 9597 17728
rect 9180 17688 9186 17700
rect 9585 17697 9597 17700
rect 9631 17697 9643 17731
rect 9585 17691 9643 17697
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 11882 17728 11888 17740
rect 11471 17700 11888 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 5261 17663 5319 17669
rect 5261 17660 5273 17663
rect 4856 17632 5273 17660
rect 4856 17620 4862 17632
rect 5261 17629 5273 17632
rect 5307 17629 5319 17663
rect 7374 17660 7380 17672
rect 7335 17632 7380 17660
rect 5261 17623 5319 17629
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17629 7527 17663
rect 8386 17660 8392 17672
rect 8347 17632 8392 17660
rect 7469 17623 7527 17629
rect 6917 17595 6975 17601
rect 6917 17592 6929 17595
rect 6196 17564 6929 17592
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 6196 17524 6224 17564
rect 6917 17561 6929 17564
rect 6963 17561 6975 17595
rect 6917 17555 6975 17561
rect 6638 17524 6644 17536
rect 3752 17496 6224 17524
rect 6599 17496 6644 17524
rect 3752 17484 3758 17496
rect 6638 17484 6644 17496
rect 6696 17524 6702 17536
rect 7484 17524 7512 17623
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 9490 17660 9496 17672
rect 8619 17632 9496 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 6696 17496 7512 17524
rect 6696 17484 6702 17496
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 2133 17323 2191 17329
rect 2133 17320 2145 17323
rect 1820 17292 2145 17320
rect 1820 17280 1826 17292
rect 2133 17289 2145 17292
rect 2179 17289 2191 17323
rect 2133 17283 2191 17289
rect 2314 17280 2320 17332
rect 2372 17320 2378 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 2372 17292 2605 17320
rect 2372 17280 2378 17292
rect 2593 17289 2605 17292
rect 2639 17289 2651 17323
rect 2593 17283 2651 17289
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5592 17292 5733 17320
rect 5592 17280 5598 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 5721 17283 5779 17289
rect 2498 17212 2504 17264
rect 2556 17252 2562 17264
rect 3513 17255 3571 17261
rect 3513 17252 3525 17255
rect 2556 17224 3525 17252
rect 2556 17212 2562 17224
rect 3513 17221 3525 17224
rect 3559 17221 3571 17255
rect 3513 17215 3571 17221
rect 5736 17184 5764 17283
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 11882 17320 11888 17332
rect 11843 17292 11888 17320
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 5736 17156 6745 17184
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 11054 17184 11060 17196
rect 11015 17156 11060 17184
rect 6733 17147 6791 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17184 12587 17187
rect 13630 17184 13636 17196
rect 12575 17156 13636 17184
rect 12575 17153 12587 17156
rect 12529 17147 12587 17153
rect 13630 17144 13636 17156
rect 13688 17184 13694 17196
rect 21358 17184 21364 17196
rect 13688 17156 21220 17184
rect 21319 17156 21364 17184
rect 13688 17144 13694 17156
rect 2314 17116 2320 17128
rect 2275 17088 2320 17116
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 1578 17048 1584 17060
rect 1539 17020 1584 17048
rect 1578 17008 1584 17020
rect 1636 17008 1642 17060
rect 1762 17048 1768 17060
rect 1723 17020 1768 17048
rect 1762 17008 1768 17020
rect 1820 17008 1826 17060
rect 2792 17048 2820 17079
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 3016 17088 3249 17116
rect 3016 17076 3022 17088
rect 3237 17085 3249 17088
rect 3283 17085 3295 17119
rect 3694 17116 3700 17128
rect 3655 17088 3700 17116
rect 3237 17079 3295 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 9122 17116 9128 17128
rect 4387 17088 4844 17116
rect 9083 17088 9128 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4816 17060 4844 17088
rect 9122 17076 9128 17088
rect 9180 17116 9186 17128
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 9180 17088 9413 17116
rect 9180 17076 9186 17088
rect 9401 17085 9413 17088
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 21192 17125 21220 17156
rect 21358 17144 21364 17156
rect 21416 17144 21422 17196
rect 9657 17119 9715 17125
rect 9657 17116 9669 17119
rect 9548 17088 9669 17116
rect 9548 17076 9554 17088
rect 9657 17085 9669 17088
rect 9703 17085 9715 17119
rect 9657 17079 9715 17085
rect 21177 17119 21235 17125
rect 21177 17085 21189 17119
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 2792 17020 3924 17048
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 2924 16952 3065 16980
rect 2924 16940 2930 16952
rect 3053 16949 3065 16952
rect 3099 16949 3111 16983
rect 3896 16980 3924 17020
rect 4062 17008 4068 17060
rect 4120 17048 4126 17060
rect 4586 17051 4644 17057
rect 4586 17048 4598 17051
rect 4120 17020 4598 17048
rect 4120 17008 4126 17020
rect 4586 17017 4598 17020
rect 4632 17017 4644 17051
rect 4586 17011 4644 17017
rect 4798 17008 4804 17060
rect 4856 17008 4862 17060
rect 6917 17051 6975 17057
rect 6917 17017 6929 17051
rect 6963 17048 6975 17051
rect 7282 17048 7288 17060
rect 6963 17020 7288 17048
rect 6963 17017 6975 17020
rect 6917 17011 6975 17017
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 8938 17057 8944 17060
rect 8880 17051 8944 17057
rect 8880 17017 8892 17051
rect 8926 17017 8944 17051
rect 8880 17011 8944 17017
rect 8938 17008 8944 17011
rect 8996 17008 9002 17060
rect 5074 16980 5080 16992
rect 3896 16952 5080 16980
rect 3053 16943 3111 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 6135 16952 7021 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 7009 16949 7021 16952
rect 7055 16980 7067 16983
rect 7466 16980 7472 16992
rect 7055 16952 7472 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16980 7803 16983
rect 9508 16980 9536 17076
rect 12250 17048 12256 17060
rect 12211 17020 12256 17048
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 7791 16952 9536 16980
rect 7791 16949 7803 16952
rect 7745 16943 7803 16949
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 9824 16952 10793 16980
rect 9824 16940 9830 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 12342 16980 12348 16992
rect 12303 16952 12348 16980
rect 10781 16943 10839 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2314 16776 2320 16788
rect 2275 16748 2320 16776
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 2777 16779 2835 16785
rect 2777 16745 2789 16779
rect 2823 16745 2835 16779
rect 4062 16776 4068 16788
rect 4023 16748 4068 16776
rect 2777 16739 2835 16745
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 2130 16640 2136 16652
rect 1811 16612 2136 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2792 16640 2820 16739
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8389 16779 8447 16785
rect 8389 16776 8401 16779
rect 8352 16748 8401 16776
rect 8352 16736 8358 16748
rect 8389 16745 8401 16748
rect 8435 16745 8447 16779
rect 8389 16739 8447 16745
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10100 16748 10333 16776
rect 10100 16736 10106 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 12526 16776 12532 16788
rect 10321 16739 10379 16745
rect 10704 16748 12532 16776
rect 3145 16711 3203 16717
rect 3145 16677 3157 16711
rect 3191 16708 3203 16711
rect 4246 16708 4252 16720
rect 3191 16680 4252 16708
rect 3191 16677 3203 16680
rect 3145 16671 3203 16677
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 4798 16668 4804 16720
rect 4856 16708 4862 16720
rect 6264 16711 6322 16717
rect 4856 16680 5488 16708
rect 4856 16668 4862 16680
rect 2547 16612 2820 16640
rect 3237 16643 3295 16649
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 4154 16640 4160 16652
rect 3283 16612 4160 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 5460 16649 5488 16680
rect 6264 16677 6276 16711
rect 6310 16708 6322 16711
rect 6638 16708 6644 16720
rect 6310 16680 6644 16708
rect 6310 16677 6322 16680
rect 6264 16671 6322 16677
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 9861 16711 9919 16717
rect 9861 16677 9873 16711
rect 9907 16708 9919 16711
rect 10704 16708 10732 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 13630 16776 13636 16788
rect 13591 16748 13636 16776
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 10870 16717 10876 16720
rect 10864 16708 10876 16717
rect 9907 16680 10732 16708
rect 10831 16680 10876 16708
rect 9907 16677 9919 16680
rect 9861 16671 9919 16677
rect 10864 16671 10876 16680
rect 10870 16668 10876 16671
rect 10928 16668 10934 16720
rect 5178 16643 5236 16649
rect 5178 16640 5190 16643
rect 4396 16612 5190 16640
rect 4396 16600 4402 16612
rect 5178 16609 5190 16612
rect 5224 16609 5236 16643
rect 5178 16603 5236 16609
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5491 16612 6009 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 5997 16609 6009 16612
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 7524 16612 9229 16640
rect 7524 16600 7530 16612
rect 9217 16609 9229 16612
rect 9263 16640 9275 16643
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9263 16612 9965 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 12509 16643 12567 16649
rect 12509 16640 12521 16643
rect 9953 16603 10011 16609
rect 11992 16612 12521 16640
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 4062 16572 4068 16584
rect 3467 16544 4068 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 9582 16504 9588 16516
rect 9180 16476 9588 16504
rect 9180 16464 9186 16476
rect 9582 16464 9588 16476
rect 9640 16504 9646 16516
rect 10612 16504 10640 16535
rect 9640 16476 10640 16504
rect 9640 16464 9646 16476
rect 7374 16436 7380 16448
rect 7335 16408 7380 16436
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 11992 16445 12020 16612
rect 12509 16609 12521 16612
rect 12555 16609 12567 16643
rect 12509 16603 12567 16609
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 12216 16544 12265 16572
rect 12216 16532 12222 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 11977 16439 12035 16445
rect 11977 16436 11989 16439
rect 11756 16408 11989 16436
rect 11756 16396 11762 16408
rect 11977 16405 11989 16408
rect 12023 16405 12035 16439
rect 11977 16399 12035 16405
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 2133 16235 2191 16241
rect 2133 16232 2145 16235
rect 1820 16204 2145 16232
rect 1820 16192 1826 16204
rect 2133 16201 2145 16204
rect 2179 16201 2191 16235
rect 4338 16232 4344 16244
rect 4299 16204 4344 16232
rect 2133 16195 2191 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5074 16232 5080 16244
rect 5035 16204 5080 16232
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 1578 16164 1584 16176
rect 1539 16136 1584 16164
rect 1578 16124 1584 16136
rect 1636 16124 1642 16176
rect 6641 16167 6699 16173
rect 6641 16133 6653 16167
rect 6687 16133 6699 16167
rect 6641 16127 6699 16133
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4617 16099 4675 16105
rect 4617 16096 4629 16099
rect 4304 16068 4629 16096
rect 4304 16056 4310 16068
rect 4617 16065 4629 16068
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 16028 2375 16031
rect 2866 16028 2872 16040
rect 2363 16000 2872 16028
rect 2363 15997 2375 16000
rect 2317 15991 2375 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 4798 16028 4804 16040
rect 3007 16000 4804 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 5261 16031 5319 16037
rect 5261 15997 5273 16031
rect 5307 16028 5319 16031
rect 6656 16028 6684 16127
rect 7190 16096 7196 16108
rect 7151 16068 7196 16096
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 8938 16096 8944 16108
rect 8899 16068 8944 16096
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12250 16096 12256 16108
rect 12115 16068 12256 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 10134 16028 10140 16040
rect 5307 16000 6684 16028
rect 6748 16000 10140 16028
rect 5307 15997 5319 16000
rect 5261 15991 5319 15997
rect 1765 15963 1823 15969
rect 1765 15929 1777 15963
rect 1811 15960 1823 15963
rect 2590 15960 2596 15972
rect 1811 15932 2596 15960
rect 1811 15929 1823 15932
rect 1765 15923 1823 15929
rect 2590 15920 2596 15932
rect 2648 15920 2654 15972
rect 3228 15963 3286 15969
rect 3228 15929 3240 15963
rect 3274 15960 3286 15963
rect 3510 15960 3516 15972
rect 3274 15932 3516 15960
rect 3274 15929 3286 15932
rect 3228 15923 3286 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 5534 15960 5540 15972
rect 5447 15932 5540 15960
rect 5534 15920 5540 15932
rect 5592 15960 5598 15972
rect 6748 15960 6776 16000
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 5592 15932 6776 15960
rect 7009 15963 7067 15969
rect 5592 15920 5598 15932
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 7055 15932 7665 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 7653 15923 7711 15929
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2774 15892 2780 15904
rect 2731 15864 2780 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 2774 15852 2780 15864
rect 2832 15892 2838 15904
rect 3050 15892 3056 15904
rect 2832 15864 3056 15892
rect 2832 15852 2838 15864
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 7098 15852 7104 15904
rect 7156 15892 7162 15904
rect 8754 15892 8760 15904
rect 7156 15864 7201 15892
rect 8715 15864 8760 15892
rect 7156 15852 7162 15864
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 11790 15892 11796 15904
rect 8895 15864 11796 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2590 15688 2596 15700
rect 2551 15660 2596 15688
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 3053 15691 3111 15697
rect 3053 15688 3065 15691
rect 2746 15660 3065 15688
rect 1578 15620 1584 15632
rect 1539 15592 1584 15620
rect 1578 15580 1584 15592
rect 1636 15580 1642 15632
rect 2746 15620 2774 15660
rect 3053 15657 3065 15660
rect 3099 15657 3111 15691
rect 4154 15688 4160 15700
rect 4115 15660 4160 15688
rect 3053 15651 3111 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4525 15691 4583 15697
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 4798 15688 4804 15700
rect 4571 15660 4804 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 4798 15648 4804 15660
rect 4856 15688 4862 15700
rect 6181 15691 6239 15697
rect 6181 15688 6193 15691
rect 4856 15660 6193 15688
rect 4856 15648 4862 15660
rect 6181 15657 6193 15660
rect 6227 15688 6239 15691
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 6227 15660 8309 15688
rect 6227 15657 6239 15660
rect 6181 15651 6239 15657
rect 8297 15657 8309 15660
rect 8343 15688 8355 15691
rect 8754 15688 8760 15700
rect 8343 15660 8760 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8996 15660 9321 15688
rect 8996 15648 9002 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 12161 15691 12219 15697
rect 12161 15657 12173 15691
rect 12207 15688 12219 15691
rect 12342 15688 12348 15700
rect 12207 15660 12348 15688
rect 12207 15657 12219 15660
rect 12161 15651 12219 15657
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 2332 15592 2774 15620
rect 1762 15552 1768 15564
rect 1723 15524 1768 15552
rect 1762 15512 1768 15524
rect 1820 15512 1826 15564
rect 2332 15561 2360 15592
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 5534 15620 5540 15632
rect 4396 15592 4752 15620
rect 5495 15592 5540 15620
rect 4396 15580 4402 15592
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 3234 15552 3240 15564
rect 2832 15524 2877 15552
rect 3195 15524 3240 15552
rect 2832 15512 2838 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 4724 15493 4752 15592
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 7662 15623 7720 15629
rect 7662 15620 7674 15623
rect 7432 15592 7674 15620
rect 7432 15580 7438 15592
rect 7662 15589 7674 15592
rect 7708 15589 7720 15623
rect 9582 15620 9588 15632
rect 7662 15583 7720 15589
rect 9416 15592 9588 15620
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 8754 15552 8760 15564
rect 5675 15524 8760 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 5810 15484 5816 15496
rect 5771 15456 5816 15484
rect 4709 15447 4767 15453
rect 4632 15416 4660 15447
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8294 15484 8300 15496
rect 7975 15456 8300 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8294 15444 8300 15456
rect 8352 15484 8358 15496
rect 9416 15484 9444 15592
rect 9582 15580 9588 15592
rect 9640 15620 9646 15632
rect 9640 15592 10732 15620
rect 9640 15580 9646 15592
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10704 15561 10732 15592
rect 10422 15555 10480 15561
rect 10422 15552 10434 15555
rect 10008 15524 10434 15552
rect 10008 15512 10014 15524
rect 10422 15521 10434 15524
rect 10468 15521 10480 15555
rect 10422 15515 10480 15521
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15521 10747 15555
rect 11793 15555 11851 15561
rect 11793 15552 11805 15555
rect 10689 15515 10747 15521
rect 11072 15524 11805 15552
rect 8352 15456 9444 15484
rect 8352 15444 8358 15456
rect 5350 15416 5356 15428
rect 4632 15388 5356 15416
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 4212 15320 5181 15348
rect 4212 15308 4218 15320
rect 5169 15317 5181 15320
rect 5215 15317 5227 15351
rect 5169 15311 5227 15317
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 7190 15348 7196 15360
rect 6595 15320 7196 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 11072 15357 11100 15524
rect 11793 15521 11805 15524
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 11606 15484 11612 15496
rect 11567 15456 11612 15484
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15484 11759 15487
rect 12342 15484 12348 15496
rect 11747 15456 12348 15484
rect 11747 15453 11759 15456
rect 11701 15447 11759 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 7616 15320 11069 15348
rect 7616 15308 7622 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 2133 15147 2191 15153
rect 2133 15144 2145 15147
rect 1820 15116 2145 15144
rect 1820 15104 1826 15116
rect 2133 15113 2145 15116
rect 2179 15113 2191 15147
rect 2133 15107 2191 15113
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 2958 15144 2964 15156
rect 2915 15116 2964 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 4890 15144 4896 15156
rect 4396 15116 4896 15144
rect 4396 15104 4402 15116
rect 4890 15104 4896 15116
rect 4948 15144 4954 15156
rect 5442 15144 5448 15156
rect 4948 15116 5448 15144
rect 4948 15104 4954 15116
rect 5442 15104 5448 15116
rect 5500 15144 5506 15156
rect 5500 15116 6132 15144
rect 5500 15104 5506 15116
rect 4709 15079 4767 15085
rect 4709 15045 4721 15079
rect 4755 15045 4767 15079
rect 4709 15039 4767 15045
rect 3510 15017 3516 15020
rect 3467 15011 3516 15017
rect 3467 14977 3479 15011
rect 3513 14977 3516 15011
rect 3467 14971 3516 14977
rect 3510 14968 3516 14971
rect 3568 15008 3574 15020
rect 4724 15008 4752 15039
rect 6104 15017 6132 15116
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 7193 15147 7251 15153
rect 7193 15144 7205 15147
rect 7156 15116 7205 15144
rect 7156 15104 7162 15116
rect 7193 15113 7205 15116
rect 7239 15113 7251 15147
rect 7193 15107 7251 15113
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 8720 15116 8769 15144
rect 8720 15104 8726 15116
rect 8757 15113 8769 15116
rect 8803 15113 8815 15147
rect 8757 15107 8815 15113
rect 3568 14980 4752 15008
rect 6089 15011 6147 15017
rect 3568 14968 3574 14980
rect 6089 14977 6101 15011
rect 6135 14977 6147 15011
rect 6089 14971 6147 14977
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7098 15008 7104 15020
rect 6972 14980 7104 15008
rect 6972 14968 6978 14980
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7432 14980 7757 15008
rect 7432 14968 7438 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 9950 15008 9956 15020
rect 9447 14980 9956 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10410 15008 10416 15020
rect 10371 14980 10416 15008
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 3142 14940 3148 14952
rect 2363 14912 3148 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14940 3387 14943
rect 4154 14940 4160 14952
rect 3375 14912 4160 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 5810 14900 5816 14952
rect 5868 14949 5874 14952
rect 5868 14940 5880 14949
rect 5868 14912 5913 14940
rect 5868 14903 5880 14912
rect 5868 14900 5874 14903
rect 1765 14875 1823 14881
rect 1765 14841 1777 14875
rect 1811 14872 1823 14875
rect 2682 14872 2688 14884
rect 1811 14844 2688 14872
rect 1811 14841 1823 14844
rect 1765 14835 1823 14841
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14872 3295 14875
rect 3881 14875 3939 14881
rect 3881 14872 3893 14875
rect 3283 14844 3893 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 3881 14841 3893 14844
rect 3927 14841 3939 14875
rect 3881 14835 3939 14841
rect 10229 14875 10287 14881
rect 10229 14841 10241 14875
rect 10275 14872 10287 14875
rect 11146 14872 11152 14884
rect 10275 14844 11152 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4798 14804 4804 14816
rect 4479 14776 4804 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4798 14764 4804 14776
rect 4856 14804 4862 14816
rect 5258 14804 5264 14816
rect 4856 14776 5264 14804
rect 4856 14764 4862 14776
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 6914 14804 6920 14816
rect 6875 14776 6920 14804
rect 6914 14764 6920 14776
rect 6972 14804 6978 14816
rect 7558 14804 7564 14816
rect 6972 14776 7564 14804
rect 6972 14764 6978 14776
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 9122 14804 9128 14816
rect 7708 14776 7753 14804
rect 9083 14776 9128 14804
rect 7708 14764 7714 14776
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9263 14776 9781 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 10134 14804 10140 14816
rect 10047 14776 10140 14804
rect 9769 14767 9827 14773
rect 10134 14764 10140 14776
rect 10192 14804 10198 14816
rect 10778 14804 10784 14816
rect 10192 14776 10784 14804
rect 10192 14764 10198 14776
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2682 14600 2688 14612
rect 2643 14572 2688 14600
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 3142 14600 3148 14612
rect 3103 14572 3148 14600
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 5721 14603 5779 14609
rect 5721 14569 5733 14603
rect 5767 14600 5779 14603
rect 5810 14600 5816 14612
rect 5767 14572 5816 14600
rect 5767 14569 5779 14572
rect 5721 14563 5779 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9493 14603 9551 14609
rect 9493 14600 9505 14603
rect 9180 14572 9505 14600
rect 9180 14560 9186 14572
rect 9493 14569 9505 14572
rect 9539 14569 9551 14603
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9493 14563 9551 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 1765 14535 1823 14541
rect 1765 14501 1777 14535
rect 1811 14532 1823 14535
rect 2590 14532 2596 14544
rect 1811 14504 2596 14532
rect 1811 14501 1823 14504
rect 1765 14495 1823 14501
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 4890 14532 4896 14544
rect 3344 14504 4896 14532
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2188 14436 2329 14464
rect 2188 14424 2194 14436
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 2866 14464 2872 14476
rect 2827 14436 2872 14464
rect 2317 14427 2375 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3344 14473 3372 14504
rect 4890 14492 4896 14504
rect 4948 14492 4954 14544
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 8030 14535 8088 14541
rect 8030 14532 8042 14535
rect 7248 14504 8042 14532
rect 7248 14492 7254 14504
rect 8030 14501 8042 14504
rect 8076 14501 8088 14535
rect 8030 14495 8088 14501
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 10962 14532 10968 14544
rect 10468 14504 10968 14532
rect 10468 14492 10474 14504
rect 10962 14492 10968 14504
rect 11020 14532 11026 14544
rect 11066 14535 11124 14541
rect 11066 14532 11078 14535
rect 11020 14504 11078 14532
rect 11020 14492 11026 14504
rect 11066 14501 11078 14504
rect 11112 14501 11124 14535
rect 11066 14495 11124 14501
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4597 14467 4655 14473
rect 4597 14464 4609 14467
rect 4028 14436 4609 14464
rect 4028 14424 4034 14436
rect 4597 14433 4609 14436
rect 4643 14433 4655 14467
rect 4597 14427 4655 14433
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 11333 14467 11391 14473
rect 11333 14464 11345 14467
rect 9640 14436 11345 14464
rect 9640 14424 9646 14436
rect 11333 14433 11345 14436
rect 11379 14433 11391 14467
rect 11333 14427 11391 14433
rect 4338 14396 4344 14408
rect 4299 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 6914 14396 6920 14408
rect 6012 14368 6920 14396
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 6012 14337 6040 14368
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 5997 14331 6055 14337
rect 5997 14328 6009 14331
rect 5592 14300 6009 14328
rect 5592 14288 5598 14300
rect 5997 14297 6009 14300
rect 6043 14297 6055 14331
rect 5997 14291 6055 14297
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14260 4031 14263
rect 5626 14260 5632 14272
rect 4019 14232 5632 14260
rect 4019 14229 4031 14232
rect 3973 14223 4031 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6914 14260 6920 14272
rect 6875 14232 6920 14260
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2130 14056 2136 14068
rect 2091 14028 2136 14056
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3234 14056 3240 14068
rect 3007 14028 3240 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 8570 14056 8576 14068
rect 8531 14028 8576 14056
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 10962 14056 10968 14068
rect 10923 14028 10968 14056
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 1544 13892 2605 13920
rect 1544 13880 1550 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3988 13920 4016 14016
rect 8294 13988 8300 14000
rect 8255 13960 8300 13988
rect 8294 13948 8300 13960
rect 8352 13988 8358 14000
rect 8352 13960 9168 13988
rect 8352 13948 8358 13960
rect 3651 13892 4016 13920
rect 5353 13923 5411 13929
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5442 13920 5448 13932
rect 5399 13892 5448 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 6362 13920 6368 13932
rect 5500 13892 6368 13920
rect 5500 13880 5506 13892
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 8202 13920 8208 13932
rect 7699 13892 8208 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 3234 13852 3240 13864
rect 2363 13824 3240 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 4798 13852 4804 13864
rect 3467 13824 4804 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 6457 13855 6515 13861
rect 6457 13852 6469 13855
rect 5684 13824 6469 13852
rect 5684 13812 5690 13824
rect 6457 13821 6469 13824
rect 6503 13821 6515 13855
rect 6457 13815 6515 13821
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 8386 13852 8392 13864
rect 8159 13824 8392 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 1762 13784 1768 13796
rect 1723 13756 1768 13784
rect 1762 13744 1768 13756
rect 1820 13744 1826 13796
rect 5074 13744 5080 13796
rect 5132 13793 5138 13796
rect 5132 13784 5144 13793
rect 6472 13784 6500 13815
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 9140 13852 9168 13960
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9263 13892 9720 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9582 13852 9588 13864
rect 9140 13824 9588 13852
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9692 13852 9720 13892
rect 9858 13861 9864 13864
rect 9841 13855 9864 13861
rect 9841 13852 9853 13855
rect 9692 13824 9853 13852
rect 9841 13821 9853 13824
rect 9916 13852 9922 13864
rect 9916 13824 9989 13852
rect 9841 13815 9864 13821
rect 9858 13812 9864 13815
rect 9916 13812 9922 13824
rect 9214 13784 9220 13796
rect 5132 13756 5177 13784
rect 6472 13756 9220 13784
rect 5132 13747 5144 13756
rect 5132 13744 5138 13747
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 3326 13716 3332 13728
rect 3287 13688 3332 13716
rect 3326 13676 3332 13688
rect 3384 13676 3390 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 5994 13716 6000 13728
rect 5955 13688 6000 13716
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 7374 13716 7380 13728
rect 7335 13688 7380 13716
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 7469 13719 7527 13725
rect 7469 13685 7481 13719
rect 7515 13716 7527 13719
rect 7742 13716 7748 13728
rect 7515 13688 7748 13716
rect 7515 13685 7527 13688
rect 7469 13679 7527 13685
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 8938 13716 8944 13728
rect 8899 13688 8944 13716
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9088 13688 9133 13716
rect 9088 13676 9094 13688
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 1820 13484 2145 13512
rect 1820 13472 1826 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 2590 13512 2596 13524
rect 2551 13484 2596 13512
rect 2133 13475 2191 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 3384 13484 4537 13512
rect 3384 13472 3390 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 4525 13475 4583 13481
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 4985 13515 5043 13521
rect 4985 13512 4997 13515
rect 4856 13484 4997 13512
rect 4856 13472 4862 13484
rect 4985 13481 4997 13484
rect 5031 13481 5043 13515
rect 4985 13475 5043 13481
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5491 13484 8064 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 4120 13416 5764 13444
rect 4120 13404 4126 13416
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3237 13379 3295 13385
rect 2832 13348 2877 13376
rect 2832 13336 2838 13348
rect 3237 13345 3249 13379
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 3252 13308 3280 13339
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4028 13348 4261 13376
rect 4028 13336 4034 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5626 13376 5632 13388
rect 5399 13348 5632 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 5736 13376 5764 13416
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7162 13447 7220 13453
rect 7162 13444 7174 13447
rect 6972 13416 7174 13444
rect 6972 13404 6978 13416
rect 7162 13413 7174 13416
rect 7208 13413 7220 13447
rect 8036 13444 8064 13484
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 8260 13484 8309 13512
rect 8260 13472 8266 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 8297 13475 8355 13481
rect 8938 13472 8944 13524
rect 8996 13512 9002 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 8996 13484 9413 13512
rect 8996 13472 9002 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9858 13512 9864 13524
rect 9819 13484 9864 13512
rect 9401 13475 9459 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10042 13444 10048 13456
rect 8036 13416 10048 13444
rect 7162 13407 7220 13413
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 5994 13376 6000 13388
rect 5736 13348 6000 13376
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 8386 13376 8392 13388
rect 6687 13348 8392 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 10974 13379 11032 13385
rect 10974 13376 10986 13379
rect 10284 13348 10986 13376
rect 10284 13336 10290 13348
rect 10974 13345 10986 13348
rect 11020 13345 11032 13379
rect 11238 13376 11244 13388
rect 11151 13348 11244 13376
rect 10974 13339 11032 13345
rect 11238 13336 11244 13348
rect 11296 13376 11302 13388
rect 12158 13376 12164 13388
rect 11296 13348 12164 13376
rect 11296 13336 11302 13348
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 4338 13308 4344 13320
rect 3252 13280 4344 13308
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 8570 13308 8576 13320
rect 8531 13280 8576 13308
rect 6917 13271 6975 13277
rect 1578 13240 1584 13252
rect 1539 13212 1584 13240
rect 1578 13200 1584 13212
rect 1636 13200 1642 13252
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3292 13212 4077 13240
rect 3292 13200 3298 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 5074 13240 5080 13252
rect 4212 13212 5080 13240
rect 4212 13200 4218 13212
rect 5074 13200 5080 13212
rect 5132 13240 5138 13252
rect 5552 13240 5580 13271
rect 5132 13212 5580 13240
rect 5132 13200 5138 13212
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 6457 13243 6515 13249
rect 6457 13240 6469 13243
rect 6420 13212 6469 13240
rect 6420 13200 6426 13212
rect 6457 13209 6469 13212
rect 6503 13240 6515 13243
rect 6932 13240 6960 13271
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 6503 13212 6960 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 3050 13132 3056 13184
rect 3108 13172 3114 13184
rect 5994 13172 6000 13184
rect 3108 13144 6000 13172
rect 3108 13132 3114 13144
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1762 12968 1768 12980
rect 1723 12940 1768 12968
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 2498 12928 2504 12980
rect 2556 12928 2562 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3697 12971 3755 12977
rect 3697 12968 3709 12971
rect 2832 12940 3709 12968
rect 2832 12928 2838 12940
rect 3697 12937 3709 12940
rect 3743 12937 3755 12971
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 3697 12931 3755 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 7432 12940 7481 12968
rect 7432 12928 7438 12940
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 7742 12968 7748 12980
rect 7703 12940 7748 12968
rect 7469 12931 7527 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 9030 12928 9036 12980
rect 9088 12968 9094 12980
rect 9585 12971 9643 12977
rect 9585 12968 9597 12971
rect 9088 12940 9597 12968
rect 9088 12928 9094 12940
rect 9585 12937 9597 12940
rect 9631 12937 9643 12971
rect 9585 12931 9643 12937
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 2516 12841 2544 12928
rect 2961 12903 3019 12909
rect 2961 12869 2973 12903
rect 3007 12900 3019 12903
rect 4246 12900 4252 12912
rect 3007 12872 4252 12900
rect 3007 12869 3019 12872
rect 2961 12863 3019 12869
rect 4246 12860 4252 12872
rect 4304 12860 4310 12912
rect 5997 12903 6055 12909
rect 5997 12869 6009 12903
rect 6043 12900 6055 12903
rect 6043 12872 12434 12900
rect 6043 12869 6055 12872
rect 5997 12863 6055 12869
rect 2317 12835 2375 12841
rect 2317 12832 2329 12835
rect 1912 12804 2329 12832
rect 1912 12792 1918 12804
rect 2317 12801 2329 12804
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 5534 12832 5540 12844
rect 2648 12804 3924 12832
rect 5447 12804 5540 12832
rect 2648 12792 2654 12804
rect 3896 12773 3924 12804
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 6362 12832 6368 12844
rect 5592 12804 6368 12832
rect 5592 12792 5598 12804
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 6914 12832 6920 12844
rect 6875 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12832 6978 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 6972 12804 8309 12832
rect 6972 12792 6978 12804
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 9214 12832 9220 12844
rect 8996 12804 9220 12832
rect 8996 12792 9002 12804
rect 9214 12792 9220 12804
rect 9272 12832 9278 12844
rect 10226 12832 10232 12844
rect 9272 12804 9996 12832
rect 10187 12804 10232 12832
rect 9272 12792 9278 12804
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 3421 12767 3479 12773
rect 1995 12736 3372 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2314 12656 2320 12708
rect 2372 12696 2378 12708
rect 2372 12668 3280 12696
rect 2372 12656 2378 12668
rect 1394 12628 1400 12640
rect 1355 12600 1400 12628
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 2590 12628 2596 12640
rect 2551 12600 2596 12628
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 3252 12637 3280 12668
rect 3237 12631 3295 12637
rect 3237 12597 3249 12631
rect 3283 12597 3295 12631
rect 3344 12628 3372 12736
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 3436 12696 3464 12727
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 5776 12736 5825 12764
rect 5776 12724 5782 12736
rect 5813 12733 5825 12736
rect 5859 12733 5871 12767
rect 5813 12727 5871 12733
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 8570 12764 8576 12776
rect 7147 12736 8576 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9968 12773 9996 12804
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 4172 12696 4200 12724
rect 3436 12668 4200 12696
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5270 12699 5328 12705
rect 5270 12696 5282 12699
rect 5040 12668 5282 12696
rect 5040 12656 5046 12668
rect 5270 12665 5282 12668
rect 5316 12665 5328 12699
rect 5270 12659 5328 12665
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 8113 12699 8171 12705
rect 8113 12696 8125 12699
rect 6052 12668 8125 12696
rect 6052 12656 6058 12668
rect 8113 12665 8125 12668
rect 8159 12665 8171 12699
rect 8113 12659 8171 12665
rect 8205 12699 8263 12705
rect 8205 12665 8217 12699
rect 8251 12696 8263 12699
rect 8846 12696 8852 12708
rect 8251 12668 8852 12696
rect 8251 12665 8263 12668
rect 8205 12659 8263 12665
rect 5718 12628 5724 12640
rect 3344 12600 5724 12628
rect 3237 12591 3295 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6972 12600 7021 12628
rect 6972 12588 6978 12600
rect 7009 12597 7021 12600
rect 7055 12628 7067 12631
rect 7742 12628 7748 12640
rect 7055 12600 7748 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8128 12628 8156 12659
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 12406 12696 12434 12872
rect 19150 12696 19156 12708
rect 12406 12668 19156 12696
rect 19150 12656 19156 12668
rect 19208 12656 19214 12708
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8128 12600 8769 12628
rect 8757 12597 8769 12600
rect 8803 12628 8815 12631
rect 9858 12628 9864 12640
rect 8803 12600 9864 12628
rect 8803 12597 8815 12600
rect 8757 12591 8815 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10134 12628 10140 12640
rect 10091 12600 10140 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 2924 12396 4077 12424
rect 2924 12384 2930 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4982 12424 4988 12436
rect 4943 12396 4988 12424
rect 4065 12387 4123 12393
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 9861 12427 9919 12433
rect 5500 12396 8340 12424
rect 5500 12384 5506 12396
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 2970 12359 3028 12365
rect 2970 12356 2982 12359
rect 2832 12328 2982 12356
rect 2832 12316 2838 12328
rect 2970 12325 2982 12328
rect 3016 12325 3028 12359
rect 2970 12319 3028 12325
rect 3878 12316 3884 12368
rect 3936 12356 3942 12368
rect 5810 12356 5816 12368
rect 3936 12328 5816 12356
rect 3936 12316 3942 12328
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 6178 12316 6184 12368
rect 6236 12316 6242 12368
rect 7000 12359 7058 12365
rect 7000 12325 7012 12359
rect 7046 12356 7058 12359
rect 8202 12356 8208 12368
rect 7046 12328 8208 12356
rect 7046 12325 7058 12328
rect 7000 12319 7058 12325
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8312 12365 8340 12396
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 10226 12424 10232 12436
rect 9907 12396 10232 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12325 8355 12359
rect 8297 12319 8355 12325
rect 8404 12328 12434 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1486 12288 1492 12300
rect 1443 12260 1492 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 4246 12288 4252 12300
rect 4207 12260 4252 12288
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 5626 12288 5632 12300
rect 4356 12260 5632 12288
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 4356 12220 4384 12260
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 6086 12288 6092 12300
rect 6144 12297 6150 12300
rect 6056 12260 6092 12288
rect 6086 12248 6092 12260
rect 6144 12251 6156 12297
rect 6196 12288 6224 12316
rect 8404 12288 8432 12328
rect 8570 12288 8576 12300
rect 6196 12260 8432 12288
rect 8531 12260 8576 12288
rect 6144 12248 6150 12251
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 10974 12291 11032 12297
rect 10974 12288 10986 12291
rect 10652 12260 10986 12288
rect 10652 12248 10658 12260
rect 10974 12257 10986 12260
rect 11020 12257 11032 12291
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 10974 12251 11032 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 12406 12288 12434 12328
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 12406 12260 19809 12288
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 3283 12192 4384 12220
rect 4709 12223 4767 12229
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4890 12220 4896 12232
rect 4755 12192 4896 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 1670 12084 1676 12096
rect 1627 12056 1676 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3252 12084 3280 12183
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6730 12220 6736 12232
rect 6420 12192 6736 12220
rect 6420 12180 6426 12192
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8343 12192 9137 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 8036 12124 10364 12152
rect 2924 12056 3280 12084
rect 2924 12044 2930 12056
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 8036 12084 8064 12124
rect 3936 12056 8064 12084
rect 8113 12087 8171 12093
rect 3936 12044 3942 12056
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8202 12084 8208 12096
rect 8159 12056 8208 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8386 12084 8392 12096
rect 8347 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 10336 12084 10364 12124
rect 11698 12084 11704 12096
rect 10336 12056 11704 12084
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20806 12084 20812 12096
rect 20027 12056 20812 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20806 12044 20812 12056
rect 20864 12044 20870 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2648 11852 2697 11880
rect 2648 11840 2654 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 2685 11843 2743 11849
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3200 11852 4292 11880
rect 3200 11840 3206 11852
rect 4264 11812 4292 11852
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 4396 11852 4629 11880
rect 4396 11840 4402 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7098 11880 7104 11892
rect 7055 11852 7104 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 9950 11880 9956 11892
rect 9911 11852 9956 11880
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 12066 11880 12072 11892
rect 11296 11852 12072 11880
rect 11296 11840 11302 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 6546 11812 6552 11824
rect 4264 11784 6552 11812
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11744 2191 11747
rect 2774 11744 2780 11756
rect 2179 11716 2780 11744
rect 2179 11713 2191 11716
rect 2133 11707 2191 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 2866 11704 2872 11756
rect 2924 11744 2930 11756
rect 2968 11747 3026 11753
rect 2968 11744 2980 11747
rect 2924 11716 2980 11744
rect 2924 11704 2930 11716
rect 2968 11713 2980 11716
rect 3014 11713 3026 11747
rect 2968 11707 3026 11713
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 5040 11716 5181 11744
rect 5040 11704 5046 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 10594 11744 10600 11756
rect 7699 11716 8432 11744
rect 10555 11716 10600 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 1489 11679 1547 11685
rect 1489 11645 1501 11679
rect 1535 11676 1547 11679
rect 1578 11676 1584 11688
rect 1535 11648 1584 11676
rect 1535 11645 1547 11648
rect 1489 11639 1547 11645
rect 1578 11636 1584 11648
rect 1636 11676 1642 11688
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 1636 11648 5641 11676
rect 1636 11636 1642 11648
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 8294 11676 8300 11688
rect 8255 11648 8300 11676
rect 5629 11639 5687 11645
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8404 11676 8432 11716
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 8553 11679 8611 11685
rect 8553 11676 8565 11679
rect 8404 11648 8565 11676
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 3206 11611 3264 11617
rect 3206 11608 3218 11611
rect 1912 11580 3218 11608
rect 1912 11568 1918 11580
rect 3206 11577 3218 11580
rect 3252 11577 3264 11611
rect 3206 11571 3264 11577
rect 4890 11568 4896 11620
rect 4948 11608 4954 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 4948 11580 4997 11608
rect 4948 11568 4954 11580
rect 4985 11577 4997 11580
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 6457 11611 6515 11617
rect 6457 11608 6469 11611
rect 5960 11580 6469 11608
rect 5960 11568 5966 11580
rect 6457 11577 6469 11580
rect 6503 11577 6515 11611
rect 6457 11571 6515 11577
rect 8496 11552 8524 11648
rect 8553 11645 8565 11648
rect 8599 11645 8611 11679
rect 8553 11639 8611 11645
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10778 11676 10784 11688
rect 9916 11648 10784 11676
rect 9916 11636 9922 11648
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 10928 11648 11897 11676
rect 10928 11636 10934 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 19150 11676 19156 11688
rect 19111 11648 19156 11676
rect 11885 11639 11943 11645
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 10321 11611 10379 11617
rect 10321 11577 10333 11611
rect 10367 11608 10379 11611
rect 10965 11611 11023 11617
rect 10965 11608 10977 11611
rect 10367 11580 10977 11608
rect 10367 11577 10379 11580
rect 10321 11571 10379 11577
rect 10965 11577 10977 11580
rect 11011 11577 11023 11611
rect 10965 11571 11023 11577
rect 1673 11543 1731 11549
rect 1673 11509 1685 11543
rect 1719 11540 1731 11543
rect 2038 11540 2044 11552
rect 1719 11512 2044 11540
rect 1719 11509 1731 11512
rect 1673 11503 1731 11509
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 4338 11540 4344 11552
rect 2372 11512 2417 11540
rect 4299 11512 4344 11540
rect 2372 11500 2378 11512
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5534 11540 5540 11552
rect 5123 11512 5540 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5994 11540 6000 11552
rect 5955 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6880 11512 7389 11540
rect 6880 11500 6886 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7524 11512 7569 11540
rect 7524 11500 7530 11512
rect 8478 11500 8484 11552
rect 8536 11500 8542 11552
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 9766 11540 9772 11552
rect 9723 11512 9772 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 19334 11540 19340 11552
rect 19295 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2130 11336 2136 11348
rect 1627 11308 2136 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 2314 11336 2320 11348
rect 2271 11308 2320 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2685 11339 2743 11345
rect 2685 11336 2697 11339
rect 2556 11308 2697 11336
rect 2556 11296 2562 11308
rect 2685 11305 2697 11308
rect 2731 11305 2743 11339
rect 3142 11336 3148 11348
rect 3103 11308 3148 11336
rect 2685 11299 2743 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5626 11336 5632 11348
rect 4672 11308 5632 11336
rect 4672 11296 4678 11308
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 5997 11339 6055 11345
rect 5997 11305 6009 11339
rect 6043 11336 6055 11339
rect 6086 11336 6092 11348
rect 6043 11308 6092 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10652 11308 10885 11336
rect 10652 11296 10658 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 3878 11268 3884 11280
rect 2096 11240 3884 11268
rect 2096 11228 2102 11240
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 6273 11271 6331 11277
rect 6273 11268 6285 11271
rect 4080 11240 6285 11268
rect 4080 11212 4108 11240
rect 6273 11237 6285 11240
rect 6319 11237 6331 11271
rect 6273 11231 6331 11237
rect 7368 11271 7426 11277
rect 7368 11237 7380 11271
rect 7414 11268 7426 11271
rect 8202 11268 8208 11280
rect 7414 11240 8208 11268
rect 7414 11237 7426 11240
rect 7368 11231 7426 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 8444 11240 12434 11268
rect 8444 11228 8450 11240
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 3050 11200 3056 11212
rect 2963 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11200 3114 11212
rect 3602 11200 3608 11212
rect 3108 11172 3608 11200
rect 3108 11160 3114 11172
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4890 11209 4896 11212
rect 4884 11163 4896 11209
rect 4948 11200 4954 11212
rect 4948 11172 4984 11200
rect 4890 11160 4896 11163
rect 4948 11160 4954 11172
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6788 11172 7113 11200
rect 6788 11160 6794 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 9766 11209 9772 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8352 11172 9505 11200
rect 8352 11160 8358 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9760 11200 9772 11209
rect 9679 11172 9772 11200
rect 9493 11163 9551 11169
rect 9760 11163 9772 11172
rect 9824 11200 9830 11212
rect 10594 11200 10600 11212
rect 9824 11172 10600 11200
rect 9766 11160 9772 11163
rect 9824 11160 9830 11172
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 12406 11200 12434 11240
rect 18693 11203 18751 11209
rect 18693 11200 18705 11203
rect 12406 11172 18705 11200
rect 18693 11169 18705 11172
rect 18739 11169 18751 11203
rect 18693 11163 18751 11169
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 4614 11132 4620 11144
rect 3292 11104 3337 11132
rect 4575 11104 4620 11132
rect 3292 11092 3298 11104
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 1486 11024 1492 11076
rect 1544 11064 1550 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1544 11036 1869 11064
rect 1544 11024 1550 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 9122 11064 9128 11076
rect 9083 11036 9128 11064
rect 1857 11027 1915 11033
rect 9122 11024 9128 11036
rect 9180 11024 9186 11076
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 10836 11036 11161 11064
rect 10836 11024 10842 11036
rect 11149 11033 11161 11036
rect 11195 11033 11207 11067
rect 11149 11027 11207 11033
rect 18877 11067 18935 11073
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 19886 11064 19892 11076
rect 18923 11036 19892 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 11974 10996 11980 11008
rect 1728 10968 11980 10996
rect 1728 10956 1734 10968
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2832 10764 3065 10792
rect 2832 10752 2838 10764
rect 3053 10761 3065 10764
rect 3099 10792 3111 10795
rect 3234 10792 3240 10804
rect 3099 10764 3240 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3329 10795 3387 10801
rect 3329 10761 3341 10795
rect 3375 10792 3387 10795
rect 4798 10792 4804 10804
rect 3375 10764 4804 10792
rect 3375 10761 3387 10764
rect 3329 10755 3387 10761
rect 4798 10752 4804 10764
rect 4856 10792 4862 10804
rect 4856 10764 5028 10792
rect 4856 10752 4862 10764
rect 5000 10724 5028 10764
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5442 10792 5448 10804
rect 5132 10764 5448 10792
rect 5132 10752 5138 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 5776 10764 6837 10792
rect 5776 10752 5782 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7466 10792 7472 10804
rect 7423 10764 7472 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10410 10792 10416 10804
rect 10091 10764 10416 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 9490 10724 9496 10736
rect 5000 10696 5304 10724
rect 2746 10628 4108 10656
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2746 10588 2774 10628
rect 4080 10600 4108 10628
rect 1719 10560 2774 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 3513 10591 3571 10597
rect 3513 10588 3525 10591
rect 3292 10560 3525 10588
rect 3292 10548 3298 10560
rect 3513 10557 3525 10560
rect 3559 10557 3571 10591
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 3513 10551 3571 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4338 10597 4344 10600
rect 4332 10588 4344 10597
rect 4299 10560 4344 10588
rect 4332 10551 4344 10560
rect 4396 10588 4402 10600
rect 5166 10588 5172 10600
rect 4396 10560 5172 10588
rect 4338 10548 4344 10551
rect 4396 10548 4402 10560
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5276 10588 5304 10696
rect 7944 10696 9496 10724
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 7944 10656 7972 10696
rect 9490 10684 9496 10696
rect 9548 10724 9554 10736
rect 9548 10696 9720 10724
rect 9548 10684 9554 10696
rect 5500 10628 7972 10656
rect 8021 10659 8079 10665
rect 5500 10616 5506 10628
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8202 10656 8208 10668
rect 8067 10628 8208 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9364 10628 9597 10656
rect 9364 10616 9370 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9692 10656 9720 10696
rect 9766 10684 9772 10736
rect 9824 10724 9830 10736
rect 10962 10724 10968 10736
rect 9824 10696 10968 10724
rect 9824 10684 9830 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 10410 10656 10416 10668
rect 9692 10628 10416 10656
rect 9585 10619 9643 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 5626 10588 5632 10600
rect 5276 10560 5632 10588
rect 5626 10548 5632 10560
rect 5684 10588 5690 10600
rect 7006 10588 7012 10600
rect 5684 10560 6592 10588
rect 6967 10560 7012 10588
rect 5684 10548 5690 10560
rect 1946 10529 1952 10532
rect 1940 10520 1952 10529
rect 1907 10492 1952 10520
rect 1940 10483 1952 10492
rect 1946 10480 1952 10483
rect 2004 10480 2010 10532
rect 6457 10523 6515 10529
rect 6457 10520 6469 10523
rect 4448 10492 6469 10520
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 4448 10452 4476 10492
rect 6457 10489 6469 10492
rect 6503 10489 6515 10523
rect 6564 10520 6592 10560
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 8803 10560 11897 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 7745 10523 7803 10529
rect 7745 10520 7757 10523
rect 6564 10492 7757 10520
rect 6457 10483 6515 10489
rect 7745 10489 7757 10492
rect 7791 10489 7803 10523
rect 7745 10483 7803 10489
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 7883 10492 9812 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 3384 10424 4476 10452
rect 3384 10412 3390 10424
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 4948 10424 5457 10452
rect 4948 10412 4954 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5445 10415 5503 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9398 10452 9404 10464
rect 9359 10424 9404 10452
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9674 10452 9680 10464
rect 9539 10424 9680 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9784 10452 9812 10492
rect 9858 10480 9864 10532
rect 9916 10520 9922 10532
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9916 10492 10517 10520
rect 9916 10480 9922 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 11900 10520 11928 10551
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 18233 10591 18291 10597
rect 18233 10588 18245 10591
rect 12032 10560 18245 10588
rect 12032 10548 12038 10560
rect 18233 10557 18245 10560
rect 18279 10588 18291 10591
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18279 10560 18705 10588
rect 18279 10557 18291 10560
rect 18233 10551 18291 10557
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 12894 10520 12900 10532
rect 11900 10492 12900 10520
rect 10505 10483 10563 10489
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 13630 10520 13636 10532
rect 13591 10492 13636 10520
rect 13630 10480 13636 10492
rect 13688 10480 13694 10532
rect 10226 10452 10232 10464
rect 9784 10424 10232 10452
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 11054 10452 11060 10464
rect 11015 10424 11060 10452
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 19426 10452 19432 10464
rect 18463 10424 19432 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 7006 10248 7012 10260
rect 2087 10220 6868 10248
rect 6967 10220 7012 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 3878 10180 3884 10192
rect 1872 10152 3884 10180
rect 1872 10124 1900 10152
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 4985 10183 5043 10189
rect 4985 10180 4997 10183
rect 4856 10152 4997 10180
rect 4856 10140 4862 10152
rect 4985 10149 4997 10152
rect 5031 10149 5043 10183
rect 4985 10143 5043 10149
rect 5077 10183 5135 10189
rect 5077 10149 5089 10183
rect 5123 10180 5135 10183
rect 5123 10152 5396 10180
rect 5123 10149 5135 10152
rect 5077 10143 5135 10149
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2498 10112 2504 10124
rect 2424 10084 2504 10112
rect 2424 10053 2452 10084
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 3326 10112 3332 10124
rect 3287 10084 3332 10112
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5224 10084 5313 10112
rect 5224 10072 5230 10084
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10013 2467 10047
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2409 10007 2467 10013
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 5285 10053 5313 10084
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5368 10044 5396 10152
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 5997 10183 6055 10189
rect 5997 10180 6009 10183
rect 5500 10152 6009 10180
rect 5500 10140 5506 10152
rect 5997 10149 6009 10152
rect 6043 10149 6055 10183
rect 6840 10180 6868 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7374 10248 7380 10260
rect 7156 10220 7380 10248
rect 7156 10208 7162 10220
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 9030 10248 9036 10260
rect 7515 10220 9036 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 9720 10248
rect 9548 10208 9554 10220
rect 9582 10180 9588 10192
rect 6840 10152 9588 10180
rect 5997 10143 6055 10149
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 9692 10180 9720 10220
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 9824 10220 9869 10248
rect 9824 10208 9830 10220
rect 9861 10183 9919 10189
rect 9861 10180 9873 10183
rect 9692 10152 9873 10180
rect 9861 10149 9873 10152
rect 9907 10149 9919 10183
rect 11054 10180 11060 10192
rect 9861 10143 9919 10149
rect 10244 10152 11060 10180
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6730 10112 6736 10124
rect 6135 10084 6736 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 8389 10115 8447 10121
rect 8389 10112 8401 10115
rect 7800 10084 8401 10112
rect 7800 10072 7806 10084
rect 8389 10081 8401 10084
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 9214 10112 9220 10124
rect 8527 10084 9220 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 9214 10072 9220 10084
rect 9272 10112 9278 10124
rect 10244 10112 10272 10152
rect 11054 10140 11060 10152
rect 11112 10180 11118 10192
rect 13538 10180 13544 10192
rect 11112 10152 13544 10180
rect 11112 10140 11118 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 9272 10084 10272 10112
rect 10321 10115 10379 10121
rect 9272 10072 9278 10084
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10367 10084 10793 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10781 10081 10793 10084
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 12825 10115 12883 10121
rect 12825 10081 12837 10115
rect 12871 10112 12883 10115
rect 13262 10112 13268 10124
rect 12871 10084 13268 10112
rect 12871 10081 12883 10084
rect 12825 10075 12883 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 5368 10016 6141 10044
rect 5261 10007 5319 10013
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9976 1639 9979
rect 5442 9976 5448 9988
rect 1627 9948 5448 9976
rect 1627 9945 1639 9948
rect 1581 9939 1639 9945
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 5592 9948 5641 9976
rect 5592 9936 5598 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 6113 9976 6141 10016
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 7561 10047 7619 10053
rect 6236 10016 6281 10044
rect 6236 10004 6242 10016
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 7466 9976 7472 9988
rect 6113 9948 7472 9976
rect 5629 9939 5687 9945
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 3418 9908 3424 9920
rect 3099 9880 3424 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 4617 9911 4675 9917
rect 3568 9880 3613 9908
rect 3568 9868 3574 9880
rect 4617 9877 4629 9911
rect 4663 9908 4675 9911
rect 4798 9908 4804 9920
rect 4663 9880 4804 9908
rect 4663 9877 4675 9880
rect 4617 9871 4675 9877
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 7576 9908 7604 10007
rect 8680 9976 8708 10007
rect 8938 10004 8944 10056
rect 8996 10044 9002 10056
rect 9582 10044 9588 10056
rect 8996 10016 9588 10044
rect 8996 10004 9002 10016
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 9968 9976 9996 10007
rect 10502 9976 10508 9988
rect 8680 9948 10508 9976
rect 10502 9936 10508 9948
rect 10560 9976 10566 9988
rect 11701 9979 11759 9985
rect 11701 9976 11713 9979
rect 10560 9948 11713 9976
rect 10560 9936 10566 9948
rect 11701 9945 11713 9948
rect 11747 9945 11759 9979
rect 11701 9939 11759 9945
rect 7650 9908 7656 9920
rect 6696 9880 6741 9908
rect 7576 9880 7656 9908
rect 6696 9868 6702 9880
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 8021 9911 8079 9917
rect 8021 9877 8033 9911
rect 8067 9908 8079 9911
rect 8386 9908 8392 9920
rect 8067 9880 8392 9908
rect 8067 9877 8079 9880
rect 8021 9871 8079 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9858 9908 9864 9920
rect 8536 9880 9864 9908
rect 8536 9868 8542 9880
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10008 9880 10333 9908
rect 10008 9868 10014 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 10321 9871 10379 9877
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10594 9908 10600 9920
rect 10459 9880 10600 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 11112 9880 11161 9908
rect 11112 9868 11118 9880
rect 11149 9877 11161 9880
rect 11195 9877 11207 9911
rect 11149 9871 11207 9877
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12066 9908 12072 9920
rect 11940 9880 12072 9908
rect 11940 9868 11946 9880
rect 12066 9868 12072 9880
rect 12124 9908 12130 9920
rect 13096 9908 13124 10007
rect 12124 9880 13124 9908
rect 12124 9868 12130 9880
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 3142 9704 3148 9716
rect 2648 9676 3148 9704
rect 2648 9664 2654 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3292 9676 5396 9704
rect 3292 9664 3298 9676
rect 3970 9636 3976 9648
rect 2976 9608 3464 9636
rect 3931 9608 3976 9636
rect 2976 9577 3004 9608
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3436 9568 3464 9608
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 4249 9639 4307 9645
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 4982 9636 4988 9648
rect 4295 9608 4988 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5368 9636 5396 9676
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 13538 9704 13544 9716
rect 5500 9676 13400 9704
rect 13499 9676 13544 9704
rect 5500 9664 5506 9676
rect 5994 9636 6000 9648
rect 5368 9608 6000 9636
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6825 9639 6883 9645
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 6871 9608 7236 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 4706 9568 4712 9580
rect 3436 9540 4108 9568
rect 4667 9540 4712 9568
rect 3329 9531 3387 9537
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 2694 9435 2752 9441
rect 2694 9432 2706 9435
rect 2648 9404 2706 9432
rect 2648 9392 2654 9404
rect 2694 9401 2706 9404
rect 2740 9401 2752 9435
rect 2694 9395 2752 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1946 9364 1952 9376
rect 1627 9336 1952 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1946 9324 1952 9336
rect 2004 9364 2010 9376
rect 3344 9364 3372 9531
rect 4080 9512 4108 9540
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4890 9568 4896 9580
rect 4851 9540 4896 9568
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3476 9472 3617 9500
rect 3476 9460 3482 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4246 9500 4252 9512
rect 4120 9472 4252 9500
rect 4120 9460 4126 9472
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4396 9472 4629 9500
rect 4396 9460 4402 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 6086 9500 6092 9512
rect 6047 9472 6092 9500
rect 4617 9463 4675 9469
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 7208 9500 7236 9608
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 9306 9636 9312 9648
rect 8352 9608 8524 9636
rect 9267 9608 9312 9636
rect 8352 9596 8358 9608
rect 8496 9577 8524 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 10965 9639 11023 9645
rect 10965 9636 10977 9639
rect 10928 9608 10977 9636
rect 10928 9596 10934 9608
rect 10965 9605 10977 9608
rect 11011 9605 11023 9639
rect 13372 9636 13400 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 15838 9704 15844 9716
rect 13648 9676 15844 9704
rect 13648 9636 13676 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 13372 9608 13676 9636
rect 10965 9599 11023 9605
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8938 9568 8944 9580
rect 8899 9540 8944 9568
rect 8481 9531 8539 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 11164 9540 12020 9568
rect 7650 9500 7656 9512
rect 7208 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8202 9500 8208 9512
rect 8163 9472 8208 9500
rect 8202 9460 8208 9472
rect 8260 9500 8266 9512
rect 11164 9509 11192 9540
rect 10689 9503 10747 9509
rect 10689 9500 10701 9503
rect 8260 9472 10701 9500
rect 8260 9460 8266 9472
rect 10689 9469 10701 9472
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11882 9500 11888 9512
rect 11843 9472 11888 9500
rect 11149 9463 11207 9469
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 11992 9500 12020 9540
rect 13078 9500 13084 9512
rect 11992 9472 13084 9500
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 4028 9404 6469 9432
rect 4028 9392 4034 9404
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 7960 9435 8018 9441
rect 7960 9401 7972 9435
rect 8006 9432 8018 9435
rect 9306 9432 9312 9444
rect 8006 9404 9312 9432
rect 8006 9401 8018 9404
rect 7960 9395 8018 9401
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9582 9392 9588 9444
rect 9640 9432 9646 9444
rect 9950 9432 9956 9444
rect 9640 9404 9956 9432
rect 9640 9392 9646 9404
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10502 9441 10508 9444
rect 10444 9435 10508 9441
rect 10444 9401 10456 9435
rect 10490 9401 10508 9435
rect 10444 9395 10508 9401
rect 10502 9392 10508 9395
rect 10560 9392 10566 9444
rect 11238 9392 11244 9444
rect 11296 9432 11302 9444
rect 12130 9435 12188 9441
rect 12130 9432 12142 9435
rect 11296 9404 12142 9432
rect 11296 9392 11302 9404
rect 12130 9401 12142 9404
rect 12176 9432 12188 9435
rect 14550 9432 14556 9444
rect 12176 9404 14556 9432
rect 12176 9401 12188 9404
rect 12130 9395 12188 9401
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 3510 9364 3516 9376
rect 2004 9336 3372 9364
rect 3471 9336 3516 9364
rect 2004 9324 2010 9336
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4856 9336 5457 9364
rect 4856 9324 4862 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5592 9336 5917 9364
rect 5592 9324 5598 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 10962 9364 10968 9376
rect 6052 9336 10968 9364
rect 6052 9324 6058 9336
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 12986 9364 12992 9376
rect 11480 9336 12992 9364
rect 11480 9324 11486 9336
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 2682 9160 2688 9172
rect 2179 9132 2688 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 3510 9160 3516 9172
rect 3191 9132 3516 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4798 9160 4804 9172
rect 4759 9132 4804 9160
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6328 9132 7328 9160
rect 6328 9120 6334 9132
rect 3421 9095 3479 9101
rect 3421 9092 3433 9095
rect 1412 9064 3433 9092
rect 1412 9036 1440 9064
rect 3421 9061 3433 9064
rect 3467 9061 3479 9095
rect 5994 9092 6000 9104
rect 3421 9055 3479 9061
rect 3528 9064 6000 9092
rect 3528 9036 3556 9064
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 7300 9092 7328 9132
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7432 9132 7941 9160
rect 7432 9120 7438 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 7929 9123 7987 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9674 9160 9680 9172
rect 8444 9132 8489 9160
rect 9635 9132 9680 9160
rect 8444 9120 8450 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11698 9160 11704 9172
rect 11471 9132 11704 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 11839 9132 12357 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13044 9132 13553 9160
rect 13044 9120 13050 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 14550 9160 14556 9172
rect 14511 9132 14556 9160
rect 13541 9123 13599 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 9398 9092 9404 9104
rect 6144 9064 7236 9092
rect 7300 9064 9404 9092
rect 6144 9052 6150 9064
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 3510 8984 3516 9036
rect 3568 8984 3574 9036
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 4396 8996 5856 9024
rect 4396 8984 4402 8996
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2866 8956 2872 8968
rect 2731 8928 2872 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 3200 8928 4905 8956
rect 3200 8916 3206 8928
rect 4893 8925 4905 8928
rect 4939 8956 4951 8959
rect 4982 8956 4988 8968
rect 4939 8928 4988 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5123 8928 5488 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5258 8888 5264 8900
rect 2700 8860 5264 8888
rect 2700 8832 2728 8860
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2038 8820 2044 8832
rect 1627 8792 2044 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2682 8780 2688 8832
rect 2740 8780 2746 8832
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4798 8820 4804 8832
rect 4479 8792 4804 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5460 8829 5488 8928
rect 5445 8823 5503 8829
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 5718 8820 5724 8832
rect 5491 8792 5724 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5828 8820 5856 8996
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6558 9027 6616 9033
rect 6558 9024 6570 9027
rect 6236 8996 6570 9024
rect 6236 8984 6242 8996
rect 6558 8993 6570 8996
rect 6604 8993 6616 9027
rect 7208 9024 7236 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 10137 9095 10195 9101
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 12158 9092 12164 9104
rect 10183 9064 12164 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 7208 8996 7297 9024
rect 6558 8987 6616 8993
rect 7285 8993 7297 8996
rect 7331 9024 7343 9027
rect 9122 9024 9128 9036
rect 7331 8996 9128 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10778 9024 10784 9036
rect 10091 8996 10784 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 9024 12495 9027
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 12483 8996 13093 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 15286 8984 15292 9036
rect 15344 9024 15350 9036
rect 15666 9027 15724 9033
rect 15666 9024 15678 9027
rect 15344 8996 15678 9024
rect 15344 8984 15350 8996
rect 15666 8993 15678 8996
rect 15712 8993 15724 9027
rect 15666 8987 15724 8993
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6871 8928 6929 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 8294 8956 8300 8968
rect 7524 8928 8300 8956
rect 7524 8916 7530 8928
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9306 8956 9312 8968
rect 8619 8928 9312 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8956 10287 8959
rect 10502 8956 10508 8968
rect 10275 8928 10508 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 11238 8956 11244 8968
rect 11199 8928 11244 8956
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8956 11391 8959
rect 12066 8956 12072 8968
rect 11379 8928 12072 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8956 12311 8959
rect 13262 8956 13268 8968
rect 12299 8928 13268 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8925 15991 8959
rect 15933 8919 15991 8925
rect 7561 8891 7619 8897
rect 7561 8888 7573 8891
rect 6840 8860 7573 8888
rect 6840 8820 6868 8860
rect 7561 8857 7573 8860
rect 7607 8857 7619 8891
rect 11422 8888 11428 8900
rect 7561 8851 7619 8857
rect 7668 8860 11428 8888
rect 5828 8792 6868 8820
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 6972 8792 7113 8820
rect 6972 8780 6978 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 7101 8783 7159 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7668 8820 7696 8860
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 7432 8792 7696 8820
rect 7432 8780 7438 8792
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8720 8792 9137 8820
rect 8720 8780 8726 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9214 8780 9220 8832
rect 9272 8820 9278 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 9272 8792 10701 8820
rect 9272 8780 9278 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 12805 8823 12863 8829
rect 12805 8789 12817 8823
rect 12851 8820 12863 8823
rect 13538 8820 13544 8832
rect 12851 8792 13544 8820
rect 12851 8789 12863 8792
rect 12805 8783 12863 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 14001 8823 14059 8829
rect 14001 8789 14013 8823
rect 14047 8820 14059 8823
rect 14090 8820 14096 8832
rect 14047 8792 14096 8820
rect 14047 8789 14059 8792
rect 14001 8783 14059 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 15948 8820 15976 8919
rect 15620 8792 15976 8820
rect 15620 8780 15626 8792
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 3510 8616 3516 8628
rect 1627 8588 3516 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 8665 8619 8723 8625
rect 3835 8588 8616 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 3329 8551 3387 8557
rect 3329 8517 3341 8551
rect 3375 8517 3387 8551
rect 3329 8511 3387 8517
rect 5721 8551 5779 8557
rect 5721 8517 5733 8551
rect 5767 8548 5779 8551
rect 5810 8548 5816 8560
rect 5767 8520 5816 8548
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 1964 8276 1992 8375
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 3344 8412 3372 8511
rect 5810 8508 5816 8520
rect 5868 8508 5874 8560
rect 8588 8548 8616 8588
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8754 8616 8760 8628
rect 8711 8588 8760 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 9548 8588 10609 8616
rect 9548 8576 9554 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 13078 8616 13084 8628
rect 13039 8588 13084 8616
rect 10597 8579 10655 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 11882 8548 11888 8560
rect 8588 8520 11888 8548
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 12621 8551 12679 8557
rect 12621 8517 12633 8551
rect 12667 8548 12679 8551
rect 13354 8548 13360 8560
rect 12667 8520 13360 8548
rect 12667 8517 12679 8520
rect 12621 8511 12679 8517
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 14829 8551 14887 8557
rect 14829 8517 14841 8551
rect 14875 8548 14887 8551
rect 17313 8551 17371 8557
rect 14875 8520 15332 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 15304 8492 15332 8520
rect 17313 8517 17325 8551
rect 17359 8548 17371 8551
rect 18690 8548 18696 8560
rect 17359 8520 18696 8548
rect 17359 8517 17371 8520
rect 17313 8511 17371 8517
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6914 8480 6920 8492
rect 6512 8452 6920 8480
rect 6512 8440 6518 8452
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 8628 8452 9352 8480
rect 8628 8440 8634 8452
rect 2648 8384 3372 8412
rect 3605 8415 3663 8421
rect 2648 8372 2654 8384
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 3694 8412 3700 8424
rect 3651 8384 3700 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4304 8384 4353 8412
rect 4304 8372 4310 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 4608 8415 4666 8421
rect 4608 8381 4620 8415
rect 4654 8412 4666 8415
rect 5718 8412 5724 8424
rect 4654 8384 5724 8412
rect 4654 8381 4666 8384
rect 4608 8375 4666 8381
rect 2222 8353 2228 8356
rect 2216 8344 2228 8353
rect 2183 8316 2228 8344
rect 2216 8307 2228 8316
rect 2222 8304 2228 8307
rect 2280 8304 2286 8356
rect 4356 8344 4384 8375
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 6420 8384 7604 8412
rect 6420 8372 6426 8384
rect 5442 8344 5448 8356
rect 2746 8316 5448 8344
rect 2746 8276 2774 8316
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 5994 8344 6000 8356
rect 5955 8316 6000 8344
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 6144 8316 6469 8344
rect 6144 8304 6150 8316
rect 6457 8313 6469 8316
rect 6503 8313 6515 8347
rect 7374 8344 7380 8356
rect 6457 8307 6515 8313
rect 6932 8316 7380 8344
rect 6932 8288 6960 8316
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7576 8344 7604 8384
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8122 8415 8180 8421
rect 8122 8412 8134 8415
rect 7708 8384 8134 8412
rect 7708 8372 7714 8384
rect 8122 8381 8134 8384
rect 8168 8381 8180 8415
rect 8122 8375 8180 8381
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8527 8384 8861 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8849 8381 8861 8384
rect 8895 8412 8907 8415
rect 9214 8412 9220 8424
rect 8895 8384 9220 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 7576 8316 7696 8344
rect 1820 8248 2774 8276
rect 1820 8236 1826 8248
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 6914 8276 6920 8288
rect 5316 8248 6920 8276
rect 5316 8236 5322 8248
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 7009 8279 7067 8285
rect 7009 8245 7021 8279
rect 7055 8276 7067 8279
rect 7190 8276 7196 8288
rect 7055 8248 7196 8276
rect 7055 8245 7067 8248
rect 7009 8239 7067 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7668 8276 7696 8316
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 8202 8344 8208 8356
rect 7800 8316 8208 8344
rect 7800 8304 7806 8316
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 8404 8344 8432 8375
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 9324 8421 9352 8452
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 9456 8452 10241 8480
rect 9456 8440 9462 8452
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10468 8452 11069 8480
rect 10468 8440 10474 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11974 8480 11980 8492
rect 11935 8452 11980 8480
rect 11057 8443 11115 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 13449 8483 13507 8489
rect 13449 8480 13461 8483
rect 12406 8452 13461 8480
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 10870 8412 10876 8424
rect 9999 8384 10876 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 12406 8412 12434 8452
rect 13449 8449 13461 8452
rect 13495 8449 13507 8483
rect 15286 8480 15292 8492
rect 15247 8452 15292 8480
rect 13449 8443 13507 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 12894 8412 12900 8424
rect 10980 8384 12434 8412
rect 12855 8384 12900 8412
rect 8260 8316 9812 8344
rect 8260 8304 8266 8316
rect 9784 8285 9812 8316
rect 8481 8279 8539 8285
rect 8481 8276 8493 8279
rect 7668 8248 8493 8276
rect 8481 8245 8493 8248
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8276 9827 8279
rect 10502 8276 10508 8288
rect 9815 8248 10508 8276
rect 9815 8245 9827 8248
rect 9769 8239 9827 8245
rect 10502 8236 10508 8248
rect 10560 8276 10566 8288
rect 10980 8276 11008 8384
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 13596 8384 17141 8412
rect 13596 8372 13602 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 12434 8344 12440 8356
rect 12207 8316 12440 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 13716 8347 13774 8353
rect 13716 8313 13728 8347
rect 13762 8344 13774 8347
rect 14734 8344 14740 8356
rect 13762 8316 14740 8344
rect 13762 8313 13774 8316
rect 13716 8307 13774 8313
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 15473 8347 15531 8353
rect 15473 8313 15485 8347
rect 15519 8344 15531 8347
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15519 8316 16129 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 16117 8313 16129 8316
rect 16163 8313 16175 8347
rect 16117 8307 16175 8313
rect 10560 8248 11008 8276
rect 10560 8236 10566 8248
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 11756 8248 12265 8276
rect 11756 8236 11762 8248
rect 12253 8245 12265 8248
rect 12299 8245 12311 8279
rect 15378 8276 15384 8288
rect 15339 8248 15384 8276
rect 12253 8239 12311 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 15746 8236 15752 8288
rect 15804 8276 15810 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15804 8248 15853 8276
rect 15804 8236 15810 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1394 8072 1400 8084
rect 1355 8044 1400 8072
rect 1394 8032 1400 8044
rect 1452 8032 1458 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2866 8072 2872 8084
rect 2823 8044 2872 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4212 8044 4353 8072
rect 4212 8032 4218 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 4341 8035 4399 8041
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 4798 8072 4804 8084
rect 4755 8044 4804 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5626 8072 5632 8084
rect 4908 8044 5632 8072
rect 3145 8007 3203 8013
rect 2056 7976 3096 8004
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 2056 7945 2084 7976
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 1728 7908 2053 7936
rect 1728 7896 1734 7908
rect 2041 7905 2053 7908
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2590 7936 2596 7948
rect 2179 7908 2596 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 3068 7936 3096 7976
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 4908 8004 4936 8044
rect 5626 8032 5632 8044
rect 5684 8072 5690 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5684 8044 5733 8072
rect 5684 8032 5690 8044
rect 5721 8041 5733 8044
rect 5767 8041 5779 8075
rect 5721 8035 5779 8041
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 6595 8044 7665 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8067 8044 9597 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 11974 8072 11980 8084
rect 11931 8044 11980 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 11974 8032 11980 8044
rect 12032 8072 12038 8084
rect 13909 8075 13967 8081
rect 12032 8044 12434 8072
rect 12032 8032 12038 8044
rect 5810 8004 5816 8016
rect 3191 7976 4936 8004
rect 5000 7976 5816 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 4890 7936 4896 7948
rect 3068 7908 4896 7936
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 2774 7868 2780 7880
rect 1949 7831 2007 7837
rect 1964 7732 1992 7831
rect 2746 7828 2780 7868
rect 2832 7828 2838 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 2746 7800 2774 7828
rect 2547 7772 2774 7800
rect 3252 7800 3280 7831
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4798 7868 4804 7880
rect 3384 7840 3429 7868
rect 4759 7840 4804 7868
rect 3384 7828 3390 7840
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5000 7877 5028 7976
rect 5810 7964 5816 7976
rect 5868 7964 5874 8016
rect 7926 8004 7932 8016
rect 7576 7976 7932 8004
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 5307 7908 6377 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 6365 7905 6377 7908
rect 6411 7936 6423 7939
rect 6638 7936 6644 7948
rect 6411 7908 6644 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7098 7936 7104 7948
rect 7055 7908 7104 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7576 7936 7604 7976
rect 7926 7964 7932 7976
rect 7984 8004 7990 8016
rect 12406 8004 12434 8044
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 14090 8072 14096 8084
rect 13955 8044 14096 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 14090 8032 14096 8044
rect 14148 8072 14154 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14148 8044 14841 8072
rect 14148 8032 14154 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 15378 8072 15384 8084
rect 15335 8044 15384 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 13274 8007 13332 8013
rect 13274 8004 13286 8007
rect 7984 7976 12204 8004
rect 12406 7976 13286 8004
rect 7984 7964 7990 7976
rect 7484 7908 7604 7936
rect 8481 7939 8539 7945
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6178 7868 6184 7880
rect 6043 7840 6184 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 5534 7800 5540 7812
rect 3252 7772 5540 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 5828 7800 5856 7831
rect 6178 7828 6184 7840
rect 6236 7868 6242 7880
rect 7190 7868 7196 7880
rect 6236 7840 7196 7868
rect 6236 7828 6242 7840
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7484 7877 7512 7908
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8938 7936 8944 7948
rect 8527 7908 8944 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8938 7896 8944 7908
rect 8996 7936 9002 7948
rect 9490 7936 9496 7948
rect 8996 7908 9496 7936
rect 8996 7896 9002 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10502 7936 10508 7948
rect 10463 7908 10508 7936
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10772 7939 10830 7945
rect 10772 7905 10784 7939
rect 10818 7936 10830 7939
rect 11974 7936 11980 7948
rect 10818 7908 11980 7936
rect 10818 7905 10830 7908
rect 10772 7899 10830 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 9398 7868 9404 7880
rect 9359 7840 9404 7868
rect 7561 7831 7619 7837
rect 6638 7800 6644 7812
rect 5828 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 7374 7760 7380 7812
rect 7432 7800 7438 7812
rect 7576 7800 7604 7831
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 8294 7800 8300 7812
rect 7432 7772 7604 7800
rect 8255 7772 8300 7800
rect 7432 7760 7438 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 12176 7809 12204 7976
rect 13274 7973 13286 7976
rect 13320 7973 13332 8007
rect 14918 8004 14924 8016
rect 14879 7976 14924 8004
rect 13274 7967 13332 7973
rect 14918 7964 14924 7976
rect 14976 7964 14982 8016
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 15562 7936 15568 7948
rect 13587 7908 15568 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7769 12219 7803
rect 12161 7763 12219 7769
rect 2222 7732 2228 7744
rect 1964 7704 2228 7732
rect 2222 7692 2228 7704
rect 2280 7732 2286 7744
rect 3326 7732 3332 7744
rect 2280 7704 3332 7732
rect 2280 7692 2286 7704
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3844 7704 3985 7732
rect 3844 7692 3850 7704
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 4120 7704 5273 7732
rect 4120 7692 4126 7704
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7732 5411 7735
rect 5626 7732 5632 7744
rect 5399 7704 5632 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 6604 7704 6837 7732
rect 6604 7692 6610 7704
rect 6825 7701 6837 7704
rect 6871 7701 6883 7735
rect 6825 7695 6883 7701
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7732 10103 7735
rect 11238 7732 11244 7744
rect 10091 7704 11244 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13556 7732 13584 7899
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15746 7936 15752 7948
rect 15707 7908 15752 7936
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17322 7939 17380 7945
rect 17322 7936 17334 7939
rect 16632 7908 17334 7936
rect 16632 7896 16638 7908
rect 17322 7905 17334 7908
rect 17368 7905 17380 7939
rect 17322 7899 17380 7905
rect 14734 7868 14740 7880
rect 14647 7840 14740 7868
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17678 7868 17684 7880
rect 17635 7840 17684 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 14752 7800 14780 7828
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 14752 7772 16221 7800
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16209 7763 16267 7769
rect 13320 7704 13584 7732
rect 15933 7735 15991 7741
rect 13320 7692 13326 7704
rect 15933 7701 15945 7735
rect 15979 7732 15991 7735
rect 17862 7732 17868 7744
rect 15979 7704 17868 7732
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3326 7528 3332 7540
rect 3191 7500 3332 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5169 7531 5227 7537
rect 5169 7528 5181 7531
rect 4856 7500 5181 7528
rect 4856 7488 4862 7500
rect 5169 7497 5181 7500
rect 5215 7497 5227 7531
rect 5169 7491 5227 7497
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6503 7500 6653 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12032 7500 12388 7528
rect 12032 7488 12038 7500
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 6822 7460 6828 7472
rect 3651 7432 6828 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 9033 7463 9091 7469
rect 9033 7429 9045 7463
rect 9079 7429 9091 7463
rect 9033 7423 9091 7429
rect 5626 7392 5632 7404
rect 5587 7364 5632 7392
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 7190 7392 7196 7404
rect 5776 7364 5821 7392
rect 7151 7364 7196 7392
rect 5776 7352 5782 7364
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 9048 7392 9076 7423
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12360 7460 12388 7500
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12621 7531 12679 7537
rect 12621 7528 12633 7531
rect 12492 7500 12633 7528
rect 12492 7488 12498 7500
rect 12621 7497 12633 7500
rect 12667 7497 12679 7531
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 12621 7491 12679 7497
rect 13372 7500 15025 7528
rect 13372 7460 13400 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 11940 7432 12296 7460
rect 12360 7432 13400 7460
rect 11940 7420 11946 7432
rect 11333 7395 11391 7401
rect 9048 7364 9444 7392
rect 9416 7336 9444 7364
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 11698 7392 11704 7404
rect 11379 7364 11704 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 11974 7392 11980 7404
rect 11935 7364 11980 7392
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 2746 7296 3433 7324
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 2010 7259 2068 7265
rect 2010 7256 2022 7259
rect 1544 7228 2022 7256
rect 1544 7216 1550 7228
rect 2010 7225 2022 7228
rect 2056 7225 2068 7259
rect 2010 7219 2068 7225
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7188 1458 7200
rect 2746 7188 2774 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 3970 7324 3976 7336
rect 3927 7296 3976 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4338 7324 4344 7336
rect 4299 7296 4344 7324
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 4430 7284 4436 7336
rect 4488 7324 4494 7336
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4488 7296 4813 7324
rect 4488 7284 4494 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 7653 7327 7711 7333
rect 4801 7287 4859 7293
rect 5460 7296 7604 7324
rect 5460 7256 5488 7296
rect 4080 7228 5488 7256
rect 5537 7259 5595 7265
rect 4080 7197 4108 7228
rect 5537 7225 5549 7259
rect 5583 7256 5595 7259
rect 6457 7259 6515 7265
rect 6457 7256 6469 7259
rect 5583 7228 6469 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 6457 7225 6469 7228
rect 6503 7225 6515 7259
rect 6457 7219 6515 7225
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 6972 7228 7021 7256
rect 6972 7216 6978 7228
rect 7009 7225 7021 7228
rect 7055 7225 7067 7259
rect 7576 7256 7604 7296
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7742 7324 7748 7336
rect 7699 7296 7748 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7926 7333 7932 7336
rect 7920 7324 7932 7333
rect 7887 7296 7932 7324
rect 7920 7287 7932 7296
rect 7926 7284 7932 7287
rect 7984 7284 7990 7336
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9214 7256 9220 7268
rect 7576 7228 9220 7256
rect 7009 7219 7067 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 9324 7256 9352 7287
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9565 7327 9623 7333
rect 9565 7324 9577 7327
rect 9456 7296 9577 7324
rect 9456 7284 9462 7296
rect 9565 7293 9577 7296
rect 9611 7293 9623 7327
rect 9565 7287 9623 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12268 7333 12296 7432
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13320 7364 13369 7392
rect 13320 7352 13326 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 12124 7296 12173 7324
rect 12124 7284 12130 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7293 12311 7327
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12253 7287 12311 7293
rect 12406 7296 12909 7324
rect 10502 7256 10508 7268
rect 9324 7228 10508 7256
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 12406 7256 12434 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 16393 7327 16451 7333
rect 12897 7287 12955 7293
rect 14568 7296 16252 7324
rect 11940 7228 12434 7256
rect 11940 7216 11946 7228
rect 13538 7216 13544 7268
rect 13596 7265 13602 7268
rect 13596 7259 13660 7265
rect 13596 7225 13614 7259
rect 13648 7225 13660 7259
rect 13596 7219 13660 7225
rect 13596 7216 13602 7219
rect 1452 7160 2774 7188
rect 4065 7191 4123 7197
rect 1452 7148 1458 7160
rect 4065 7157 4077 7191
rect 4111 7157 4123 7191
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4065 7151 4123 7157
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 4948 7160 7113 7188
rect 4948 7148 4954 7160
rect 7101 7157 7113 7160
rect 7147 7188 7159 7191
rect 9582 7188 9588 7200
rect 7147 7160 9588 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 14568 7188 14596 7296
rect 16126 7259 16184 7265
rect 16126 7256 16138 7259
rect 14752 7228 16138 7256
rect 14752 7200 14780 7228
rect 16126 7225 16138 7228
rect 16172 7225 16184 7259
rect 16224 7256 16252 7296
rect 16393 7293 16405 7327
rect 16439 7324 16451 7327
rect 17678 7324 17684 7336
rect 16439 7296 17684 7324
rect 16439 7293 16451 7296
rect 16393 7287 16451 7293
rect 17678 7284 17684 7296
rect 17736 7284 17742 7336
rect 16945 7259 17003 7265
rect 16945 7256 16957 7259
rect 16224 7228 16957 7256
rect 16126 7219 16184 7225
rect 16945 7225 16957 7228
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 14734 7188 14740 7200
rect 10836 7160 14596 7188
rect 14647 7160 14740 7188
rect 10836 7148 10842 7160
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 2372 6956 3157 6984
rect 2372 6944 2378 6956
rect 3145 6953 3157 6956
rect 3191 6953 3203 6987
rect 3145 6947 3203 6953
rect 4522 6944 4528 6996
rect 4580 6984 4586 6996
rect 14182 6984 14188 6996
rect 4580 6956 14188 6984
rect 4580 6944 4586 6956
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 2133 6919 2191 6925
rect 2133 6885 2145 6919
rect 2179 6916 2191 6919
rect 3050 6916 3056 6928
rect 2179 6888 3056 6916
rect 2179 6885 2191 6888
rect 2133 6879 2191 6885
rect 3050 6876 3056 6888
rect 3108 6876 3114 6928
rect 4080 6888 5304 6916
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6848 1547 6851
rect 2774 6848 2780 6860
rect 1535 6820 2780 6848
rect 1535 6817 1547 6820
rect 1489 6811 1547 6817
rect 2774 6808 2780 6820
rect 2832 6848 2838 6860
rect 4080 6848 4108 6888
rect 5178 6851 5236 6857
rect 5178 6848 5190 6851
rect 2832 6820 4108 6848
rect 4172 6820 5190 6848
rect 2832 6808 2838 6820
rect 4172 6792 4200 6820
rect 5178 6817 5190 6820
rect 5224 6817 5236 6851
rect 5276 6848 5304 6888
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 5408 6888 6040 6916
rect 5408 6876 5414 6888
rect 5905 6851 5963 6857
rect 5905 6848 5917 6851
rect 5276 6820 5917 6848
rect 5178 6811 5236 6817
rect 5905 6817 5917 6820
rect 5951 6817 5963 6851
rect 6012 6848 6040 6888
rect 9416 6888 11008 6916
rect 6178 6848 6184 6860
rect 6012 6820 6184 6848
rect 5905 6811 5963 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 6328 6820 6377 6848
rect 6328 6808 6334 6820
rect 6365 6817 6377 6820
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6880 6820 7021 6848
rect 6880 6808 6886 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6848 7159 6851
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7147 6820 7757 6848
rect 7147 6817 7159 6820
rect 7101 6811 7159 6817
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8260 6820 8401 6848
rect 8260 6808 8266 6820
rect 8389 6817 8401 6820
rect 8435 6848 8447 6851
rect 9416 6848 9444 6888
rect 8435 6820 9444 6848
rect 9493 6851 9551 6857
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9674 6848 9680 6860
rect 9539 6820 9680 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2958 6780 2964 6792
rect 2455 6752 2964 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2240 6712 2268 6743
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3421 6783 3479 6789
rect 3283 6752 3372 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2240 6684 2789 6712
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 2130 6644 2136 6656
rect 1811 6616 2136 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 3344 6644 3372 6752
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 4154 6780 4160 6792
rect 3467 6752 4160 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6914 6780 6920 6792
rect 5552 6752 6316 6780
rect 6875 6752 6920 6780
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3752 6684 4077 6712
rect 3752 6672 3758 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 5166 6644 5172 6656
rect 3344 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5552 6644 5580 6752
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5684 6684 6193 6712
rect 5684 6672 5690 6684
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 6288 6712 6316 6752
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 8665 6783 8723 6789
rect 8665 6780 8677 6783
rect 7024 6752 8677 6780
rect 7024 6712 7052 6752
rect 8665 6749 8677 6752
rect 8711 6749 8723 6783
rect 9968 6780 9996 6811
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10853 6851 10911 6857
rect 10853 6848 10865 6851
rect 10376 6820 10865 6848
rect 10376 6808 10382 6820
rect 10853 6817 10865 6820
rect 10899 6817 10911 6851
rect 10980 6848 11008 6888
rect 11238 6876 11244 6928
rect 11296 6916 11302 6928
rect 11296 6888 13216 6916
rect 11296 6876 11302 6888
rect 12437 6851 12495 6857
rect 10980 6820 12388 6848
rect 10853 6811 10911 6817
rect 10410 6780 10416 6792
rect 8665 6743 8723 6749
rect 9692 6752 10416 6780
rect 9692 6724 9720 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10560 6752 10609 6780
rect 10560 6740 10566 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 6288 6684 7052 6712
rect 7469 6715 7527 6721
rect 6181 6675 6239 6681
rect 7469 6681 7481 6715
rect 7515 6712 7527 6715
rect 8478 6712 8484 6724
rect 7515 6684 8484 6712
rect 7515 6681 7527 6684
rect 7469 6675 7527 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 9674 6672 9680 6724
rect 9732 6672 9738 6724
rect 9769 6715 9827 6721
rect 9769 6681 9781 6715
rect 9815 6712 9827 6715
rect 10042 6712 10048 6724
rect 9815 6684 10048 6712
rect 9815 6681 9827 6684
rect 9769 6675 9827 6681
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 5718 6644 5724 6656
rect 5316 6616 5580 6644
rect 5679 6616 5724 6644
rect 5316 6604 5322 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 6788 6616 8217 6644
rect 6788 6604 6794 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 8812 6616 10241 6644
rect 8812 6604 8818 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 11974 6644 11980 6656
rect 11935 6616 11980 6644
rect 10229 6607 10287 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12250 6644 12256 6656
rect 12211 6616 12256 6644
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12360 6644 12388 6820
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12483 6820 12909 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 13078 6848 13084 6860
rect 13039 6820 13084 6848
rect 12897 6811 12955 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13188 6712 13216 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14792 6888 15148 6916
rect 14792 6876 14798 6888
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13412 6820 13553 6848
rect 13412 6808 13418 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 14918 6848 14924 6860
rect 14879 6820 14924 6848
rect 13541 6811 13599 6817
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15120 6789 15148 6888
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 16942 6848 16948 6860
rect 15565 6811 15623 6817
rect 15764 6820 16948 6848
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 15580 6712 15608 6811
rect 15764 6721 15792 6820
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17218 6808 17224 6860
rect 17276 6857 17282 6860
rect 17276 6848 17288 6857
rect 17276 6820 17321 6848
rect 17276 6811 17288 6820
rect 17276 6808 17282 6811
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17678 6780 17684 6792
rect 17543 6752 17684 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 13188 6684 15608 6712
rect 15749 6715 15807 6721
rect 15749 6681 15761 6715
rect 15795 6681 15807 6715
rect 15749 6675 15807 6681
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12360 6616 12725 6644
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13262 6644 13268 6656
rect 12943 6616 13268 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 14366 6644 14372 6656
rect 13771 6616 14372 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 16117 6647 16175 6653
rect 16117 6613 16129 6647
rect 16163 6644 16175 6647
rect 16574 6644 16580 6656
rect 16163 6616 16580 6644
rect 16163 6613 16175 6616
rect 16117 6607 16175 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 1486 6440 1492 6452
rect 1443 6412 1492 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 1486 6400 1492 6412
rect 1544 6400 1550 6452
rect 8386 6440 8392 6452
rect 6840 6412 8392 6440
rect 2958 6372 2964 6384
rect 2871 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6372 3022 6384
rect 3694 6372 3700 6384
rect 3016 6344 3700 6372
rect 3016 6332 3022 6344
rect 3694 6332 3700 6344
rect 3752 6332 3758 6384
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6341 4675 6375
rect 4617 6335 4675 6341
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 4154 6304 4160 6316
rect 4115 6276 4160 6304
rect 4154 6264 4160 6276
rect 4212 6304 4218 6316
rect 4632 6304 4660 6335
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 6840 6372 6868 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 13354 6440 13360 6452
rect 8720 6412 13360 6440
rect 8720 6400 8726 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13538 6440 13544 6452
rect 13499 6412 13544 6440
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 15010 6440 15016 6452
rect 14599 6412 15016 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6440 16635 6443
rect 18598 6440 18604 6452
rect 16623 6412 18604 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 6236 6344 6868 6372
rect 9861 6375 9919 6381
rect 6236 6332 6242 6344
rect 9861 6341 9873 6375
rect 9907 6372 9919 6375
rect 9907 6344 10364 6372
rect 9907 6341 9919 6344
rect 9861 6335 9919 6341
rect 10336 6316 10364 6344
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 10560 6344 10916 6372
rect 10560 6332 10566 6344
rect 4212 6276 4660 6304
rect 5997 6307 6055 6313
rect 4212 6264 4218 6276
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6454 6304 6460 6316
rect 6043 6276 6460 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6454 6264 6460 6276
rect 6512 6304 6518 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6512 6276 6837 6304
rect 6512 6264 6518 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 6825 6267 6883 6273
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10778 6304 10784 6316
rect 10459 6276 10784 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10888 6304 10916 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11238 6372 11244 6384
rect 11112 6344 11244 6372
rect 11112 6332 11118 6344
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 10888 6276 11928 6304
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2866 6236 2872 6248
rect 2823 6208 2872 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3660 6208 3985 6236
rect 3660 6196 3666 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 4856 6208 6561 6236
rect 4856 6196 4862 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7081 6239 7139 6245
rect 7081 6236 7093 6239
rect 6972 6208 7093 6236
rect 6972 6196 6978 6208
rect 7081 6205 7093 6208
rect 7127 6205 7139 6239
rect 7081 6199 7139 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 9122 6236 9128 6248
rect 8527 6208 9128 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9272 6208 10517 6236
rect 9272 6196 9278 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 11333 6239 11391 6245
rect 11333 6236 11345 6239
rect 10505 6199 10563 6205
rect 10704 6208 11345 6236
rect 2532 6171 2590 6177
rect 2532 6137 2544 6171
rect 2578 6168 2590 6171
rect 2961 6171 3019 6177
rect 2961 6168 2973 6171
rect 2578 6140 2973 6168
rect 2578 6137 2590 6140
rect 2532 6131 2590 6137
rect 2961 6137 2973 6140
rect 3007 6137 3019 6171
rect 2961 6131 3019 6137
rect 5718 6128 5724 6180
rect 5776 6177 5782 6180
rect 5776 6168 5788 6177
rect 8726 6171 8784 6177
rect 8726 6168 8738 6171
rect 5776 6140 5821 6168
rect 8312 6140 8738 6168
rect 5776 6131 5788 6140
rect 5776 6128 5782 6131
rect 8312 6112 8340 6140
rect 8726 6137 8738 6140
rect 8772 6137 8784 6171
rect 8726 6131 8784 6137
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 10410 6168 10416 6180
rect 9456 6140 10416 6168
rect 9456 6128 9462 6140
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3292 6072 3617 6100
rect 3292 6060 3298 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 6270 6100 6276 6112
rect 4111 6072 6276 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 7098 6100 7104 6112
rect 6604 6072 7104 6100
rect 6604 6060 6610 6072
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8294 6100 8300 6112
rect 8251 6072 8300 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9030 6060 9036 6112
rect 9088 6100 9094 6112
rect 10704 6100 10732 6208
rect 11333 6205 11345 6208
rect 11379 6236 11391 6239
rect 11900 6236 11928 6276
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 13556 6304 13584 6400
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 12032 6276 12296 6304
rect 13556 6276 13921 6304
rect 12032 6264 12038 6276
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11379 6208 11836 6236
rect 11900 6208 12173 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 10870 6100 10876 6112
rect 9088 6072 10732 6100
rect 10831 6072 10876 6100
rect 9088 6060 9094 6072
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11112 6072 11161 6100
rect 11112 6060 11118 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11149 6063 11207 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11808 6100 11836 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12268 6236 12296 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14976 6276 15025 6304
rect 14976 6264 14982 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 16574 6304 16580 6316
rect 16071 6276 16580 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16574 6264 16580 6276
rect 16632 6264 16638 6316
rect 17126 6264 17132 6316
rect 17184 6304 17190 6316
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 17184 6276 17693 6304
rect 17184 6264 17190 6276
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 12417 6239 12475 6245
rect 12417 6236 12429 6239
rect 12268 6208 12429 6236
rect 12161 6199 12219 6205
rect 12417 6205 12429 6208
rect 12463 6205 12475 6239
rect 12417 6199 12475 6205
rect 12176 6168 12204 6199
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 13320 6208 15393 6236
rect 13320 6196 13326 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 17586 6236 17592 6248
rect 17547 6208 17592 6236
rect 15381 6199 15439 6205
rect 17586 6196 17592 6208
rect 17644 6236 17650 6248
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 17644 6208 18153 6236
rect 17644 6196 17650 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 12250 6168 12256 6180
rect 12176 6140 12256 6168
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 14182 6168 14188 6180
rect 14143 6140 14188 6168
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 16209 6171 16267 6177
rect 16209 6137 16221 6171
rect 16255 6168 16267 6171
rect 16255 6140 17172 6168
rect 16255 6137 16267 6140
rect 16209 6131 16267 6137
rect 13906 6100 13912 6112
rect 11808 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 16117 6103 16175 6109
rect 16117 6069 16129 6103
rect 16163 6100 16175 6103
rect 16390 6100 16396 6112
rect 16163 6072 16396 6100
rect 16163 6069 16175 6072
rect 16117 6063 16175 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17144 6109 17172 6140
rect 17129 6103 17187 6109
rect 17129 6069 17141 6103
rect 17175 6069 17187 6103
rect 17494 6100 17500 6112
rect 17455 6072 17500 6100
rect 17129 6063 17187 6069
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2130 5896 2136 5908
rect 2091 5868 2136 5896
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 2464 5868 2513 5896
rect 2464 5856 2470 5868
rect 2501 5865 2513 5868
rect 2547 5865 2559 5899
rect 3234 5896 3240 5908
rect 3195 5868 3240 5896
rect 2501 5859 2559 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 4065 5899 4123 5905
rect 4065 5865 4077 5899
rect 4111 5865 4123 5899
rect 4430 5896 4436 5908
rect 4391 5868 4436 5896
rect 4065 5859 4123 5865
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 4080 5828 4108 5859
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4982 5856 4988 5908
rect 5040 5896 5046 5908
rect 6178 5896 6184 5908
rect 5040 5868 6184 5896
rect 5040 5856 5046 5868
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 6822 5896 6828 5908
rect 6420 5868 6828 5896
rect 6420 5856 6426 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6972 5868 7389 5896
rect 6972 5856 6978 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 7377 5859 7435 5865
rect 3191 5800 4108 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4212 5800 4660 5828
rect 4212 5788 4218 5800
rect 3694 5760 3700 5772
rect 3436 5732 3700 5760
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 3436 5701 3464 5732
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1544 5664 1869 5692
rect 1544 5652 1550 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 3421 5695 3479 5701
rect 2087 5664 2820 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2792 5633 2820 5664
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3878 5692 3884 5704
rect 3568 5664 3884 5692
rect 3568 5652 3574 5664
rect 3878 5652 3884 5664
rect 3936 5692 3942 5704
rect 4632 5701 4660 5800
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 4948 5800 7236 5828
rect 4948 5788 4954 5800
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 4724 5732 5089 5760
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3936 5664 4537 5692
rect 3936 5652 3942 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5593 2835 5627
rect 2777 5587 2835 5593
rect 3786 5584 3792 5636
rect 3844 5624 3850 5636
rect 4724 5624 4752 5732
rect 5077 5729 5089 5732
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 5684 5732 5733 5760
rect 5684 5720 5690 5732
rect 5721 5729 5733 5732
rect 5767 5760 5779 5763
rect 6086 5760 6092 5772
rect 5767 5732 6092 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6264 5763 6322 5769
rect 6264 5729 6276 5763
rect 6310 5760 6322 5763
rect 7098 5760 7104 5772
rect 6310 5732 7104 5760
rect 6310 5729 6322 5732
rect 6264 5723 6322 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5500 5664 6009 5692
rect 5500 5652 5506 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 3844 5596 4752 5624
rect 5261 5627 5319 5633
rect 3844 5584 3850 5596
rect 5261 5593 5273 5627
rect 5307 5624 5319 5627
rect 7208 5624 7236 5800
rect 7392 5692 7420 5859
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7524 5868 10824 5896
rect 7524 5856 7530 5868
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 9674 5837 9680 5840
rect 8021 5831 8079 5837
rect 8021 5828 8033 5831
rect 7800 5800 8033 5828
rect 7800 5788 7806 5800
rect 8021 5797 8033 5800
rect 8067 5797 8079 5831
rect 9668 5828 9680 5837
rect 9587 5800 9680 5828
rect 8021 5791 8079 5797
rect 9668 5791 9680 5800
rect 9732 5828 9738 5840
rect 10686 5828 10692 5840
rect 9732 5800 10692 5828
rect 9674 5788 9680 5791
rect 9732 5788 9738 5800
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 10796 5828 10824 5868
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 10928 5868 12357 5896
rect 10928 5856 10934 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13412 5868 13860 5896
rect 13412 5856 13418 5868
rect 11054 5828 11060 5840
rect 10796 5800 11060 5828
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 12308 5800 13553 5828
rect 12308 5788 12314 5800
rect 13541 5797 13553 5800
rect 13587 5797 13599 5831
rect 13832 5828 13860 5868
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 15381 5899 15439 5905
rect 15381 5896 15393 5899
rect 13964 5868 15393 5896
rect 13964 5856 13970 5868
rect 15381 5865 15393 5868
rect 15427 5865 15439 5899
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 15381 5859 15439 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 17494 5856 17500 5908
rect 17552 5896 17558 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 17552 5868 17601 5896
rect 17552 5856 17558 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 16761 5831 16819 5837
rect 16761 5828 16773 5831
rect 13832 5800 16773 5828
rect 13541 5791 13599 5797
rect 16761 5797 16773 5800
rect 16807 5797 16819 5831
rect 16761 5791 16819 5797
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 8202 5760 8208 5772
rect 7524 5732 8208 5760
rect 7524 5720 7530 5732
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 9180 5732 9413 5760
rect 9180 5720 9186 5732
rect 9401 5729 9413 5732
rect 9447 5760 9459 5763
rect 9950 5760 9956 5772
rect 9447 5732 9956 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 11238 5760 11244 5772
rect 10468 5732 11244 5760
rect 10468 5720 10474 5732
rect 11238 5720 11244 5732
rect 11296 5760 11302 5772
rect 11701 5763 11759 5769
rect 11296 5732 11652 5760
rect 11296 5720 11302 5732
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7392 5664 7757 5692
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7745 5655 7803 5661
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 11054 5692 11060 5704
rect 8444 5664 8800 5692
rect 11015 5664 11060 5692
rect 8444 5652 8450 5664
rect 8665 5627 8723 5633
rect 8665 5624 8677 5627
rect 5307 5596 6040 5624
rect 7208 5596 8677 5624
rect 5307 5593 5319 5596
rect 5261 5587 5319 5593
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 1578 5556 1584 5568
rect 1535 5528 1584 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6012 5556 6040 5596
rect 8665 5593 8677 5596
rect 8711 5593 8723 5627
rect 8665 5587 8723 5593
rect 8202 5556 8208 5568
rect 6012 5528 8208 5556
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8386 5556 8392 5568
rect 8347 5528 8392 5556
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8772 5556 8800 5664
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 10336 5596 11529 5624
rect 10336 5556 10364 5596
rect 11517 5593 11529 5596
rect 11563 5593 11575 5627
rect 11624 5624 11652 5732
rect 11701 5729 11713 5763
rect 11747 5760 11759 5763
rect 11882 5760 11888 5772
rect 11747 5732 11888 5760
rect 11747 5729 11759 5732
rect 11701 5723 11759 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12483 5732 13093 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 14550 5760 14556 5772
rect 13320 5732 14044 5760
rect 14511 5732 14556 5760
rect 13320 5720 13326 5732
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 12032 5664 12173 5692
rect 12032 5652 12038 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 12676 5664 13921 5692
rect 12676 5652 12682 5664
rect 13909 5661 13921 5664
rect 13955 5661 13967 5695
rect 14016 5692 14044 5732
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 17957 5763 18015 5769
rect 17957 5760 17969 5763
rect 15896 5732 17969 5760
rect 15896 5720 15902 5732
rect 17957 5729 17969 5732
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5760 20959 5763
rect 21358 5760 21364 5772
rect 20947 5732 21364 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14016 5664 15025 5692
rect 13909 5655 13967 5661
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16724 5664 16865 5692
rect 16724 5652 16730 5664
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17126 5692 17132 5704
rect 17083 5664 17132 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 18233 5627 18291 5633
rect 18233 5624 18245 5627
rect 11624 5596 18245 5624
rect 11517 5587 11575 5593
rect 18233 5593 18245 5596
rect 18279 5593 18291 5627
rect 18233 5587 18291 5593
rect 10778 5556 10784 5568
rect 8772 5528 10364 5556
rect 10739 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 12805 5559 12863 5565
rect 12805 5525 12817 5559
rect 12851 5556 12863 5559
rect 12894 5556 12900 5568
rect 12851 5528 12900 5556
rect 12851 5525 12863 5528
rect 12805 5519 12863 5525
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14608 5528 14749 5556
rect 14608 5516 14614 5528
rect 14737 5525 14749 5528
rect 14783 5525 14795 5559
rect 15746 5556 15752 5568
rect 15707 5528 15752 5556
rect 14737 5519 14795 5525
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 21174 5556 21180 5568
rect 21135 5528 21180 5556
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 5626 5352 5632 5364
rect 4028 5324 5632 5352
rect 4028 5312 4034 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 5902 5352 5908 5364
rect 5863 5324 5908 5352
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 7926 5352 7932 5364
rect 7791 5324 7932 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8294 5312 8300 5364
rect 8352 5312 8358 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 11238 5352 11244 5364
rect 8803 5324 11244 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11848 5324 11897 5352
rect 11848 5312 11854 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 12342 5352 12348 5364
rect 12303 5324 12348 5352
rect 11885 5315 11943 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 17126 5352 17132 5364
rect 17087 5324 17132 5352
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5284 1915 5287
rect 2314 5284 2320 5296
rect 1903 5256 2320 5284
rect 1903 5253 1915 5256
rect 1857 5247 1915 5253
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 4525 5287 4583 5293
rect 2424 5256 3464 5284
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2424 5216 2452 5256
rect 2004 5188 2452 5216
rect 2593 5219 2651 5225
rect 2004 5176 2010 5188
rect 2593 5185 2605 5219
rect 2639 5216 2651 5219
rect 3326 5216 3332 5228
rect 2639 5188 3332 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3436 5225 3464 5256
rect 4525 5253 4537 5287
rect 4571 5284 4583 5287
rect 7190 5284 7196 5296
rect 4571 5256 7196 5284
rect 4571 5253 4583 5256
rect 4525 5247 4583 5253
rect 7190 5244 7196 5256
rect 7248 5284 7254 5296
rect 8312 5284 8340 5312
rect 7248 5256 7880 5284
rect 7248 5244 7254 5256
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 4120 5188 6469 5216
rect 4120 5176 4126 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 7098 5216 7104 5228
rect 7059 5188 7104 5216
rect 6457 5179 6515 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 3694 5148 3700 5160
rect 1719 5120 3700 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 3878 5148 3884 5160
rect 3839 5120 3884 5148
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4338 5148 4344 5160
rect 4299 5120 4344 5148
rect 4338 5108 4344 5120
rect 4396 5108 4402 5160
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 4890 5148 4896 5160
rect 4847 5120 4896 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5258 5148 5264 5160
rect 5219 5120 5264 5148
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5500 5120 5733 5148
rect 5500 5108 5506 5120
rect 5721 5117 5733 5120
rect 5767 5148 5779 5151
rect 5994 5148 6000 5160
rect 5767 5120 6000 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 7374 5148 7380 5160
rect 7335 5120 7380 5148
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7852 5148 7880 5256
rect 8220 5256 8340 5284
rect 11057 5287 11115 5293
rect 8220 5225 8248 5256
rect 11057 5253 11069 5287
rect 11103 5253 11115 5287
rect 11057 5247 11115 5253
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9674 5216 9680 5228
rect 9539 5188 9680 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10778 5216 10784 5228
rect 10551 5188 10784 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 11072 5216 11100 5247
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 14093 5287 14151 5293
rect 14093 5284 14105 5287
rect 12124 5256 14105 5284
rect 12124 5244 12130 5256
rect 14093 5253 14105 5256
rect 14139 5253 14151 5287
rect 14093 5247 14151 5253
rect 16209 5287 16267 5293
rect 16209 5253 16221 5287
rect 16255 5284 16267 5287
rect 17402 5284 17408 5296
rect 16255 5256 17408 5284
rect 16255 5253 16267 5256
rect 16209 5247 16267 5253
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 15654 5216 15660 5228
rect 11072 5188 14504 5216
rect 15615 5188 15660 5216
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 7852 5120 9597 5148
rect 9585 5117 9597 5120
rect 9631 5148 9643 5151
rect 10042 5148 10048 5160
rect 9631 5120 10048 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11054 5148 11060 5160
rect 10735 5120 11060 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 12066 5148 12072 5160
rect 12027 5120 12072 5148
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12529 5151 12587 5157
rect 12529 5117 12541 5151
rect 12575 5148 12587 5151
rect 12618 5148 12624 5160
rect 12575 5120 12624 5148
rect 12575 5117 12587 5120
rect 12529 5111 12587 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12894 5148 12900 5160
rect 12855 5120 12900 5148
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 14476 5157 14504 5188
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 14700 5120 14933 5148
rect 14700 5108 14706 5120
rect 14921 5117 14933 5120
rect 14967 5117 14979 5151
rect 15838 5148 15844 5160
rect 15799 5120 15844 5148
rect 14921 5111 14979 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 18506 5148 18512 5160
rect 17736 5120 18512 5148
rect 17736 5108 17742 5120
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 2130 5040 2136 5092
rect 2188 5080 2194 5092
rect 2777 5083 2835 5089
rect 2777 5080 2789 5083
rect 2188 5052 2789 5080
rect 2188 5040 2194 5052
rect 2777 5049 2789 5052
rect 2823 5049 2835 5083
rect 2777 5043 2835 5049
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 7392 5080 7420 5108
rect 4304 5052 7420 5080
rect 8389 5083 8447 5089
rect 4304 5040 4310 5052
rect 8389 5049 8401 5083
rect 8435 5080 8447 5083
rect 8478 5080 8484 5092
rect 8435 5052 8484 5080
rect 8435 5049 8447 5052
rect 8389 5043 8447 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 9677 5083 9735 5089
rect 9677 5049 9689 5083
rect 9723 5080 9735 5083
rect 9858 5080 9864 5092
rect 9723 5052 9864 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 10318 5040 10324 5092
rect 10376 5080 10382 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 10376 5052 15761 5080
rect 10376 5040 10382 5052
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15749 5043 15807 5049
rect 17218 5040 17224 5092
rect 17276 5080 17282 5092
rect 18242 5083 18300 5089
rect 18242 5080 18254 5083
rect 17276 5052 18254 5080
rect 17276 5040 17282 5052
rect 18242 5049 18254 5052
rect 18288 5049 18300 5083
rect 18242 5043 18300 5049
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 2464 4984 2697 5012
rect 2464 4972 2470 4984
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 3142 5012 3148 5024
rect 3103 4984 3148 5012
rect 2685 4975 2743 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4706 5012 4712 5024
rect 4111 4984 4712 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4985 5015 5043 5021
rect 4985 4981 4997 5015
rect 5031 5012 5043 5015
rect 5350 5012 5356 5024
rect 5031 4984 5356 5012
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5626 5012 5632 5024
rect 5491 4984 5632 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7650 5012 7656 5024
rect 7331 4984 7656 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7650 4972 7656 4984
rect 7708 5012 7714 5024
rect 9306 5012 9312 5024
rect 7708 4984 9312 5012
rect 7708 4972 7714 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 10045 5015 10103 5021
rect 10045 4981 10057 5015
rect 10091 5012 10103 5015
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 10091 4984 10609 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 10597 4975 10655 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13722 5012 13728 5024
rect 13683 4984 13728 5012
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 14645 5015 14703 5021
rect 14645 4981 14657 5015
rect 14691 5012 14703 5015
rect 14734 5012 14740 5024
rect 14691 4984 14740 5012
rect 14691 4981 14703 4984
rect 14645 4975 14703 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 15105 5015 15163 5021
rect 15105 4981 15117 5015
rect 15151 5012 15163 5015
rect 15378 5012 15384 5024
rect 15151 4984 15384 5012
rect 15151 4981 15163 4984
rect 15105 4975 15163 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16574 5012 16580 5024
rect 16535 4984 16580 5012
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1946 4808 1952 4820
rect 1811 4780 1952 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2130 4808 2136 4820
rect 2091 4780 2136 4808
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 5534 4808 5540 4820
rect 2516 4780 5540 4808
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 2516 4672 2544 4780
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 5684 4780 7512 4808
rect 5684 4768 5690 4780
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 2869 4743 2927 4749
rect 2869 4740 2881 4743
rect 2740 4712 2881 4740
rect 2740 4700 2746 4712
rect 2869 4709 2881 4712
rect 2915 4709 2927 4743
rect 5902 4740 5908 4752
rect 2869 4703 2927 4709
rect 5368 4712 5908 4740
rect 1719 4644 2544 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 4062 4672 4068 4684
rect 2832 4644 2877 4672
rect 4023 4644 4068 4672
rect 2832 4632 2838 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4706 4672 4712 4684
rect 4667 4644 4712 4672
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 5368 4613 5396 4712
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 6086 4700 6092 4752
rect 6144 4740 6150 4752
rect 7484 4749 7512 4780
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7800 4780 7849 4808
rect 7800 4768 7806 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8846 4808 8852 4820
rect 8619 4780 8852 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 9766 4808 9772 4820
rect 9631 4780 9772 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10134 4808 10140 4820
rect 10091 4780 10140 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 12161 4811 12219 4817
rect 12161 4808 12173 4811
rect 11204 4780 12173 4808
rect 11204 4768 11210 4780
rect 12161 4777 12173 4780
rect 12207 4777 12219 4811
rect 13722 4808 13728 4820
rect 12161 4771 12219 4777
rect 12268 4780 13728 4808
rect 7469 4743 7527 4749
rect 6144 4712 6868 4740
rect 6144 4700 6150 4712
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5626 4672 5632 4684
rect 5583 4644 5632 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6840 4681 6868 4712
rect 7469 4709 7481 4743
rect 7515 4740 7527 4743
rect 10318 4740 10324 4752
rect 7515 4712 10324 4740
rect 7515 4709 7527 4712
rect 7469 4703 7527 4709
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 10778 4749 10784 4752
rect 10772 4740 10784 4749
rect 10739 4712 10784 4740
rect 10772 4703 10784 4712
rect 10778 4700 10784 4703
rect 10836 4700 10842 4752
rect 12268 4740 12296 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 17218 4808 17224 4820
rect 14148 4780 16528 4808
rect 17179 4780 17224 4808
rect 14148 4768 14154 4780
rect 10980 4712 12296 4740
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4641 6883 4675
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6825 4635 6883 4641
rect 6932 4644 7389 4672
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 6932 4604 6960 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8386 4672 8392 4684
rect 8343 4644 8392 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 5491 4576 5580 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 1596 4536 1624 4567
rect 2222 4536 2228 4548
rect 1596 4508 2228 4536
rect 2222 4496 2228 4508
rect 2280 4536 2286 4548
rect 2976 4536 3004 4567
rect 5552 4548 5580 4576
rect 5736 4576 6960 4604
rect 2280 4508 3004 4536
rect 2280 4496 2286 4508
rect 5534 4496 5540 4548
rect 5592 4496 5598 4548
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 3108 4440 3433 4468
rect 3108 4428 3114 4440
rect 3421 4437 3433 4440
rect 3467 4468 3479 4471
rect 3878 4468 3884 4480
rect 3467 4440 3884 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 4798 4468 4804 4480
rect 4571 4440 4804 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 4798 4428 4804 4440
rect 4856 4468 4862 4480
rect 5736 4468 5764 4576
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 7156 4576 7205 4604
rect 7156 4564 7162 4576
rect 7193 4573 7205 4576
rect 7239 4604 7251 4607
rect 7282 4604 7288 4616
rect 7239 4576 7288 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 7392 4604 7420 4635
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8754 4672 8760 4684
rect 8715 4644 8760 4672
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9398 4672 9404 4684
rect 9359 4644 9404 4672
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 10410 4672 10416 4684
rect 9907 4644 10416 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10410 4632 10416 4644
rect 10468 4672 10474 4684
rect 10980 4672 11008 4712
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 13136 4712 13676 4740
rect 13136 4700 13142 4712
rect 10468 4644 11008 4672
rect 10468 4632 10474 4644
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11974 4672 11980 4684
rect 11112 4644 11980 4672
rect 11112 4632 11118 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12308 4644 12357 4672
rect 12308 4632 12314 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 13170 4672 13176 4684
rect 12851 4644 13176 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 13648 4681 13676 4712
rect 15654 4700 15660 4752
rect 15712 4740 15718 4752
rect 16086 4743 16144 4749
rect 16086 4740 16098 4743
rect 15712 4712 16098 4740
rect 15712 4700 15718 4712
rect 16086 4709 16098 4712
rect 16132 4740 16144 4743
rect 16390 4740 16396 4752
rect 16132 4712 16396 4740
rect 16132 4709 16144 4712
rect 16086 4703 16144 4709
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 16500 4740 16528 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 21174 4749 21180 4752
rect 18693 4743 18751 4749
rect 18693 4740 18705 4743
rect 16500 4712 18705 4740
rect 18693 4709 18705 4712
rect 18739 4709 18751 4743
rect 18693 4703 18751 4709
rect 21116 4743 21180 4749
rect 21116 4709 21128 4743
rect 21162 4709 21180 4743
rect 21116 4703 21180 4709
rect 21174 4700 21180 4703
rect 21232 4700 21238 4752
rect 13633 4675 13691 4681
rect 13320 4644 13365 4672
rect 13320 4632 13326 4644
rect 13633 4641 13645 4675
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14424 4644 14565 4672
rect 14424 4632 14430 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15381 4675 15439 4681
rect 15381 4672 15393 4675
rect 14792 4644 15393 4672
rect 14792 4632 14798 4644
rect 15381 4641 15393 4644
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15620 4644 15853 4672
rect 15620 4632 15626 4644
rect 15841 4641 15853 4644
rect 15887 4672 15899 4675
rect 18506 4672 18512 4684
rect 15887 4644 18512 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 18506 4632 18512 4644
rect 18564 4672 18570 4684
rect 21361 4675 21419 4681
rect 21361 4672 21373 4675
rect 18564 4644 21373 4672
rect 18564 4632 18570 4644
rect 21361 4641 21373 4644
rect 21407 4641 21419 4675
rect 21361 4635 21419 4641
rect 9582 4604 9588 4616
rect 7392 4576 9588 4604
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10502 4604 10508 4616
rect 10008 4576 10508 4604
rect 10008 4564 10014 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 13354 4604 13360 4616
rect 12483 4576 13360 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 13464 4576 15025 4604
rect 6270 4496 6276 4548
rect 6328 4536 6334 4548
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 6328 4508 8125 4536
rect 6328 4496 6334 4508
rect 8113 4505 8125 4508
rect 8159 4505 8171 4539
rect 8113 4499 8171 4505
rect 9306 4496 9312 4548
rect 9364 4536 9370 4548
rect 9766 4536 9772 4548
rect 9364 4508 9772 4536
rect 9364 4496 9370 4508
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 11716 4508 12020 4536
rect 4856 4440 5764 4468
rect 4856 4428 4862 4440
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5868 4440 5917 4468
rect 5868 4428 5874 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 6362 4468 6368 4480
rect 6323 4440 6368 4468
rect 5905 4431 5963 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 11716 4468 11744 4508
rect 9456 4440 11744 4468
rect 9456 4428 9462 4440
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 11885 4471 11943 4477
rect 11885 4468 11897 4471
rect 11848 4440 11897 4468
rect 11848 4428 11854 4440
rect 11885 4437 11897 4440
rect 11931 4437 11943 4471
rect 11992 4468 12020 4508
rect 12158 4496 12164 4548
rect 12216 4536 12222 4548
rect 13081 4539 13139 4545
rect 13081 4536 13093 4539
rect 12216 4508 13093 4536
rect 12216 4496 12222 4508
rect 13081 4505 13093 4508
rect 13127 4505 13139 4539
rect 13081 4499 13139 4505
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 13464 4536 13492 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 15013 4567 15071 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 13228 4508 13492 4536
rect 13817 4539 13875 4545
rect 13228 4496 13234 4508
rect 13817 4505 13829 4539
rect 13863 4536 13875 4539
rect 15470 4536 15476 4548
rect 13863 4508 15476 4536
rect 13863 4505 13875 4508
rect 13817 4499 13875 4505
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 16776 4508 19993 4536
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 11992 4440 12449 4468
rect 11885 4431 11943 4437
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 12526 4428 12532 4480
rect 12584 4468 12590 4480
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 12584 4440 12633 4468
rect 12584 4428 12590 4440
rect 12621 4437 12633 4440
rect 12667 4437 12679 4471
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 12621 4431 12679 4437
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16776 4468 16804 4508
rect 19981 4505 19993 4508
rect 20027 4505 20039 4539
rect 19981 4499 20039 4505
rect 18046 4468 18052 4480
rect 16264 4440 16804 4468
rect 18007 4440 18052 4468
rect 16264 4428 16270 4440
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 18196 4440 18337 4468
rect 18196 4428 18202 4440
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18325 4431 18383 4437
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1581 4267 1639 4273
rect 1581 4233 1593 4267
rect 1627 4264 1639 4267
rect 2866 4264 2872 4276
rect 1627 4236 2872 4264
rect 1627 4233 1639 4236
rect 1581 4227 1639 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 4890 4264 4896 4276
rect 3620 4236 4896 4264
rect 1854 4128 1860 4140
rect 1504 4100 1860 4128
rect 1504 4069 1532 4100
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 3620 4128 3648 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 7006 4264 7012 4276
rect 5408 4236 7012 4264
rect 5408 4224 5414 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7340 4236 8033 4264
rect 7340 4224 7346 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 11054 4264 11060 4276
rect 8021 4227 8079 4233
rect 8128 4236 11060 4264
rect 4985 4199 5043 4205
rect 4985 4165 4997 4199
rect 5031 4196 5043 4199
rect 5031 4168 5856 4196
rect 5031 4165 5043 4168
rect 4985 4159 5043 4165
rect 5718 4128 5724 4140
rect 3528 4100 3648 4128
rect 5644 4100 5724 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4029 1547 4063
rect 1489 4023 1547 4029
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2222 4069 2228 4072
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1820 4032 1961 4060
rect 1820 4020 1826 4032
rect 1949 4029 1961 4032
rect 1995 4029 2007 4063
rect 2216 4060 2228 4069
rect 2183 4032 2228 4060
rect 1949 4023 2007 4029
rect 2216 4023 2228 4032
rect 1964 3992 1992 4023
rect 2222 4020 2228 4023
rect 2280 4020 2286 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 3528 4060 3556 4100
rect 2556 4032 3556 4060
rect 3605 4063 3663 4069
rect 2556 4020 2562 4032
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 4430 4060 4436 4072
rect 3651 4032 4436 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3620 3992 3648 4023
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 3850 3995 3908 4001
rect 3850 3992 3862 3995
rect 1964 3964 3648 3992
rect 3712 3964 3862 3992
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3712 3924 3740 3964
rect 3850 3961 3862 3964
rect 3896 3961 3908 3995
rect 3850 3955 3908 3961
rect 3384 3896 3740 3924
rect 5261 3927 5319 3933
rect 3384 3884 3390 3896
rect 5261 3893 5273 3927
rect 5307 3924 5319 3927
rect 5534 3924 5540 3936
rect 5307 3896 5540 3924
rect 5307 3893 5319 3896
rect 5261 3887 5319 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5644 3933 5672 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 5828 4128 5856 4168
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5828 4100 5917 4128
rect 5905 4097 5917 4100
rect 5951 4128 5963 4131
rect 5994 4128 6000 4140
rect 5951 4100 6000 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 8128 4137 8156 4236
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 14090 4264 14096 4276
rect 11164 4236 14096 4264
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 11164 4196 11192 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 16390 4264 16396 4276
rect 16351 4236 16396 4264
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 9824 4168 11192 4196
rect 9824 4156 9830 4168
rect 17218 4156 17224 4208
rect 17276 4196 17282 4208
rect 17865 4199 17923 4205
rect 17276 4168 17356 4196
rect 17276 4156 17282 4168
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 6512 4100 6653 4128
rect 6512 4088 6518 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 10781 4131 10839 4137
rect 8113 4091 8171 4097
rect 9600 4100 9904 4128
rect 9600 4072 9628 4100
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 9030 4060 9036 4072
rect 7708 4032 9036 4060
rect 7708 4020 7714 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 9766 4060 9772 4072
rect 9723 4032 9772 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9876 4060 9904 4100
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 11790 4128 11796 4140
rect 10827 4100 11796 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 11790 4088 11796 4100
rect 11848 4128 11854 4140
rect 13725 4131 13783 4137
rect 11848 4100 12020 4128
rect 11848 4088 11854 4100
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 9876 4032 10885 4060
rect 10873 4029 10885 4032
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11020 4032 11065 4060
rect 11624 4032 11897 4060
rect 11020 4020 11026 4032
rect 6914 4001 6920 4004
rect 6908 3992 6920 4001
rect 6875 3964 6920 3992
rect 6908 3955 6920 3964
rect 6914 3952 6920 3955
rect 6972 3952 6978 4004
rect 9432 3995 9490 4001
rect 9432 3961 9444 3995
rect 9478 3992 9490 3995
rect 10134 3992 10140 4004
rect 9478 3964 10140 3992
rect 9478 3961 9490 3964
rect 9432 3955 9490 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 11514 3992 11520 4004
rect 10652 3964 11520 3992
rect 10652 3952 10658 3964
rect 11514 3952 11520 3964
rect 11572 3992 11578 4004
rect 11624 3992 11652 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 11992 4060 12020 4100
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 13998 4128 14004 4140
rect 13771 4100 14004 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 17328 4137 17356 4168
rect 17865 4165 17877 4199
rect 17911 4196 17923 4199
rect 19242 4196 19248 4208
rect 17911 4168 19248 4196
rect 17911 4165 17923 4168
rect 17865 4159 17923 4165
rect 19242 4156 19248 4168
rect 19300 4156 19306 4208
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 21818 4128 21824 4140
rect 17460 4100 17505 4128
rect 20456 4100 21824 4128
rect 17460 4088 17466 4100
rect 12141 4063 12199 4069
rect 12141 4060 12153 4063
rect 11992 4032 12153 4060
rect 11885 4023 11943 4029
rect 12141 4029 12153 4032
rect 12187 4029 12199 4063
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 12141 4023 12199 4029
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15654 4060 15660 4072
rect 15059 4032 15660 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 17494 4060 17500 4072
rect 17455 4032 17500 4060
rect 17494 4020 17500 4032
rect 17552 4020 17558 4072
rect 17586 4020 17592 4072
rect 17644 4060 17650 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17644 4032 18153 4060
rect 17644 4020 17650 4032
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18598 4060 18604 4072
rect 18559 4032 18604 4060
rect 18141 4023 18199 4029
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 20456 4069 20484 4100
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 20211 4032 20453 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 20441 4023 20499 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 20588 4032 21097 4060
rect 20588 4020 20594 4032
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 21085 4023 21143 4029
rect 11572 3964 11652 3992
rect 11572 3952 11578 3964
rect 11698 3952 11704 4004
rect 11756 3992 11762 4004
rect 12618 3992 12624 4004
rect 11756 3964 12624 3992
rect 11756 3952 11762 3964
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 13906 3992 13912 4004
rect 13867 3964 13912 3992
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 15280 3995 15338 4001
rect 15280 3961 15292 3995
rect 15326 3992 15338 3995
rect 15930 3992 15936 4004
rect 15326 3964 15936 3992
rect 15326 3961 15338 3964
rect 15280 3955 15338 3961
rect 15930 3952 15936 3964
rect 15988 3952 15994 4004
rect 20714 3992 20720 4004
rect 20548 3964 20720 3992
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3924 5779 3927
rect 6730 3924 6736 3936
rect 5767 3896 6736 3924
rect 5767 3893 5779 3896
rect 5721 3887 5779 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 7156 3896 8125 3924
rect 7156 3884 7162 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 8294 3924 8300 3936
rect 8255 3896 8300 3924
rect 8113 3887 8171 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 8536 3896 9965 3924
rect 8536 3884 8542 3896
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 12802 3924 12808 3936
rect 11379 3896 12808 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13814 3924 13820 3936
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14274 3924 14280 3936
rect 14235 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 16022 3924 16028 3936
rect 14783 3896 16028 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18325 3927 18383 3933
rect 18325 3924 18337 3927
rect 18012 3896 18337 3924
rect 18012 3884 18018 3896
rect 18325 3893 18337 3896
rect 18371 3893 18383 3927
rect 18782 3924 18788 3936
rect 18743 3896 18788 3924
rect 18325 3887 18383 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19058 3924 19064 3936
rect 19019 3896 19064 3924
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 20548 3924 20576 3964
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 20898 3992 20904 4004
rect 20859 3964 20904 3992
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 19843 3896 20576 3924
rect 20625 3927 20683 3933
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 21358 3924 21364 3936
rect 20671 3896 21364 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1489 3723 1547 3729
rect 1489 3689 1501 3723
rect 1535 3720 1547 3723
rect 2222 3720 2228 3732
rect 1535 3692 2228 3720
rect 1535 3689 1547 3692
rect 1489 3683 1547 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 4062 3720 4068 3732
rect 2332 3692 4068 3720
rect 1026 3612 1032 3664
rect 1084 3652 1090 3664
rect 2332 3652 2360 3692
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 5166 3720 5172 3732
rect 4212 3692 5172 3720
rect 4212 3680 4218 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5902 3720 5908 3732
rect 5863 3692 5908 3720
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 6144 3692 6592 3720
rect 6144 3680 6150 3692
rect 1084 3624 2360 3652
rect 2624 3655 2682 3661
rect 1084 3612 1090 3624
rect 2624 3621 2636 3655
rect 2670 3652 2682 3655
rect 2866 3652 2872 3664
rect 2670 3624 2872 3652
rect 2670 3621 2682 3624
rect 2624 3615 2682 3621
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 5258 3652 5264 3664
rect 3200 3624 4108 3652
rect 3200 3612 3206 3624
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 3326 3584 3332 3596
rect 1544 3556 3188 3584
rect 3287 3556 3332 3584
rect 1544 3544 1550 3556
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 2958 3516 2964 3528
rect 2915 3488 2964 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3160 3516 3188 3556
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3878 3584 3884 3596
rect 3568 3556 3884 3584
rect 3568 3544 3574 3556
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 4080 3593 4108 3624
rect 4632 3624 5264 3652
rect 4057 3587 4115 3593
rect 4057 3553 4069 3587
rect 4103 3553 4115 3587
rect 4057 3547 4115 3553
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4488 3556 4537 3584
rect 4488 3544 4494 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 4338 3516 4344 3528
rect 3160 3488 4344 3516
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4632 3516 4660 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 5920 3652 5948 3680
rect 6426 3655 6484 3661
rect 6426 3652 6438 3655
rect 5920 3624 6438 3652
rect 6426 3621 6438 3624
rect 6472 3621 6484 3655
rect 6564 3652 6592 3692
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7374 3720 7380 3732
rect 7064 3692 7380 3720
rect 7064 3680 7070 3692
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 8260 3692 8401 3720
rect 8260 3680 8266 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8389 3683 8447 3689
rect 8496 3692 9137 3720
rect 8496 3652 8524 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9732 3692 10057 3720
rect 9732 3680 9738 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10284 3692 10701 3720
rect 10284 3680 10290 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 12066 3720 12072 3732
rect 10836 3692 12072 3720
rect 10836 3680 10842 3692
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 15654 3720 15660 3732
rect 15304 3692 15660 3720
rect 6564 3624 8524 3652
rect 6426 3615 6484 3621
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 11606 3652 11612 3664
rect 9088 3624 11612 3652
rect 9088 3612 9094 3624
rect 4792 3587 4850 3593
rect 4792 3553 4804 3587
rect 4838 3584 4850 3587
rect 5994 3584 6000 3596
rect 4838 3556 6000 3584
rect 4838 3553 4850 3556
rect 4792 3547 4850 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 9766 3584 9772 3596
rect 6104 3556 9772 3584
rect 4448 3488 4660 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 624 3420 1716 3448
rect 624 3408 630 3420
rect 1688 3380 1716 3420
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4448 3448 4476 3488
rect 3844 3420 4476 3448
rect 3844 3408 3850 3420
rect 3050 3380 3056 3392
rect 1688 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3234 3380 3240 3392
rect 3195 3352 3240 3380
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 4249 3383 4307 3389
rect 4249 3349 4261 3383
rect 4295 3380 4307 3383
rect 6104 3380 6132 3556
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10888 3593 10916 3624
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 12888 3655 12946 3661
rect 12888 3621 12900 3655
rect 12934 3652 12946 3655
rect 13262 3652 13268 3664
rect 12934 3624 13268 3652
rect 12934 3621 12946 3624
rect 12888 3615 12946 3621
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 14016 3652 14044 3680
rect 14798 3655 14856 3661
rect 14798 3652 14810 3655
rect 14016 3624 14810 3652
rect 14798 3621 14810 3624
rect 14844 3621 14856 3655
rect 14798 3615 14856 3621
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 10100 3556 10149 3584
rect 10100 3544 10106 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3553 10931 3587
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 10873 3547 10931 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11701 3587 11759 3593
rect 11701 3553 11713 3587
rect 11747 3553 11759 3587
rect 11701 3547 11759 3553
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 8570 3516 8576 3528
rect 8527 3488 8576 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 4295 3352 6132 3380
rect 6196 3380 6224 3479
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9674 3516 9680 3528
rect 8987 3488 9680 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 8680 3448 8708 3479
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 11716 3516 11744 3547
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 13354 3584 13360 3596
rect 12124 3556 13360 3584
rect 12124 3544 12130 3556
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 15304 3584 15332 3692
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15930 3720 15936 3732
rect 15891 3692 15936 3720
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 19061 3723 19119 3729
rect 19061 3689 19073 3723
rect 19107 3689 19119 3723
rect 19061 3683 19119 3689
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 16393 3655 16451 3661
rect 16393 3652 16405 3655
rect 15620 3624 16405 3652
rect 15620 3612 15626 3624
rect 16393 3621 16405 3624
rect 16439 3621 16451 3655
rect 19076 3652 19104 3683
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 21177 3723 21235 3729
rect 21177 3720 21189 3723
rect 20680 3692 21189 3720
rect 20680 3680 20686 3692
rect 21177 3689 21189 3692
rect 21223 3689 21235 3723
rect 21177 3683 21235 3689
rect 16393 3615 16451 3621
rect 17696 3624 19104 3652
rect 14599 3556 15332 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 17696 3593 17724 3624
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 20257 3655 20315 3661
rect 20257 3652 20269 3655
rect 19392 3624 20269 3652
rect 19392 3612 19398 3624
rect 20257 3621 20269 3624
rect 20303 3621 20315 3655
rect 20806 3652 20812 3664
rect 20767 3624 20812 3652
rect 20257 3615 20315 3621
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 15436 3556 17417 3584
rect 15436 3544 15442 3556
rect 17405 3553 17417 3556
rect 17451 3553 17463 3587
rect 17405 3547 17463 3553
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 17920 3556 18153 3584
rect 17920 3544 17926 3556
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 18748 3556 18797 3584
rect 18748 3544 18754 3556
rect 18785 3553 18797 3556
rect 18831 3553 18843 3587
rect 19242 3584 19248 3596
rect 19203 3556 19248 3584
rect 18785 3547 18843 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 21358 3584 21364 3596
rect 21319 3556 21364 3584
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 12342 3516 12348 3528
rect 11256 3488 11744 3516
rect 12303 3488 12348 3516
rect 10244 3448 10272 3476
rect 7432 3420 8616 3448
rect 8680 3420 10272 3448
rect 7432 3408 7438 3420
rect 6454 3380 6460 3392
rect 6196 3352 6460 3380
rect 4295 3349 4307 3352
rect 4249 3343 4307 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 6972 3352 7573 3380
rect 6972 3340 6978 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 8021 3383 8079 3389
rect 8021 3380 8033 3383
rect 7984 3352 8033 3380
rect 7984 3340 7990 3352
rect 8021 3349 8033 3352
rect 8067 3349 8079 3383
rect 8588 3380 8616 3420
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8588 3352 8953 3380
rect 8021 3343 8079 3349
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 9858 3380 9864 3392
rect 9723 3352 9864 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 11256 3380 11284 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 16758 3516 16764 3528
rect 16719 3488 16764 3516
rect 12621 3479 12679 3485
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 12636 3448 12664 3479
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 11572 3420 12664 3448
rect 11572 3408 11578 3420
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 16209 3451 16267 3457
rect 16209 3448 16221 3451
rect 16172 3420 16221 3448
rect 16172 3408 16178 3420
rect 16209 3417 16221 3420
rect 16255 3417 16267 3451
rect 16209 3411 16267 3417
rect 18325 3451 18383 3457
rect 18325 3417 18337 3451
rect 18371 3448 18383 3451
rect 19242 3448 19248 3460
rect 18371 3420 19248 3448
rect 18371 3417 18383 3420
rect 18325 3411 18383 3417
rect 19242 3408 19248 3420
rect 19300 3408 19306 3460
rect 20070 3448 20076 3460
rect 20031 3420 20076 3448
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 20530 3408 20536 3460
rect 20588 3448 20594 3460
rect 20625 3451 20683 3457
rect 20625 3448 20637 3451
rect 20588 3420 20637 3448
rect 20588 3408 20594 3420
rect 20625 3417 20637 3420
rect 20671 3417 20683 3451
rect 20625 3411 20683 3417
rect 10008 3352 11284 3380
rect 11333 3383 11391 3389
rect 10008 3340 10014 3352
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11790 3380 11796 3392
rect 11379 3352 11796 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 13538 3380 13544 3392
rect 11931 3352 13544 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 17310 3380 17316 3392
rect 17267 3352 17316 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17865 3383 17923 3389
rect 17865 3349 17877 3383
rect 17911 3380 17923 3383
rect 18138 3380 18144 3392
rect 17911 3352 18144 3380
rect 17911 3349 17923 3352
rect 17865 3343 17923 3349
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 18598 3380 18604 3392
rect 18559 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19797 3383 19855 3389
rect 19797 3349 19809 3383
rect 19843 3380 19855 3383
rect 21358 3380 21364 3392
rect 19843 3352 21364 3380
rect 19843 3349 19855 3352
rect 19797 3343 19855 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1765 3179 1823 3185
rect 1765 3176 1777 3179
rect 1728 3148 1777 3176
rect 1728 3136 1734 3148
rect 1765 3145 1777 3148
rect 1811 3145 1823 3179
rect 1765 3139 1823 3145
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2832 3148 2881 3176
rect 2832 3136 2838 3148
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 4798 3176 4804 3188
rect 3099 3148 4804 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5000 3148 7696 3176
rect 2961 3111 3019 3117
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 3007 3080 3556 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2866 3040 2872 3052
rect 2363 3012 2872 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2866 3000 2872 3012
rect 2924 3040 2930 3052
rect 3234 3040 3240 3052
rect 2924 3012 3240 3040
rect 2924 3000 2930 3012
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 3418 2972 3424 2984
rect 1719 2944 3424 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3528 2972 3556 3080
rect 5000 3040 5028 3148
rect 5169 3111 5227 3117
rect 5169 3077 5181 3111
rect 5215 3108 5227 3111
rect 6454 3108 6460 3120
rect 5215 3080 6460 3108
rect 5215 3077 5227 3080
rect 5169 3071 5227 3077
rect 6454 3068 6460 3080
rect 6512 3068 6518 3120
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 7466 3108 7472 3120
rect 6696 3080 7472 3108
rect 6696 3068 6702 3080
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 4448 3012 5028 3040
rect 5077 3043 5135 3049
rect 3970 2972 3976 2984
rect 3528 2944 3976 2972
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4269 2975 4327 2981
rect 4269 2941 4281 2975
rect 4315 2972 4327 2975
rect 4448 2972 4476 3012
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5442 3040 5448 3052
rect 5123 3012 5448 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5902 3040 5908 3052
rect 5583 3012 5908 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 5994 3000 6000 3052
rect 6052 3040 6058 3052
rect 7282 3040 7288 3052
rect 6052 3012 7288 3040
rect 6052 3000 6058 3012
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 4315 2944 4476 2972
rect 4315 2941 4327 2944
rect 4269 2935 4327 2941
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 4580 2944 5181 2972
rect 4580 2932 4586 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6730 2972 6736 2984
rect 5767 2944 6736 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 3053 2907 3111 2913
rect 3053 2904 3065 2907
rect 2455 2876 3065 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 3053 2873 3065 2876
rect 3099 2873 3111 2907
rect 5534 2904 5540 2916
rect 3053 2867 3111 2873
rect 3344 2876 5540 2904
rect 3344 2848 3372 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5629 2907 5687 2913
rect 5629 2873 5641 2907
rect 5675 2904 5687 2907
rect 7006 2904 7012 2916
rect 5675 2876 6684 2904
rect 6967 2876 7012 2904
rect 5675 2873 5687 2876
rect 5629 2867 5687 2873
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1578 2836 1584 2848
rect 256 2808 1584 2836
rect 256 2796 262 2808
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 2501 2839 2559 2845
rect 2501 2805 2513 2839
rect 2547 2836 2559 2839
rect 2961 2839 3019 2845
rect 2961 2836 2973 2839
rect 2547 2808 2973 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 2961 2805 2973 2808
rect 3007 2805 3019 2839
rect 2961 2799 3019 2805
rect 3145 2839 3203 2845
rect 3145 2805 3157 2839
rect 3191 2836 3203 2839
rect 3234 2836 3240 2848
rect 3191 2808 3240 2836
rect 3191 2805 3203 2808
rect 3145 2799 3203 2805
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 3326 2796 3332 2848
rect 3384 2796 3390 2848
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 5902 2836 5908 2848
rect 3752 2808 5908 2836
rect 3752 2796 3758 2808
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6086 2836 6092 2848
rect 6047 2808 6092 2836
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 6656 2845 6684 2876
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2805 6699 2839
rect 7668 2836 7696 3148
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 13265 3179 13323 3185
rect 9824 3148 10088 3176
rect 9824 3136 9830 3148
rect 8573 3111 8631 3117
rect 8573 3108 8585 3111
rect 7760 3080 8585 3108
rect 7760 3049 7788 3080
rect 8573 3077 8585 3080
rect 8619 3077 8631 3111
rect 10060 3108 10088 3148
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 14642 3176 14648 3188
rect 13311 3148 14648 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 15841 3179 15899 3185
rect 15841 3145 15853 3179
rect 15887 3176 15899 3179
rect 17586 3176 17592 3188
rect 15887 3148 17592 3176
rect 15887 3145 15899 3148
rect 15841 3139 15899 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 11054 3108 11060 3120
rect 10060 3080 11060 3108
rect 8573 3071 8631 3077
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 13170 3108 13176 3120
rect 11388 3080 13176 3108
rect 11388 3068 11394 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13630 3068 13636 3120
rect 13688 3108 13694 3120
rect 13688 3080 20576 3108
rect 13688 3068 13694 3080
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7926 3040 7932 3052
rect 7887 3012 7932 3040
rect 7745 3003 7803 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10594 3040 10600 3052
rect 10091 3012 10600 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 13262 3040 13268 3052
rect 12759 3012 13268 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8478 2972 8484 2984
rect 8067 2944 8484 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10744 2944 10793 2972
rect 10744 2932 10750 2944
rect 10781 2941 10793 2944
rect 10827 2972 10839 2975
rect 10870 2972 10876 2984
rect 10827 2944 10876 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 9674 2904 9680 2916
rect 8260 2876 9680 2904
rect 8260 2864 8266 2876
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 9800 2907 9858 2913
rect 9800 2873 9812 2907
rect 9846 2904 9858 2907
rect 10226 2904 10232 2916
rect 9846 2876 10232 2904
rect 9846 2873 9858 2876
rect 9800 2867 9858 2873
rect 10226 2864 10232 2876
rect 10284 2904 10290 2916
rect 10980 2904 11008 3003
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 15289 3043 15347 3049
rect 14332 3012 14872 3040
rect 14332 3000 14338 3012
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11848 2944 11897 2972
rect 11848 2932 11854 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12400 2944 12909 2972
rect 12400 2932 12406 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 12897 2935 12955 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13780 2944 14013 2972
rect 13780 2932 13786 2944
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2972 14703 2975
rect 14734 2972 14740 2984
rect 14691 2944 14740 2972
rect 14691 2941 14703 2944
rect 14645 2935 14703 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14844 2972 14872 3012
rect 15289 3009 15301 3043
rect 15335 3040 15347 3043
rect 15930 3040 15936 3052
rect 15335 3012 15936 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 20548 3049 20576 3080
rect 20533 3043 20591 3049
rect 17000 3012 17908 3040
rect 17000 3000 17006 3012
rect 15381 2975 15439 2981
rect 15381 2972 15393 2975
rect 14844 2944 15393 2972
rect 15381 2941 15393 2944
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 16758 2972 16764 2984
rect 15519 2944 16764 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 17880 2981 17908 3012
rect 20533 3009 20545 3043
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 18012 2944 18337 2972
rect 18012 2932 18018 2944
rect 18325 2941 18337 2944
rect 18371 2941 18383 2975
rect 18782 2972 18788 2984
rect 18743 2944 18788 2972
rect 18325 2935 18383 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19426 2972 19432 2984
rect 19383 2944 19432 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19886 2972 19892 2984
rect 19847 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 20772 2944 21189 2972
rect 20772 2932 20778 2944
rect 21177 2941 21189 2944
rect 21223 2972 21235 2975
rect 22738 2972 22744 2984
rect 21223 2944 22744 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 14829 2907 14887 2913
rect 10284 2876 14780 2904
rect 10284 2864 10290 2876
rect 8294 2836 8300 2848
rect 7668 2808 8300 2836
rect 6641 2799 6699 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8478 2836 8484 2848
rect 8435 2808 8484 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8619 2808 8677 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 8665 2805 8677 2808
rect 8711 2836 8723 2839
rect 10042 2836 10048 2848
rect 8711 2808 10048 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10192 2808 10333 2836
rect 10192 2796 10198 2808
rect 10321 2805 10333 2808
rect 10367 2805 10379 2839
rect 10686 2836 10692 2848
rect 10647 2808 10692 2836
rect 10321 2799 10379 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11882 2836 11888 2848
rect 10928 2808 11888 2836
rect 10928 2796 10934 2808
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12710 2836 12716 2848
rect 12115 2808 12716 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 13725 2839 13783 2845
rect 12860 2808 12905 2836
rect 12860 2796 12866 2808
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 13814 2836 13820 2848
rect 13771 2808 13820 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14182 2836 14188 2848
rect 14143 2808 14188 2836
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 14752 2836 14780 2876
rect 14829 2873 14841 2907
rect 14875 2904 14887 2907
rect 15194 2904 15200 2916
rect 14875 2876 15200 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 16117 2907 16175 2913
rect 16117 2904 16129 2907
rect 15712 2876 16129 2904
rect 15712 2864 15718 2876
rect 16117 2873 16129 2876
rect 16163 2873 16175 2907
rect 16117 2867 16175 2873
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2873 16359 2907
rect 16301 2867 16359 2873
rect 16206 2836 16212 2848
rect 14752 2808 16212 2836
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16316 2836 16344 2867
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 17129 2907 17187 2913
rect 17129 2904 17141 2907
rect 16540 2876 17141 2904
rect 16540 2864 16546 2876
rect 17129 2873 17141 2876
rect 17175 2873 17187 2907
rect 19150 2904 19156 2916
rect 19111 2876 19156 2904
rect 17129 2867 17187 2873
rect 19150 2864 19156 2876
rect 19208 2864 19214 2916
rect 19610 2864 19616 2916
rect 19668 2904 19674 2916
rect 19705 2907 19763 2913
rect 19705 2904 19717 2907
rect 19668 2876 19717 2904
rect 19668 2864 19674 2876
rect 19705 2873 19717 2876
rect 19751 2873 19763 2907
rect 19705 2867 19763 2873
rect 17681 2839 17739 2845
rect 17681 2836 17693 2839
rect 16316 2808 17693 2836
rect 17681 2805 17693 2808
rect 17727 2805 17739 2839
rect 17681 2799 17739 2805
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 18141 2839 18199 2845
rect 18141 2836 18153 2839
rect 18012 2808 18153 2836
rect 18012 2796 18018 2808
rect 18141 2805 18153 2808
rect 18187 2805 18199 2839
rect 18598 2836 18604 2848
rect 18559 2808 18604 2836
rect 18141 2799 18199 2805
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2682 2632 2688 2644
rect 2643 2604 2688 2632
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 4062 2632 4068 2644
rect 3099 2604 4068 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5074 2632 5080 2644
rect 4755 2604 5080 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7190 2632 7196 2644
rect 7151 2604 7196 2632
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 8849 2635 8907 2641
rect 8849 2601 8861 2635
rect 8895 2601 8907 2635
rect 9858 2632 9864 2644
rect 9819 2604 9864 2632
rect 8849 2595 8907 2601
rect 1578 2524 1584 2576
rect 1636 2564 1642 2576
rect 1673 2567 1731 2573
rect 1673 2564 1685 2567
rect 1636 2536 1685 2564
rect 1636 2524 1642 2536
rect 1673 2533 1685 2536
rect 1719 2533 1731 2567
rect 1673 2527 1731 2533
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 3878 2564 3884 2576
rect 2455 2536 3884 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 5721 2567 5779 2573
rect 4028 2536 4844 2564
rect 4028 2524 4034 2536
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 2958 2496 2964 2508
rect 2271 2468 2964 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3191 2468 3740 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 1857 2363 1915 2369
rect 1857 2329 1869 2363
rect 1903 2360 1915 2363
rect 3160 2360 3188 2459
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3292 2400 3337 2428
rect 3292 2388 3298 2400
rect 1903 2332 3188 2360
rect 3712 2360 3740 2468
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4816 2505 4844 2536
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 6086 2564 6092 2576
rect 5767 2536 6092 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 6086 2524 6092 2536
rect 6144 2524 6150 2576
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 7374 2564 7380 2576
rect 7147 2536 7380 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 8864 2564 8892 2595
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10134 2632 10140 2644
rect 9999 2604 10140 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 11146 2632 11152 2644
rect 10428 2604 11152 2632
rect 10428 2564 10456 2604
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12253 2635 12311 2641
rect 12253 2601 12265 2635
rect 12299 2601 12311 2635
rect 12253 2595 12311 2601
rect 12345 2635 12403 2641
rect 12345 2601 12357 2635
rect 12391 2632 12403 2635
rect 20257 2635 20315 2641
rect 12391 2604 20116 2632
rect 12391 2601 12403 2604
rect 12345 2595 12403 2601
rect 8864 2536 10456 2564
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 12268 2564 12296 2595
rect 12710 2564 12716 2576
rect 11112 2536 12112 2564
rect 12268 2536 12434 2564
rect 12671 2536 12716 2564
rect 11112 2524 11118 2536
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4120 2468 4261 2496
rect 4120 2456 4126 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 4890 2496 4896 2508
rect 4847 2468 4896 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 6236 2468 7757 2496
rect 6236 2456 6242 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 7852 2468 9628 2496
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 6914 2428 6920 2440
rect 5675 2400 6920 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7282 2428 7288 2440
rect 7243 2400 7288 2428
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 3712 2332 6316 2360
rect 1903 2329 1915 2332
rect 1857 2323 1915 2329
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 2648 2264 4169 2292
rect 2648 2252 2654 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 6178 2292 6184 2304
rect 6139 2264 6184 2292
rect 4157 2255 4215 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 6288 2292 6316 2332
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 7852 2360 7880 2468
rect 8294 2428 8300 2440
rect 8255 2400 8300 2428
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8435 2400 9536 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 9508 2369 9536 2400
rect 6420 2332 7880 2360
rect 9493 2363 9551 2369
rect 6420 2320 6426 2332
rect 9493 2329 9505 2363
rect 9539 2329 9551 2363
rect 9600 2360 9628 2468
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 9732 2468 10701 2496
rect 9732 2456 9738 2468
rect 10689 2465 10701 2468
rect 10735 2496 10747 2499
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10735 2468 10977 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 12084 2505 12112 2536
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 11296 2468 11345 2496
rect 11296 2456 11302 2468
rect 11333 2465 11345 2468
rect 11379 2465 11391 2499
rect 11333 2459 11391 2465
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2465 12127 2499
rect 12406 2496 12434 2536
rect 12710 2524 12716 2536
rect 12768 2524 12774 2576
rect 13814 2564 13820 2576
rect 13775 2536 13820 2564
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 14182 2524 14188 2576
rect 14240 2564 14246 2576
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14240 2536 14933 2564
rect 14240 2524 14246 2536
rect 14921 2533 14933 2536
rect 14967 2533 14979 2567
rect 15470 2564 15476 2576
rect 15431 2536 15476 2564
rect 14921 2527 14979 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 16022 2564 16028 2576
rect 15983 2536 16028 2564
rect 16022 2524 16028 2536
rect 16080 2524 16086 2576
rect 17589 2567 17647 2573
rect 17589 2533 17601 2567
rect 17635 2564 17647 2567
rect 17954 2564 17960 2576
rect 17635 2536 17960 2564
rect 17635 2533 17647 2536
rect 17589 2527 17647 2533
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 18138 2564 18144 2576
rect 18099 2536 18144 2564
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 18693 2567 18751 2573
rect 18693 2564 18705 2567
rect 18656 2536 18705 2564
rect 18656 2524 18662 2536
rect 18693 2533 18705 2536
rect 18739 2533 18751 2567
rect 19242 2564 19248 2576
rect 19203 2536 19248 2564
rect 18693 2527 18751 2533
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 12406 2468 13277 2496
rect 12069 2459 12127 2465
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13265 2459 13323 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 18506 2496 18512 2508
rect 16715 2468 18512 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 20088 2505 20116 2604
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20346 2632 20352 2644
rect 20303 2604 20352 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 20622 2564 20628 2576
rect 20583 2536 20628 2564
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 20073 2499 20131 2505
rect 20073 2465 20085 2499
rect 20119 2465 20131 2499
rect 20073 2459 20131 2465
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 21358 2496 21364 2508
rect 21315 2468 21364 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 21358 2456 21364 2468
rect 21416 2456 21422 2508
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 10152 2400 12357 2428
rect 10152 2360 10180 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 16899 2400 18552 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 9600 2332 10180 2360
rect 11517 2363 11575 2369
rect 9493 2323 9551 2329
rect 11517 2329 11529 2363
rect 11563 2360 11575 2363
rect 12526 2360 12532 2372
rect 11563 2332 12434 2360
rect 12487 2332 12532 2360
rect 11563 2329 11575 2332
rect 11517 2323 11575 2329
rect 7006 2292 7012 2304
rect 6288 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7558 2252 7564 2304
rect 7616 2292 7622 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 7616 2264 10517 2292
rect 7616 2252 7622 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 12406 2292 12434 2332
rect 12526 2320 12532 2332
rect 12584 2320 12590 2372
rect 12986 2320 12992 2372
rect 13044 2360 13050 2372
rect 13081 2363 13139 2369
rect 13081 2360 13093 2363
rect 13044 2332 13093 2360
rect 13044 2320 13050 2332
rect 13081 2329 13093 2332
rect 13127 2329 13139 2363
rect 13081 2323 13139 2329
rect 13446 2320 13452 2372
rect 13504 2360 13510 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13504 2332 13645 2360
rect 13504 2320 13510 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13633 2323 13691 2329
rect 13906 2320 13912 2372
rect 13964 2360 13970 2372
rect 14737 2363 14795 2369
rect 14737 2360 14749 2363
rect 13964 2332 14749 2360
rect 13964 2320 13970 2332
rect 14737 2329 14749 2332
rect 14783 2329 14795 2363
rect 14737 2323 14795 2329
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 15841 2363 15899 2369
rect 15841 2360 15853 2363
rect 14884 2332 15853 2360
rect 14884 2320 14890 2332
rect 15841 2329 15853 2332
rect 15887 2329 15899 2363
rect 15841 2323 15899 2329
rect 16942 2320 16948 2372
rect 17000 2360 17006 2372
rect 17405 2363 17463 2369
rect 17405 2360 17417 2363
rect 17000 2332 17417 2360
rect 17000 2320 17006 2332
rect 17405 2329 17417 2332
rect 17451 2329 17463 2363
rect 17405 2323 17463 2329
rect 17494 2320 17500 2372
rect 17552 2360 17558 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17552 2332 17969 2360
rect 17552 2320 17558 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 18524 2360 18552 2400
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 18656 2400 19073 2428
rect 18656 2388 18662 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 18690 2360 18696 2372
rect 18524 2332 18696 2360
rect 17957 2323 18015 2329
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 20809 2363 20867 2369
rect 20809 2329 20821 2363
rect 20855 2360 20867 2363
rect 22278 2360 22284 2372
rect 20855 2332 22284 2360
rect 20855 2329 20867 2332
rect 20809 2323 20867 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 13722 2292 13728 2304
rect 12406 2264 13728 2292
rect 10505 2255 10563 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 14332 2264 15393 2292
rect 14332 2252 14338 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18601 2295 18659 2301
rect 18601 2292 18613 2295
rect 17920 2264 18613 2292
rect 17920 2252 17926 2264
rect 18601 2261 18613 2264
rect 18647 2261 18659 2295
rect 21174 2292 21180 2304
rect 21135 2264 21180 2292
rect 18601 2255 18659 2261
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 6178 2048 6184 2100
rect 6236 2088 6242 2100
rect 9950 2088 9956 2100
rect 6236 2060 9956 2088
rect 6236 2048 6242 2060
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 10060 2060 14044 2088
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 10060 2020 10088 2060
rect 13909 2023 13967 2029
rect 13909 2020 13921 2023
rect 4120 1992 10088 2020
rect 10152 1992 13921 2020
rect 4120 1980 4126 1992
rect 4890 1912 4896 1964
rect 4948 1952 4954 1964
rect 10152 1952 10180 1992
rect 13909 1989 13921 1992
rect 13955 1989 13967 2023
rect 14016 2020 14044 2060
rect 16666 2048 16672 2100
rect 16724 2088 16730 2100
rect 21174 2088 21180 2100
rect 16724 2060 21180 2088
rect 16724 2048 16730 2060
rect 21174 2048 21180 2060
rect 21232 2048 21238 2100
rect 18046 2020 18052 2032
rect 14016 1992 18052 2020
rect 13909 1983 13967 1989
rect 18046 1980 18052 1992
rect 18104 1980 18110 2032
rect 4948 1924 10180 1952
rect 4948 1912 4954 1924
rect 10318 1912 10324 1964
rect 10376 1952 10382 1964
rect 12250 1952 12256 1964
rect 10376 1924 12256 1952
rect 10376 1912 10382 1924
rect 12250 1912 12256 1924
rect 12308 1912 12314 1964
rect 16574 1952 16580 1964
rect 12406 1924 16580 1952
rect 2958 1844 2964 1896
rect 3016 1884 3022 1896
rect 12406 1884 12434 1924
rect 16574 1912 16580 1924
rect 16632 1912 16638 1964
rect 3016 1856 12434 1884
rect 13909 1887 13967 1893
rect 3016 1844 3022 1856
rect 13909 1853 13921 1887
rect 13955 1884 13967 1887
rect 19058 1884 19064 1896
rect 13955 1856 19064 1884
rect 13955 1853 13967 1856
rect 13909 1847 13967 1853
rect 19058 1844 19064 1856
rect 19116 1844 19122 1896
rect 4154 1776 4160 1828
rect 4212 1816 4218 1828
rect 8386 1816 8392 1828
rect 4212 1788 8392 1816
rect 4212 1776 4218 1788
rect 8386 1776 8392 1788
rect 8444 1776 8450 1828
rect 4982 1708 4988 1760
rect 5040 1748 5046 1760
rect 6546 1748 6552 1760
rect 5040 1720 6552 1748
rect 5040 1708 5046 1720
rect 6546 1708 6552 1720
rect 6604 1708 6610 1760
rect 2774 1368 2780 1420
rect 2832 1408 2838 1420
rect 3786 1408 3792 1420
rect 2832 1380 3792 1408
rect 2832 1368 2838 1380
rect 3786 1368 3792 1380
rect 3844 1368 3850 1420
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2780 20476 2832 20528
rect 3240 20519 3292 20528
rect 3240 20485 3249 20519
rect 3249 20485 3283 20519
rect 3283 20485 3292 20519
rect 3240 20476 3292 20485
rect 4068 20519 4120 20528
rect 4068 20485 4077 20519
rect 4077 20485 4111 20519
rect 4111 20485 4120 20519
rect 4068 20476 4120 20485
rect 2872 20408 2924 20460
rect 2136 20315 2188 20324
rect 2136 20281 2145 20315
rect 2145 20281 2179 20315
rect 2179 20281 2188 20315
rect 2136 20272 2188 20281
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 2872 20315 2924 20324
rect 2872 20281 2881 20315
rect 2881 20281 2915 20315
rect 2915 20281 2924 20315
rect 2872 20272 2924 20281
rect 3424 20315 3476 20324
rect 3424 20281 3433 20315
rect 3433 20281 3467 20315
rect 3467 20281 3476 20315
rect 3424 20272 3476 20281
rect 10600 20272 10652 20324
rect 2780 20204 2832 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2228 20043 2280 20052
rect 2228 20009 2237 20043
rect 2237 20009 2271 20043
rect 2271 20009 2280 20043
rect 2228 20000 2280 20009
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 2964 20000 3016 20052
rect 2228 19864 2280 19916
rect 2596 19864 2648 19916
rect 4068 19864 4120 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 2596 19456 2648 19465
rect 3424 19456 3476 19508
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 1768 19227 1820 19236
rect 1768 19193 1777 19227
rect 1777 19193 1811 19227
rect 1811 19193 1820 19227
rect 1768 19184 1820 19193
rect 2964 19252 3016 19304
rect 3608 19252 3660 19304
rect 8576 19252 8628 19304
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1768 18912 1820 18964
rect 2228 18912 2280 18964
rect 2964 18912 3016 18964
rect 3608 18912 3660 18964
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 1584 18887 1636 18896
rect 1584 18853 1593 18887
rect 1593 18853 1627 18887
rect 1627 18853 1636 18887
rect 1584 18844 1636 18853
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 3148 18776 3200 18828
rect 8668 18844 8720 18896
rect 3056 18708 3108 18760
rect 9588 18776 9640 18828
rect 11244 18776 11296 18828
rect 6828 18708 6880 18760
rect 4068 18683 4120 18692
rect 4068 18649 4077 18683
rect 4077 18649 4111 18683
rect 4111 18649 4120 18683
rect 4068 18640 4120 18649
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 9588 18411 9640 18420
rect 9588 18377 9597 18411
rect 9597 18377 9631 18411
rect 9631 18377 9640 18411
rect 9588 18368 9640 18377
rect 1768 18300 1820 18352
rect 10232 18275 10284 18284
rect 10232 18241 10241 18275
rect 10241 18241 10275 18275
rect 10275 18241 10284 18275
rect 10232 18232 10284 18241
rect 2872 18207 2924 18216
rect 2872 18173 2881 18207
rect 2881 18173 2915 18207
rect 2915 18173 2924 18207
rect 2872 18164 2924 18173
rect 9864 18164 9916 18216
rect 1768 18139 1820 18148
rect 1768 18105 1777 18139
rect 1777 18105 1811 18139
rect 1811 18105 1820 18139
rect 1768 18096 1820 18105
rect 2320 18139 2372 18148
rect 2320 18105 2329 18139
rect 2329 18105 2363 18139
rect 2363 18105 2372 18139
rect 2320 18096 2372 18105
rect 11060 18096 11112 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 7288 18028 7340 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1768 17824 1820 17876
rect 2872 17824 2924 17876
rect 3056 17867 3108 17876
rect 3056 17833 3065 17867
rect 3065 17833 3099 17867
rect 3099 17833 3108 17867
rect 3056 17824 3108 17833
rect 6920 17824 6972 17876
rect 7288 17867 7340 17876
rect 7288 17833 7297 17867
rect 7297 17833 7331 17867
rect 7331 17833 7340 17867
rect 7288 17824 7340 17833
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 2504 17688 2556 17740
rect 5540 17731 5592 17740
rect 5540 17697 5574 17731
rect 5574 17697 5592 17731
rect 6828 17756 6880 17808
rect 10232 17824 10284 17876
rect 10876 17824 10928 17876
rect 11244 17867 11296 17876
rect 11244 17833 11253 17867
rect 11253 17833 11287 17867
rect 11287 17833 11296 17867
rect 11244 17824 11296 17833
rect 9772 17756 9824 17808
rect 5540 17688 5592 17697
rect 7012 17688 7064 17740
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 9128 17688 9180 17740
rect 11888 17688 11940 17740
rect 4804 17620 4856 17672
rect 7380 17663 7432 17672
rect 7380 17629 7389 17663
rect 7389 17629 7423 17663
rect 7423 17629 7432 17663
rect 7380 17620 7432 17629
rect 8392 17663 8444 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 3700 17484 3752 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 9496 17620 9548 17672
rect 6644 17484 6696 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1768 17280 1820 17332
rect 2320 17280 2372 17332
rect 5540 17280 5592 17332
rect 7380 17323 7432 17332
rect 2504 17212 2556 17264
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 13636 17144 13688 17196
rect 21364 17187 21416 17196
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 1768 17051 1820 17060
rect 1768 17017 1777 17051
rect 1777 17017 1811 17051
rect 1811 17017 1820 17051
rect 1768 17008 1820 17017
rect 2964 17076 3016 17128
rect 3700 17119 3752 17128
rect 3700 17085 3709 17119
rect 3709 17085 3743 17119
rect 3743 17085 3752 17119
rect 3700 17076 3752 17085
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 9496 17076 9548 17128
rect 21364 17153 21373 17187
rect 21373 17153 21407 17187
rect 21407 17153 21416 17187
rect 21364 17144 21416 17153
rect 2872 16940 2924 16992
rect 4068 17008 4120 17060
rect 4804 17008 4856 17060
rect 7288 17008 7340 17060
rect 8944 17008 8996 17060
rect 5080 16940 5132 16992
rect 7472 16940 7524 16992
rect 12256 17051 12308 17060
rect 12256 17017 12265 17051
rect 12265 17017 12299 17051
rect 12299 17017 12308 17051
rect 12256 17008 12308 17017
rect 9772 16940 9824 16992
rect 12348 16983 12400 16992
rect 12348 16949 12357 16983
rect 12357 16949 12391 16983
rect 12391 16949 12400 16983
rect 12348 16940 12400 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 4068 16779 4120 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 2136 16600 2188 16652
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 4068 16736 4120 16745
rect 8300 16736 8352 16788
rect 10048 16736 10100 16788
rect 4252 16668 4304 16720
rect 4804 16668 4856 16720
rect 4160 16600 4212 16652
rect 4344 16600 4396 16652
rect 6644 16668 6696 16720
rect 12532 16736 12584 16788
rect 13636 16779 13688 16788
rect 13636 16745 13645 16779
rect 13645 16745 13679 16779
rect 13679 16745 13688 16779
rect 13636 16736 13688 16745
rect 10876 16711 10928 16720
rect 10876 16677 10910 16711
rect 10910 16677 10928 16711
rect 10876 16668 10928 16677
rect 7472 16600 7524 16652
rect 4068 16532 4120 16584
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 9128 16464 9180 16516
rect 9588 16464 9640 16516
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 11704 16396 11756 16448
rect 12164 16532 12216 16584
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1768 16192 1820 16244
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 5080 16235 5132 16244
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 1584 16167 1636 16176
rect 1584 16133 1593 16167
rect 1593 16133 1627 16167
rect 1627 16133 1636 16167
rect 1584 16124 1636 16133
rect 4252 16056 4304 16108
rect 2872 15988 2924 16040
rect 4804 15988 4856 16040
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 12256 16056 12308 16108
rect 2596 15920 2648 15972
rect 3516 15920 3568 15972
rect 5540 15963 5592 15972
rect 5540 15929 5549 15963
rect 5549 15929 5583 15963
rect 5583 15929 5592 15963
rect 10140 15988 10192 16040
rect 5540 15920 5592 15929
rect 2780 15852 2832 15904
rect 3056 15852 3108 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 8760 15895 8812 15904
rect 7104 15852 7156 15861
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 11796 15852 11848 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 2596 15691 2648 15700
rect 2596 15657 2605 15691
rect 2605 15657 2639 15691
rect 2639 15657 2648 15691
rect 2596 15648 2648 15657
rect 1584 15623 1636 15632
rect 1584 15589 1593 15623
rect 1593 15589 1627 15623
rect 1627 15589 1636 15623
rect 1584 15580 1636 15589
rect 4160 15691 4212 15700
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 4804 15648 4856 15700
rect 8760 15648 8812 15700
rect 8944 15648 8996 15700
rect 12348 15648 12400 15700
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 4344 15580 4396 15632
rect 5540 15623 5592 15632
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 3240 15555 3292 15564
rect 2780 15512 2832 15521
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 5540 15589 5549 15623
rect 5549 15589 5583 15623
rect 5583 15589 5592 15623
rect 5540 15580 5592 15589
rect 7380 15580 7432 15632
rect 8760 15512 8812 15564
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 8300 15444 8352 15496
rect 9588 15580 9640 15632
rect 9956 15512 10008 15564
rect 5356 15376 5408 15428
rect 4160 15308 4212 15360
rect 7196 15308 7248 15360
rect 7564 15308 7616 15360
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 12348 15444 12400 15496
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 1768 15104 1820 15156
rect 2964 15104 3016 15156
rect 4344 15104 4396 15156
rect 4896 15104 4948 15156
rect 5448 15104 5500 15156
rect 3516 14968 3568 15020
rect 7104 15104 7156 15156
rect 8668 15104 8720 15156
rect 6920 14968 6972 15020
rect 7104 14968 7156 15020
rect 7380 14968 7432 15020
rect 9956 14968 10008 15020
rect 10416 15011 10468 15020
rect 10416 14977 10425 15011
rect 10425 14977 10459 15011
rect 10459 14977 10468 15011
rect 10416 14968 10468 14977
rect 3148 14900 3200 14952
rect 4160 14900 4212 14952
rect 5816 14943 5868 14952
rect 5816 14909 5834 14943
rect 5834 14909 5868 14943
rect 5816 14900 5868 14909
rect 2688 14832 2740 14884
rect 11152 14832 11204 14884
rect 4804 14764 4856 14816
rect 5264 14764 5316 14816
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 7564 14807 7616 14816
rect 6920 14764 6972 14773
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 9128 14807 9180 14816
rect 7656 14764 7708 14773
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 10140 14807 10192 14816
rect 10140 14773 10149 14807
rect 10149 14773 10183 14807
rect 10183 14773 10192 14807
rect 10784 14807 10836 14816
rect 10140 14764 10192 14773
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2688 14603 2740 14612
rect 2688 14569 2697 14603
rect 2697 14569 2731 14603
rect 2731 14569 2740 14603
rect 2688 14560 2740 14569
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 5816 14560 5868 14612
rect 9128 14560 9180 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 2596 14492 2648 14544
rect 2136 14424 2188 14476
rect 2872 14467 2924 14476
rect 2872 14433 2881 14467
rect 2881 14433 2915 14467
rect 2915 14433 2924 14467
rect 2872 14424 2924 14433
rect 4896 14492 4948 14544
rect 7196 14492 7248 14544
rect 10416 14492 10468 14544
rect 10968 14492 11020 14544
rect 3976 14424 4028 14476
rect 9588 14424 9640 14476
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 5540 14288 5592 14340
rect 6920 14356 6972 14408
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 5632 14220 5684 14272
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2136 14059 2188 14068
rect 2136 14025 2145 14059
rect 2145 14025 2179 14059
rect 2179 14025 2188 14059
rect 2136 14016 2188 14025
rect 3240 14016 3292 14068
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 8576 14059 8628 14068
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 10968 14059 11020 14068
rect 10968 14025 10977 14059
rect 10977 14025 11011 14059
rect 11011 14025 11020 14059
rect 10968 14016 11020 14025
rect 1492 13880 1544 13932
rect 8300 13991 8352 14000
rect 8300 13957 8309 13991
rect 8309 13957 8343 13991
rect 8343 13957 8352 13991
rect 8300 13948 8352 13957
rect 5448 13880 5500 13932
rect 6368 13880 6420 13932
rect 8208 13880 8260 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 3240 13812 3292 13864
rect 4804 13812 4856 13864
rect 5632 13812 5684 13864
rect 1768 13787 1820 13796
rect 1768 13753 1777 13787
rect 1777 13753 1811 13787
rect 1811 13753 1820 13787
rect 1768 13744 1820 13753
rect 5080 13787 5132 13796
rect 5080 13753 5098 13787
rect 5098 13753 5132 13787
rect 8392 13812 8444 13864
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 9864 13855 9916 13864
rect 9864 13821 9887 13855
rect 9887 13821 9916 13855
rect 9864 13812 9916 13821
rect 5080 13744 5132 13753
rect 9220 13744 9272 13796
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 7380 13719 7432 13728
rect 7380 13685 7389 13719
rect 7389 13685 7423 13719
rect 7423 13685 7432 13719
rect 7380 13676 7432 13685
rect 7748 13676 7800 13728
rect 8944 13719 8996 13728
rect 8944 13685 8953 13719
rect 8953 13685 8987 13719
rect 8987 13685 8996 13719
rect 8944 13676 8996 13685
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 1768 13472 1820 13524
rect 2596 13515 2648 13524
rect 2596 13481 2605 13515
rect 2605 13481 2639 13515
rect 2639 13481 2648 13515
rect 2596 13472 2648 13481
rect 2780 13472 2832 13524
rect 3332 13472 3384 13524
rect 4804 13472 4856 13524
rect 4068 13404 4120 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3976 13336 4028 13388
rect 5632 13336 5684 13388
rect 6920 13404 6972 13456
rect 8208 13472 8260 13524
rect 8944 13472 8996 13524
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 10048 13404 10100 13456
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 8392 13336 8444 13388
rect 10232 13336 10284 13388
rect 11244 13379 11296 13388
rect 11244 13345 11253 13379
rect 11253 13345 11287 13379
rect 11287 13345 11296 13379
rect 11244 13336 11296 13345
rect 12164 13336 12216 13388
rect 4344 13268 4396 13320
rect 8576 13311 8628 13320
rect 1584 13243 1636 13252
rect 1584 13209 1593 13243
rect 1593 13209 1627 13243
rect 1627 13209 1636 13243
rect 1584 13200 1636 13209
rect 3240 13200 3292 13252
rect 4160 13200 4212 13252
rect 5080 13200 5132 13252
rect 6368 13200 6420 13252
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 3056 13132 3108 13184
rect 6000 13132 6052 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 2504 12928 2556 12980
rect 2780 12928 2832 12980
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 7380 12928 7432 12980
rect 7748 12971 7800 12980
rect 7748 12937 7757 12971
rect 7757 12937 7791 12971
rect 7791 12937 7800 12971
rect 7748 12928 7800 12937
rect 9036 12928 9088 12980
rect 1860 12792 1912 12844
rect 4252 12860 4304 12912
rect 2596 12792 2648 12844
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 6368 12792 6420 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 8944 12792 8996 12844
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 10232 12835 10284 12844
rect 9220 12792 9272 12801
rect 2320 12656 2372 12708
rect 1400 12631 1452 12640
rect 1400 12597 1409 12631
rect 1409 12597 1443 12631
rect 1443 12597 1452 12631
rect 1400 12588 1452 12597
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 4160 12724 4212 12776
rect 5724 12724 5776 12776
rect 8576 12724 8628 12776
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 4988 12656 5040 12708
rect 6000 12656 6052 12708
rect 5724 12588 5776 12640
rect 6920 12588 6972 12640
rect 7748 12588 7800 12640
rect 8852 12656 8904 12708
rect 19156 12656 19208 12708
rect 9864 12588 9916 12640
rect 10140 12588 10192 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2872 12384 2924 12436
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 5448 12384 5500 12436
rect 2780 12316 2832 12368
rect 3884 12316 3936 12368
rect 5816 12316 5868 12368
rect 6184 12316 6236 12368
rect 8208 12316 8260 12368
rect 10232 12384 10284 12436
rect 1492 12248 1544 12300
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 5632 12248 5684 12300
rect 6092 12291 6144 12300
rect 6092 12257 6110 12291
rect 6110 12257 6144 12291
rect 6092 12248 6144 12257
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 10600 12248 10652 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 1676 12044 1728 12096
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 2872 12044 2924 12096
rect 4896 12180 4948 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6736 12223 6788 12232
rect 6368 12180 6420 12189
rect 6736 12189 6745 12223
rect 6745 12189 6779 12223
rect 6779 12189 6788 12223
rect 6736 12180 6788 12189
rect 3884 12044 3936 12096
rect 8208 12044 8260 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 11704 12044 11756 12096
rect 20812 12044 20864 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2596 11840 2648 11892
rect 3148 11840 3200 11892
rect 4344 11840 4396 11892
rect 7104 11840 7156 11892
rect 9956 11883 10008 11892
rect 9956 11849 9965 11883
rect 9965 11849 9999 11883
rect 9999 11849 10008 11883
rect 9956 11840 10008 11849
rect 11244 11840 11296 11892
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 6552 11772 6604 11824
rect 2780 11704 2832 11756
rect 2872 11704 2924 11756
rect 4988 11704 5040 11756
rect 10600 11747 10652 11756
rect 1584 11636 1636 11688
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 1860 11568 1912 11620
rect 4896 11568 4948 11620
rect 5908 11568 5960 11620
rect 9864 11636 9916 11688
rect 10784 11636 10836 11688
rect 10876 11636 10928 11688
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 2044 11500 2096 11552
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 4344 11543 4396 11552
rect 2320 11500 2372 11509
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 5540 11500 5592 11552
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 6828 11500 6880 11552
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 8484 11500 8536 11552
rect 9772 11500 9824 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2136 11296 2188 11348
rect 2320 11296 2372 11348
rect 2504 11296 2556 11348
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 4620 11296 4672 11348
rect 5632 11296 5684 11348
rect 6092 11296 6144 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 10600 11296 10652 11348
rect 2044 11228 2096 11280
rect 3884 11228 3936 11280
rect 8208 11228 8260 11280
rect 8392 11228 8444 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 3608 11160 3660 11212
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4896 11203 4948 11212
rect 4896 11169 4930 11203
rect 4930 11169 4948 11203
rect 4896 11160 4948 11169
rect 6736 11160 6788 11212
rect 8300 11160 8352 11212
rect 9772 11203 9824 11212
rect 9772 11169 9806 11203
rect 9806 11169 9824 11203
rect 9772 11160 9824 11169
rect 10600 11160 10652 11212
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 4620 11135 4672 11144
rect 3240 11092 3292 11101
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 1492 11024 1544 11076
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 10784 11024 10836 11076
rect 19892 11024 19944 11076
rect 1676 10956 1728 11008
rect 11980 10956 12032 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2780 10752 2832 10804
rect 3240 10752 3292 10804
rect 4804 10752 4856 10804
rect 5080 10752 5132 10804
rect 5448 10752 5500 10804
rect 5724 10752 5776 10804
rect 7472 10752 7524 10804
rect 10416 10752 10468 10804
rect 3240 10548 3292 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4344 10591 4396 10600
rect 4344 10557 4378 10591
rect 4378 10557 4396 10591
rect 4344 10548 4396 10557
rect 5172 10548 5224 10600
rect 5448 10616 5500 10668
rect 9496 10684 9548 10736
rect 8208 10616 8260 10668
rect 9312 10616 9364 10668
rect 9772 10684 9824 10736
rect 10968 10684 11020 10736
rect 10416 10616 10468 10668
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 5632 10548 5684 10600
rect 7012 10591 7064 10600
rect 1952 10523 2004 10532
rect 1952 10489 1986 10523
rect 1986 10489 2004 10523
rect 1952 10480 2004 10489
rect 3332 10412 3384 10464
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 4896 10412 4948 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 9680 10412 9732 10464
rect 9864 10480 9916 10532
rect 11980 10548 12032 10600
rect 12900 10480 12952 10532
rect 13636 10523 13688 10532
rect 13636 10489 13645 10523
rect 13645 10489 13679 10523
rect 13679 10489 13688 10523
rect 13636 10480 13688 10489
rect 10232 10412 10284 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 19432 10412 19484 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 7012 10251 7064 10260
rect 3884 10140 3936 10192
rect 4804 10140 4856 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 2504 10072 2556 10124
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 5172 10072 5224 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 5448 10140 5500 10192
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7104 10208 7156 10260
rect 7380 10208 7432 10260
rect 9036 10208 9088 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 9496 10208 9548 10260
rect 9588 10140 9640 10192
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 6736 10072 6788 10124
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 7748 10072 7800 10124
rect 9220 10072 9272 10124
rect 11060 10140 11112 10192
rect 13544 10140 13596 10192
rect 13268 10072 13320 10124
rect 5448 9936 5500 9988
rect 5540 9936 5592 9988
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 7472 9936 7524 9988
rect 3424 9868 3476 9920
rect 3516 9911 3568 9920
rect 3516 9877 3525 9911
rect 3525 9877 3559 9911
rect 3559 9877 3568 9911
rect 3516 9868 3568 9877
rect 4804 9868 4856 9920
rect 6644 9911 6696 9920
rect 6644 9877 6653 9911
rect 6653 9877 6687 9911
rect 6687 9877 6696 9911
rect 8944 10004 8996 10056
rect 9588 10004 9640 10056
rect 10508 9936 10560 9988
rect 6644 9868 6696 9877
rect 7656 9868 7708 9920
rect 8392 9868 8444 9920
rect 8484 9868 8536 9920
rect 9864 9868 9916 9920
rect 9956 9868 10008 9920
rect 10600 9868 10652 9920
rect 11060 9868 11112 9920
rect 11888 9868 11940 9920
rect 12072 9868 12124 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2596 9664 2648 9716
rect 3148 9664 3200 9716
rect 3240 9664 3292 9716
rect 3976 9639 4028 9648
rect 3976 9605 3985 9639
rect 3985 9605 4019 9639
rect 4019 9605 4028 9639
rect 3976 9596 4028 9605
rect 4988 9596 5040 9648
rect 5448 9664 5500 9716
rect 13544 9707 13596 9716
rect 6000 9596 6052 9648
rect 4712 9571 4764 9580
rect 2596 9392 2648 9444
rect 1952 9324 2004 9376
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 3424 9460 3476 9512
rect 4068 9460 4120 9512
rect 4252 9460 4304 9512
rect 4344 9460 4396 9512
rect 6092 9503 6144 9512
rect 6092 9469 6101 9503
rect 6101 9469 6135 9503
rect 6135 9469 6144 9503
rect 6092 9460 6144 9469
rect 8300 9596 8352 9648
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 10876 9596 10928 9648
rect 13544 9673 13553 9707
rect 13553 9673 13587 9707
rect 13587 9673 13596 9707
rect 13544 9664 13596 9673
rect 15844 9664 15896 9716
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 7656 9460 7708 9512
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 13084 9460 13136 9512
rect 3976 9392 4028 9444
rect 9312 9392 9364 9444
rect 9588 9392 9640 9444
rect 9956 9392 10008 9444
rect 10508 9392 10560 9444
rect 11244 9392 11296 9444
rect 14556 9392 14608 9444
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 4804 9324 4856 9376
rect 5540 9324 5592 9376
rect 6000 9324 6052 9376
rect 10968 9324 11020 9376
rect 11428 9324 11480 9376
rect 12992 9324 13044 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2688 9120 2740 9172
rect 3516 9120 3568 9172
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 4804 9163 4856 9172
rect 4804 9129 4813 9163
rect 4813 9129 4847 9163
rect 4847 9129 4856 9163
rect 4804 9120 4856 9129
rect 6276 9120 6328 9172
rect 6000 9052 6052 9104
rect 6092 9052 6144 9104
rect 7380 9120 7432 9172
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 9680 9163 9732 9172
rect 8392 9120 8444 9129
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 11704 9120 11756 9172
rect 12992 9120 13044 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 3516 8984 3568 9036
rect 4344 8984 4396 9036
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 2872 8916 2924 8968
rect 3148 8916 3200 8968
rect 4988 8916 5040 8968
rect 5264 8848 5316 8900
rect 2044 8780 2096 8832
rect 2688 8780 2740 8832
rect 4804 8780 4856 8832
rect 5724 8780 5776 8832
rect 6184 8984 6236 9036
rect 9404 9052 9456 9104
rect 12164 9052 12216 9104
rect 9128 8984 9180 9036
rect 10784 8984 10836 9036
rect 15292 8984 15344 9036
rect 7472 8916 7524 8968
rect 8300 8916 8352 8968
rect 9312 8916 9364 8968
rect 10508 8916 10560 8968
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 12072 8916 12124 8968
rect 13268 8916 13320 8968
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7380 8780 7432 8832
rect 11428 8848 11480 8900
rect 8668 8780 8720 8832
rect 9220 8780 9272 8832
rect 13544 8780 13596 8832
rect 14096 8780 14148 8832
rect 15568 8780 15620 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3516 8576 3568 8628
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 1768 8236 1820 8288
rect 2596 8372 2648 8424
rect 5816 8508 5868 8560
rect 8760 8576 8812 8628
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 9496 8576 9548 8628
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 11888 8508 11940 8560
rect 13360 8508 13412 8560
rect 18696 8508 18748 8560
rect 6460 8440 6512 8492
rect 6920 8440 6972 8492
rect 8576 8440 8628 8492
rect 3700 8372 3752 8424
rect 4252 8372 4304 8424
rect 2228 8347 2280 8356
rect 2228 8313 2262 8347
rect 2262 8313 2280 8347
rect 2228 8304 2280 8313
rect 5724 8372 5776 8424
rect 6368 8372 6420 8424
rect 5448 8304 5500 8356
rect 6000 8347 6052 8356
rect 6000 8313 6009 8347
rect 6009 8313 6043 8347
rect 6043 8313 6052 8347
rect 6000 8304 6052 8313
rect 6092 8304 6144 8356
rect 7380 8304 7432 8356
rect 7656 8372 7708 8424
rect 5264 8236 5316 8288
rect 6920 8236 6972 8288
rect 7196 8236 7248 8288
rect 7748 8304 7800 8356
rect 8208 8304 8260 8356
rect 9220 8372 9272 8424
rect 9404 8440 9456 8492
rect 10416 8440 10468 8492
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 10876 8372 10928 8424
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 12900 8415 12952 8424
rect 10508 8236 10560 8288
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 13544 8372 13596 8424
rect 12440 8304 12492 8356
rect 14740 8304 14792 8356
rect 11704 8236 11756 8288
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 15752 8236 15804 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1400 8075 1452 8084
rect 1400 8041 1409 8075
rect 1409 8041 1443 8075
rect 1443 8041 1452 8075
rect 1400 8032 1452 8041
rect 2872 8032 2924 8084
rect 4160 8032 4212 8084
rect 4804 8032 4856 8084
rect 1676 7896 1728 7948
rect 2596 7896 2648 7948
rect 5632 8032 5684 8084
rect 11980 8032 12032 8084
rect 4896 7896 4948 7948
rect 2780 7828 2832 7880
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 4804 7871 4856 7880
rect 3332 7828 3384 7837
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5816 7964 5868 8016
rect 6644 7896 6696 7948
rect 7104 7896 7156 7948
rect 7932 7964 7984 8016
rect 14096 8032 14148 8084
rect 15384 8032 15436 8084
rect 5540 7760 5592 7812
rect 6184 7828 6236 7880
rect 7196 7828 7248 7880
rect 8944 7896 8996 7948
rect 9496 7896 9548 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 11980 7896 12032 7948
rect 9404 7871 9456 7880
rect 6644 7760 6696 7812
rect 7380 7760 7432 7812
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 8300 7803 8352 7812
rect 8300 7769 8309 7803
rect 8309 7769 8343 7803
rect 8343 7769 8352 7803
rect 8300 7760 8352 7769
rect 14924 8007 14976 8016
rect 14924 7973 14933 8007
rect 14933 7973 14967 8007
rect 14967 7973 14976 8007
rect 14924 7964 14976 7973
rect 2228 7692 2280 7744
rect 3332 7692 3384 7744
rect 3792 7692 3844 7744
rect 4068 7692 4120 7744
rect 5632 7692 5684 7744
rect 6552 7692 6604 7744
rect 11244 7692 11296 7744
rect 13268 7692 13320 7744
rect 15568 7896 15620 7948
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 16580 7896 16632 7948
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 17684 7828 17736 7880
rect 17868 7692 17920 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3332 7488 3384 7540
rect 4804 7488 4856 7540
rect 11980 7488 12032 7540
rect 6828 7420 6880 7472
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 7196 7395 7248 7404
rect 5724 7352 5776 7361
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 11888 7420 11940 7472
rect 12440 7488 12492 7540
rect 11704 7352 11756 7404
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 1492 7216 1544 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 3976 7284 4028 7336
rect 4344 7327 4396 7336
rect 4344 7293 4353 7327
rect 4353 7293 4387 7327
rect 4387 7293 4396 7327
rect 4344 7284 4396 7293
rect 4436 7284 4488 7336
rect 6920 7216 6972 7268
rect 7748 7284 7800 7336
rect 7932 7327 7984 7336
rect 7932 7293 7966 7327
rect 7966 7293 7984 7327
rect 7932 7284 7984 7293
rect 9220 7216 9272 7268
rect 9404 7284 9456 7336
rect 12072 7284 12124 7336
rect 13268 7352 13320 7404
rect 10508 7216 10560 7268
rect 11888 7216 11940 7268
rect 13544 7216 13596 7268
rect 1400 7148 1452 7157
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 4896 7148 4948 7200
rect 9588 7148 9640 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 10784 7148 10836 7200
rect 17684 7284 17736 7336
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2320 6944 2372 6996
rect 4528 6944 4580 6996
rect 14188 6944 14240 6996
rect 3056 6876 3108 6928
rect 2780 6808 2832 6860
rect 5356 6876 5408 6928
rect 6184 6808 6236 6860
rect 6276 6808 6328 6860
rect 6828 6808 6880 6860
rect 8208 6808 8260 6860
rect 9680 6808 9732 6860
rect 2964 6740 3016 6792
rect 2136 6604 2188 6656
rect 4160 6740 4212 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 6920 6783 6972 6792
rect 3700 6672 3752 6724
rect 5172 6604 5224 6656
rect 5264 6604 5316 6656
rect 5632 6672 5684 6724
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 10324 6808 10376 6860
rect 11244 6876 11296 6928
rect 10416 6740 10468 6792
rect 10508 6740 10560 6792
rect 8484 6672 8536 6724
rect 9680 6672 9732 6724
rect 10048 6672 10100 6724
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 6736 6604 6788 6656
rect 8760 6604 8812 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12256 6647 12308 6656
rect 12256 6613 12265 6647
rect 12265 6613 12299 6647
rect 12299 6613 12308 6647
rect 12256 6604 12308 6613
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 14740 6876 14792 6928
rect 13360 6808 13412 6860
rect 14924 6851 14976 6860
rect 14924 6817 14933 6851
rect 14933 6817 14967 6851
rect 14967 6817 14976 6851
rect 14924 6808 14976 6817
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 16948 6808 17000 6860
rect 17224 6851 17276 6860
rect 17224 6817 17242 6851
rect 17242 6817 17276 6851
rect 17224 6808 17276 6817
rect 17684 6740 17736 6792
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 14372 6604 14424 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16580 6604 16632 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 1492 6400 1544 6452
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 3700 6332 3752 6384
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 6184 6332 6236 6384
rect 8392 6400 8444 6452
rect 8668 6400 8720 6452
rect 13360 6400 13412 6452
rect 13544 6443 13596 6452
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 15016 6400 15068 6452
rect 18604 6400 18656 6452
rect 10508 6332 10560 6384
rect 4160 6264 4212 6273
rect 6460 6264 6512 6316
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10784 6264 10836 6316
rect 11060 6332 11112 6384
rect 11244 6332 11296 6384
rect 2872 6196 2924 6248
rect 3608 6196 3660 6248
rect 4804 6196 4856 6248
rect 6920 6196 6972 6248
rect 9128 6196 9180 6248
rect 9220 6196 9272 6248
rect 5724 6171 5776 6180
rect 5724 6137 5742 6171
rect 5742 6137 5776 6171
rect 5724 6128 5776 6137
rect 9404 6128 9456 6180
rect 10416 6128 10468 6180
rect 3240 6060 3292 6112
rect 6276 6060 6328 6112
rect 6552 6060 6604 6112
rect 7104 6060 7156 6112
rect 8300 6060 8352 6112
rect 9036 6060 9088 6112
rect 11980 6264 12032 6316
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 11060 6060 11112 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 14924 6264 14976 6316
rect 16580 6264 16632 6316
rect 17132 6264 17184 6316
rect 13268 6196 13320 6248
rect 17592 6239 17644 6248
rect 17592 6205 17601 6239
rect 17601 6205 17635 6239
rect 17635 6205 17644 6239
rect 17592 6196 17644 6205
rect 12256 6128 12308 6180
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 13912 6060 13964 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16396 6060 16448 6112
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 2412 5856 2464 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 4988 5856 5040 5908
rect 6184 5856 6236 5908
rect 6368 5856 6420 5908
rect 6828 5856 6880 5908
rect 6920 5856 6972 5908
rect 4160 5788 4212 5840
rect 1492 5652 1544 5704
rect 3700 5720 3752 5772
rect 3516 5652 3568 5704
rect 3884 5652 3936 5704
rect 4896 5788 4948 5840
rect 3792 5584 3844 5636
rect 5632 5720 5684 5772
rect 6092 5720 6144 5772
rect 7104 5720 7156 5772
rect 5448 5652 5500 5704
rect 7472 5856 7524 5908
rect 7748 5788 7800 5840
rect 9680 5831 9732 5840
rect 9680 5797 9714 5831
rect 9714 5797 9732 5831
rect 9680 5788 9732 5797
rect 10692 5788 10744 5840
rect 10876 5856 10928 5908
rect 13360 5856 13412 5908
rect 11060 5788 11112 5840
rect 12256 5788 12308 5840
rect 13912 5856 13964 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 17500 5856 17552 5908
rect 7472 5720 7524 5772
rect 8208 5720 8260 5772
rect 9128 5720 9180 5772
rect 9956 5720 10008 5772
rect 10416 5720 10468 5772
rect 11244 5720 11296 5772
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8392 5652 8444 5704
rect 11060 5695 11112 5704
rect 1584 5516 1636 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 8208 5516 8260 5568
rect 8392 5559 8444 5568
rect 8392 5525 8401 5559
rect 8401 5525 8435 5559
rect 8435 5525 8444 5559
rect 8392 5516 8444 5525
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11888 5720 11940 5772
rect 13268 5720 13320 5772
rect 14556 5763 14608 5772
rect 11980 5652 12032 5704
rect 12624 5652 12676 5704
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 15844 5720 15896 5772
rect 21364 5763 21416 5772
rect 21364 5729 21373 5763
rect 21373 5729 21407 5763
rect 21407 5729 21416 5763
rect 21364 5720 21416 5729
rect 16672 5652 16724 5704
rect 17132 5652 17184 5704
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 12900 5516 12952 5568
rect 14556 5516 14608 5568
rect 15752 5559 15804 5568
rect 15752 5525 15761 5559
rect 15761 5525 15795 5559
rect 15795 5525 15804 5559
rect 15752 5516 15804 5525
rect 21180 5559 21232 5568
rect 21180 5525 21189 5559
rect 21189 5525 21223 5559
rect 21223 5525 21232 5559
rect 21180 5516 21232 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3976 5312 4028 5364
rect 5632 5312 5684 5364
rect 5908 5355 5960 5364
rect 5908 5321 5917 5355
rect 5917 5321 5951 5355
rect 5951 5321 5960 5355
rect 5908 5312 5960 5321
rect 7932 5312 7984 5364
rect 8300 5312 8352 5364
rect 11244 5312 11296 5364
rect 11796 5312 11848 5364
rect 12348 5355 12400 5364
rect 12348 5321 12357 5355
rect 12357 5321 12391 5355
rect 12391 5321 12400 5355
rect 12348 5312 12400 5321
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 2320 5244 2372 5296
rect 1952 5176 2004 5228
rect 3332 5176 3384 5228
rect 7196 5244 7248 5296
rect 4068 5176 4120 5228
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 3700 5108 3752 5160
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 4344 5108 4396 5117
rect 4896 5108 4948 5160
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 5448 5108 5500 5160
rect 6000 5108 6052 5160
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 8392 5176 8444 5228
rect 9680 5176 9732 5228
rect 10784 5176 10836 5228
rect 12072 5244 12124 5296
rect 17408 5244 17460 5296
rect 15660 5219 15712 5228
rect 10048 5108 10100 5160
rect 11060 5108 11112 5160
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 12624 5108 12676 5160
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 14648 5108 14700 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 17684 5108 17736 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 2136 5040 2188 5092
rect 4252 5040 4304 5092
rect 8484 5040 8536 5092
rect 9864 5040 9916 5092
rect 10324 5040 10376 5092
rect 17224 5040 17276 5092
rect 2412 4972 2464 5024
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 4712 4972 4764 5024
rect 5356 4972 5408 5024
rect 5632 4972 5684 5024
rect 7656 4972 7708 5024
rect 9312 4972 9364 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 14740 4972 14792 5024
rect 15384 4972 15436 5024
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1952 4768 2004 4820
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 5540 4768 5592 4820
rect 5632 4768 5684 4820
rect 2688 4700 2740 4752
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 4068 4675 4120 4684
rect 2780 4632 2832 4641
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4712 4675 4764 4684
rect 4712 4641 4721 4675
rect 4721 4641 4755 4675
rect 4755 4641 4764 4675
rect 4712 4632 4764 4641
rect 5908 4700 5960 4752
rect 6092 4700 6144 4752
rect 7748 4768 7800 4820
rect 8852 4768 8904 4820
rect 9772 4768 9824 4820
rect 10140 4768 10192 4820
rect 11152 4768 11204 4820
rect 5632 4632 5684 4684
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 10324 4700 10376 4752
rect 10784 4743 10836 4752
rect 10784 4709 10818 4743
rect 10818 4709 10836 4743
rect 10784 4700 10836 4709
rect 13728 4768 13780 4820
rect 14096 4768 14148 4820
rect 17224 4811 17276 4820
rect 2228 4496 2280 4548
rect 5540 4496 5592 4548
rect 3056 4428 3108 4480
rect 3884 4428 3936 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4804 4428 4856 4480
rect 7104 4564 7156 4616
rect 7288 4564 7340 4616
rect 8392 4632 8444 4684
rect 8760 4675 8812 4684
rect 8760 4641 8769 4675
rect 8769 4641 8803 4675
rect 8803 4641 8812 4675
rect 8760 4632 8812 4641
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 10416 4632 10468 4684
rect 13084 4700 13136 4752
rect 11060 4632 11112 4684
rect 11980 4632 12032 4684
rect 12256 4632 12308 4684
rect 13176 4632 13228 4684
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 15660 4700 15712 4752
rect 16396 4700 16448 4752
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 21180 4700 21232 4752
rect 13268 4632 13320 4641
rect 14372 4632 14424 4684
rect 14740 4632 14792 4684
rect 15568 4632 15620 4684
rect 18512 4632 18564 4684
rect 9588 4564 9640 4616
rect 9956 4564 10008 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 13360 4564 13412 4616
rect 6276 4496 6328 4548
rect 9312 4496 9364 4548
rect 9772 4496 9824 4548
rect 5816 4428 5868 4480
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 9404 4428 9456 4480
rect 11796 4428 11848 4480
rect 12164 4496 12216 4548
rect 13176 4496 13228 4548
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 15476 4496 15528 4548
rect 12532 4428 12584 4480
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16212 4428 16264 4480
rect 18052 4471 18104 4480
rect 18052 4437 18061 4471
rect 18061 4437 18095 4471
rect 18095 4437 18104 4471
rect 18052 4428 18104 4437
rect 18144 4428 18196 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2872 4224 2924 4276
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 1860 4088 1912 4140
rect 4896 4224 4948 4276
rect 5356 4224 5408 4276
rect 7012 4224 7064 4276
rect 7288 4224 7340 4276
rect 1768 4020 1820 4072
rect 2228 4063 2280 4072
rect 2228 4029 2262 4063
rect 2262 4029 2280 4063
rect 2228 4020 2280 4029
rect 2504 4020 2556 4072
rect 4436 4020 4488 4072
rect 3332 3884 3384 3936
rect 5540 3884 5592 3936
rect 5724 4088 5776 4140
rect 6000 4088 6052 4140
rect 6460 4088 6512 4140
rect 11060 4224 11112 4276
rect 9772 4156 9824 4208
rect 14096 4224 14148 4276
rect 16396 4267 16448 4276
rect 16396 4233 16405 4267
rect 16405 4233 16439 4267
rect 16439 4233 16448 4267
rect 16396 4224 16448 4233
rect 17224 4156 17276 4208
rect 7656 4020 7708 4072
rect 9036 4020 9088 4072
rect 9588 4020 9640 4072
rect 9772 4020 9824 4072
rect 11796 4088 11848 4140
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 6920 3995 6972 4004
rect 6920 3961 6954 3995
rect 6954 3961 6972 3995
rect 6920 3952 6972 3961
rect 10140 3952 10192 4004
rect 10600 3952 10652 4004
rect 11520 3952 11572 4004
rect 14004 4088 14056 4140
rect 19248 4156 19300 4208
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 15660 4020 15712 4072
rect 17500 4063 17552 4072
rect 17500 4029 17509 4063
rect 17509 4029 17543 4063
rect 17543 4029 17552 4063
rect 17500 4020 17552 4029
rect 17592 4020 17644 4072
rect 18604 4063 18656 4072
rect 18604 4029 18613 4063
rect 18613 4029 18647 4063
rect 18647 4029 18656 4063
rect 18604 4020 18656 4029
rect 21824 4088 21876 4140
rect 20536 4020 20588 4072
rect 11704 3952 11756 4004
rect 12624 3952 12676 4004
rect 13912 3995 13964 4004
rect 13912 3961 13921 3995
rect 13921 3961 13955 3995
rect 13955 3961 13964 3995
rect 13912 3952 13964 3961
rect 15936 3952 15988 4004
rect 6736 3884 6788 3936
rect 7104 3884 7156 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8300 3884 8352 3893
rect 8484 3884 8536 3936
rect 12808 3884 12860 3936
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 16028 3884 16080 3936
rect 17960 3884 18012 3936
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 19064 3927 19116 3936
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 20720 3952 20772 4004
rect 20904 3995 20956 4004
rect 20904 3961 20913 3995
rect 20913 3961 20947 3995
rect 20947 3961 20956 3995
rect 20904 3952 20956 3961
rect 21364 3884 21416 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2228 3680 2280 3732
rect 1032 3612 1084 3664
rect 4068 3680 4120 3732
rect 4160 3680 4212 3732
rect 5172 3680 5224 3732
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 6092 3680 6144 3732
rect 2872 3612 2924 3664
rect 3148 3612 3200 3664
rect 1492 3544 1544 3596
rect 3332 3587 3384 3596
rect 2964 3476 3016 3528
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 3516 3544 3568 3596
rect 3884 3544 3936 3596
rect 4436 3544 4488 3596
rect 4344 3476 4396 3528
rect 5264 3612 5316 3664
rect 7012 3680 7064 3732
rect 7380 3680 7432 3732
rect 8208 3680 8260 3732
rect 9680 3680 9732 3732
rect 10232 3680 10284 3732
rect 10784 3680 10836 3732
rect 12072 3680 12124 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 9036 3612 9088 3664
rect 6000 3544 6052 3596
rect 572 3408 624 3460
rect 3792 3408 3844 3460
rect 3056 3340 3108 3392
rect 3240 3383 3292 3392
rect 3240 3349 3249 3383
rect 3249 3349 3283 3383
rect 3283 3349 3292 3383
rect 3240 3340 3292 3349
rect 9772 3544 9824 3596
rect 10048 3544 10100 3596
rect 11612 3612 11664 3664
rect 13268 3612 13320 3664
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 8576 3476 8628 3528
rect 7380 3408 7432 3460
rect 9680 3476 9732 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 12072 3544 12124 3596
rect 13360 3544 13412 3596
rect 15660 3680 15712 3732
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 15568 3612 15620 3664
rect 20628 3680 20680 3732
rect 15384 3544 15436 3596
rect 19340 3612 19392 3664
rect 20812 3655 20864 3664
rect 20812 3621 20821 3655
rect 20821 3621 20855 3655
rect 20855 3621 20864 3655
rect 20812 3612 20864 3621
rect 17868 3544 17920 3596
rect 18696 3544 18748 3596
rect 19248 3587 19300 3596
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 21364 3587 21416 3596
rect 21364 3553 21373 3587
rect 21373 3553 21407 3587
rect 21407 3553 21416 3587
rect 21364 3544 21416 3553
rect 12348 3519 12400 3528
rect 6460 3340 6512 3392
rect 6920 3340 6972 3392
rect 7932 3340 7984 3392
rect 9864 3340 9916 3392
rect 9956 3340 10008 3392
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 16764 3519 16816 3528
rect 11520 3408 11572 3460
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 16120 3408 16172 3460
rect 19248 3408 19300 3460
rect 20076 3451 20128 3460
rect 20076 3417 20085 3451
rect 20085 3417 20119 3451
rect 20119 3417 20128 3451
rect 20076 3408 20128 3417
rect 20536 3408 20588 3460
rect 11796 3340 11848 3392
rect 13544 3340 13596 3392
rect 17316 3340 17368 3392
rect 18144 3340 18196 3392
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 21364 3340 21416 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 1676 3136 1728 3188
rect 2780 3136 2832 3188
rect 4804 3136 4856 3188
rect 2872 3000 2924 3052
rect 3240 3000 3292 3052
rect 3424 2932 3476 2984
rect 6460 3068 6512 3120
rect 6644 3068 6696 3120
rect 7472 3068 7524 3120
rect 3976 2932 4028 2984
rect 5448 3000 5500 3052
rect 5908 3000 5960 3052
rect 6000 3000 6052 3052
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4528 2932 4580 2941
rect 6736 2932 6788 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 5540 2864 5592 2916
rect 7012 2907 7064 2916
rect 204 2796 256 2848
rect 1584 2796 1636 2848
rect 3240 2796 3292 2848
rect 3332 2796 3384 2848
rect 3700 2796 3752 2848
rect 5908 2796 5960 2848
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 9772 3136 9824 3188
rect 14648 3136 14700 3188
rect 17592 3136 17644 3188
rect 11060 3068 11112 3120
rect 11336 3068 11388 3120
rect 13176 3068 13228 3120
rect 13636 3068 13688 3120
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 10600 3000 10652 3052
rect 8484 2932 8536 2984
rect 10692 2932 10744 2984
rect 10876 2932 10928 2984
rect 8208 2864 8260 2916
rect 9680 2864 9732 2916
rect 10232 2864 10284 2916
rect 13268 3000 13320 3052
rect 14280 3000 14332 3052
rect 11796 2932 11848 2984
rect 12348 2932 12400 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 13728 2932 13780 2984
rect 14740 2932 14792 2984
rect 15936 3000 15988 3052
rect 16948 3000 17000 3052
rect 16764 2932 16816 2984
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 17960 2932 18012 2984
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 19432 2932 19484 2984
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 20720 2932 20772 2984
rect 22744 2932 22796 2984
rect 8300 2796 8352 2848
rect 8484 2796 8536 2848
rect 10048 2796 10100 2848
rect 10140 2796 10192 2848
rect 10692 2839 10744 2848
rect 10692 2805 10701 2839
rect 10701 2805 10735 2839
rect 10735 2805 10744 2839
rect 10692 2796 10744 2805
rect 10876 2796 10928 2848
rect 11888 2796 11940 2848
rect 12716 2796 12768 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 13820 2796 13872 2848
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 15200 2864 15252 2916
rect 15660 2864 15712 2916
rect 16212 2796 16264 2848
rect 16488 2864 16540 2916
rect 19156 2907 19208 2916
rect 19156 2873 19165 2907
rect 19165 2873 19199 2907
rect 19199 2873 19208 2907
rect 19156 2864 19208 2873
rect 19616 2864 19668 2916
rect 17960 2796 18012 2848
rect 18604 2839 18656 2848
rect 18604 2805 18613 2839
rect 18613 2805 18647 2839
rect 18647 2805 18656 2839
rect 18604 2796 18656 2805
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 4068 2592 4120 2644
rect 5080 2592 5132 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 7196 2592 7248 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 9864 2635 9916 2644
rect 1584 2524 1636 2576
rect 3884 2524 3936 2576
rect 3976 2524 4028 2576
rect 2964 2456 3016 2508
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4068 2456 4120 2508
rect 6092 2524 6144 2576
rect 7380 2524 7432 2576
rect 9864 2601 9873 2635
rect 9873 2601 9907 2635
rect 9907 2601 9916 2635
rect 9864 2592 9916 2601
rect 10140 2592 10192 2644
rect 11152 2592 11204 2644
rect 11060 2524 11112 2576
rect 12716 2567 12768 2576
rect 4896 2456 4948 2508
rect 6184 2456 6236 2508
rect 6920 2388 6972 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 2596 2252 2648 2304
rect 6184 2295 6236 2304
rect 6184 2261 6193 2295
rect 6193 2261 6227 2295
rect 6227 2261 6236 2295
rect 6184 2252 6236 2261
rect 6368 2320 6420 2372
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9680 2456 9732 2508
rect 11244 2456 11296 2508
rect 12716 2533 12725 2567
rect 12725 2533 12759 2567
rect 12759 2533 12768 2567
rect 12716 2524 12768 2533
rect 13820 2567 13872 2576
rect 13820 2533 13829 2567
rect 13829 2533 13863 2567
rect 13863 2533 13872 2567
rect 13820 2524 13872 2533
rect 14188 2524 14240 2576
rect 15476 2567 15528 2576
rect 15476 2533 15485 2567
rect 15485 2533 15519 2567
rect 15519 2533 15528 2567
rect 15476 2524 15528 2533
rect 16028 2567 16080 2576
rect 16028 2533 16037 2567
rect 16037 2533 16071 2567
rect 16071 2533 16080 2567
rect 16028 2524 16080 2533
rect 17960 2524 18012 2576
rect 18144 2567 18196 2576
rect 18144 2533 18153 2567
rect 18153 2533 18187 2567
rect 18187 2533 18196 2567
rect 18144 2524 18196 2533
rect 18604 2524 18656 2576
rect 19248 2567 19300 2576
rect 19248 2533 19257 2567
rect 19257 2533 19291 2567
rect 19291 2533 19300 2567
rect 19248 2524 19300 2533
rect 18512 2456 18564 2508
rect 20352 2592 20404 2644
rect 20628 2567 20680 2576
rect 20628 2533 20637 2567
rect 20637 2533 20671 2567
rect 20671 2533 20680 2567
rect 20628 2524 20680 2533
rect 21364 2456 21416 2508
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 12532 2363 12584 2372
rect 7012 2252 7064 2304
rect 7564 2252 7616 2304
rect 12532 2329 12541 2363
rect 12541 2329 12575 2363
rect 12575 2329 12584 2363
rect 12532 2320 12584 2329
rect 12992 2320 13044 2372
rect 13452 2320 13504 2372
rect 13912 2320 13964 2372
rect 14832 2320 14884 2372
rect 16948 2320 17000 2372
rect 17500 2320 17552 2372
rect 18604 2388 18656 2440
rect 18696 2320 18748 2372
rect 22284 2320 22336 2372
rect 13728 2252 13780 2304
rect 14280 2252 14332 2304
rect 17868 2252 17920 2304
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 6184 2048 6236 2100
rect 9956 2048 10008 2100
rect 4068 1980 4120 2032
rect 4896 1912 4948 1964
rect 16672 2048 16724 2100
rect 21180 2048 21232 2100
rect 18052 1980 18104 2032
rect 10324 1912 10376 1964
rect 12256 1912 12308 1964
rect 2964 1844 3016 1896
rect 16580 1912 16632 1964
rect 19064 1844 19116 1896
rect 4160 1776 4212 1828
rect 8392 1776 8444 1828
rect 4988 1708 5040 1760
rect 6552 1708 6604 1760
rect 2780 1368 2832 1420
rect 3792 1368 3844 1420
<< metal2 >>
rect 2870 22672 2926 22681
rect 2870 22607 2926 22616
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 2226 20768 2282 20777
rect 2226 20703 2282 20712
rect 2134 20360 2190 20369
rect 2134 20295 2136 20304
rect 2188 20295 2190 20304
rect 2136 20266 2188 20272
rect 2240 20058 2268 20703
rect 2792 20534 2820 21247
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2884 20482 2912 22607
rect 4066 22264 4122 22273
rect 4066 22199 4122 22208
rect 3238 21720 3294 21729
rect 3238 21655 3294 21664
rect 3252 20534 3280 21655
rect 4080 20534 4108 22199
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 3240 20528 3292 20534
rect 2884 20466 3004 20482
rect 3240 20470 3292 20476
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 2872 20460 3004 20466
rect 2924 20454 3004 20460
rect 2872 20402 2924 20408
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 1584 19848 1636 19854
rect 1582 19816 1584 19825
rect 1636 19816 1638 19825
rect 1582 19751 1638 19760
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1596 19310 1624 19343
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1780 18970 1808 19178
rect 2240 18970 2268 19858
rect 2332 19514 2360 20266
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 19514 2636 19858
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 1584 18896 1636 18902
rect 1582 18864 1584 18873
rect 1636 18864 1638 18873
rect 1582 18799 1638 18808
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1780 18358 1808 18770
rect 2226 18456 2282 18465
rect 2226 18391 2228 18400
rect 2280 18391 2282 18400
rect 2228 18362 2280 18368
rect 1768 18352 1820 18358
rect 1768 18294 1820 18300
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 1676 18080 1728 18086
rect 1674 18048 1676 18057
rect 1728 18048 1730 18057
rect 1674 17983 1730 17992
rect 1780 17882 1808 18090
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1676 17536 1728 17542
rect 1674 17504 1676 17513
rect 1728 17504 1730 17513
rect 1674 17439 1730 17448
rect 1780 17338 1808 17682
rect 2332 17338 2360 18090
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2516 17270 2544 17682
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2320 17128 2372 17134
rect 1582 17096 1638 17105
rect 2320 17070 2372 17076
rect 1582 17031 1584 17040
rect 1636 17031 1638 17040
rect 1768 17060 1820 17066
rect 1584 17002 1636 17008
rect 1768 17002 1820 17008
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16561 1624 16594
rect 1582 16552 1638 16561
rect 1582 16487 1638 16496
rect 1780 16250 1808 17002
rect 2332 16794 2360 17070
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1584 16176 1636 16182
rect 1582 16144 1584 16153
rect 1636 16144 1638 16153
rect 1582 16079 1638 16088
rect 2148 15706 2176 16594
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 2608 15706 2636 15914
rect 2792 15910 2820 20198
rect 2884 20058 2912 20266
rect 2976 20058 3004 20454
rect 3424 20324 3476 20330
rect 3424 20266 3476 20272
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3436 19514 3464 20266
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 2976 18970 3004 19246
rect 3620 18970 3648 19246
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2884 17882 2912 18158
rect 3068 17882 3096 18702
rect 3160 18426 3188 18770
rect 4080 18698 4108 19858
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 6840 17814 6868 18702
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17882 7328 18022
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 17134 3740 17478
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16046 2912 16934
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 1584 15632 1636 15638
rect 1582 15600 1584 15609
rect 1636 15600 1638 15609
rect 1582 15535 1638 15544
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 1674 15192 1730 15201
rect 1780 15162 1808 15506
rect 1674 15127 1676 15136
rect 1728 15127 1730 15136
rect 1768 15156 1820 15162
rect 1676 15098 1728 15104
rect 1768 15098 1820 15104
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2226 14648 2282 14657
rect 2700 14618 2728 14826
rect 2226 14583 2228 14592
rect 2280 14583 2282 14592
rect 2688 14612 2740 14618
rect 2228 14554 2280 14560
rect 2688 14554 2740 14560
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 1676 14272 1728 14278
rect 1674 14240 1676 14249
rect 1728 14240 1730 14249
rect 1674 14175 1730 14184
rect 2148 14074 2176 14418
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 11218 1440 12582
rect 1504 12306 1532 13874
rect 1584 13864 1636 13870
rect 1582 13832 1584 13841
rect 1636 13832 1638 13841
rect 1582 13767 1638 13776
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1780 13530 1808 13738
rect 2608 13530 2636 14486
rect 2792 13530 2820 15506
rect 2976 15162 3004 17070
rect 4816 17066 4844 17614
rect 5552 17338 5580 17682
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4080 16794 4108 17002
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4080 16590 4108 16730
rect 4816 16726 4844 17002
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 1582 13288 1638 13297
rect 1582 13223 1584 13232
rect 1636 13223 1638 13232
rect 1584 13194 1636 13200
rect 1780 12986 1808 13330
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 11393 1532 12242
rect 1872 12102 1900 12786
rect 2332 12714 2360 13330
rect 2424 13110 2636 13138
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10441 1440 11154
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1504 10282 1532 11018
rect 1596 10985 1624 11630
rect 1688 11014 1716 12038
rect 1872 11626 1900 12038
rect 2226 11656 2282 11665
rect 1860 11620 1912 11626
rect 2226 11591 2282 11600
rect 1860 11562 1912 11568
rect 2240 11558 2268 11591
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2056 11286 2084 11494
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 1676 11008 1728 11014
rect 1582 10976 1638 10985
rect 1676 10950 1728 10956
rect 1582 10911 1638 10920
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1412 10254 1532 10282
rect 1412 10130 1440 10254
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1412 9489 1440 10066
rect 1872 10033 1900 10066
rect 1858 10024 1914 10033
rect 1858 9959 1914 9968
rect 1398 9480 1454 9489
rect 1398 9415 1454 9424
rect 1964 9382 1992 10474
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1398 9072 1454 9081
rect 1398 9007 1400 9016
rect 1452 9007 1454 9016
rect 1400 8978 1452 8984
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1398 8664 1454 8673
rect 1398 8599 1454 8608
rect 1412 8430 1440 8599
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8090 1440 8366
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 5817 1440 7142
rect 1504 6458 1532 7210
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 1504 5710 1532 6394
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1032 3664 1084 3670
rect 1032 3606 1084 3612
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 584 800 612 3402
rect 1044 800 1072 3606
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1504 800 1532 3538
rect 1596 2854 1624 5510
rect 1688 3194 1716 7890
rect 1780 7342 1808 8230
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 4078 1808 7278
rect 1858 6896 1914 6905
rect 1858 6831 1914 6840
rect 1872 4146 1900 6831
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4826 1992 5170
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1950 4584 2006 4593
rect 1950 4519 2006 4528
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2582 1624 2790
rect 1872 2774 1900 4082
rect 1688 2746 1900 2774
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 1688 1601 1716 2746
rect 1674 1592 1730 1601
rect 1674 1527 1730 1536
rect 1964 800 1992 4519
rect 2056 4049 2084 8774
rect 2148 7993 2176 11290
rect 2240 8922 2268 11494
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2240 8894 2360 8922
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2134 7984 2190 7993
rect 2134 7919 2190 7928
rect 2240 7750 2268 8298
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2332 7002 2360 8894
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 5914 2176 6598
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2332 5302 2360 6938
rect 2424 5914 2452 13110
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2516 11354 2544 12922
rect 2608 12850 2636 13110
rect 2792 12986 2820 13330
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 11898 2636 12582
rect 2884 12442 2912 14418
rect 3068 13190 3096 15846
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3160 14618 3188 14894
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3252 14074 3280 15506
rect 3528 15026 3556 15914
rect 4172 15706 4200 16594
rect 4264 16114 4292 16662
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4356 16250 4384 16594
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4356 15638 4384 16186
rect 4816 16046 4844 16662
rect 5092 16250 5120 16934
rect 6656 16726 6684 17478
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15858 4844 15982
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 4816 15830 4936 15858
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 4172 14958 4200 15302
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 14074 4016 14418
rect 4356 14414 4384 15098
rect 4816 14822 4844 15642
rect 4908 15162 4936 15830
rect 5552 15638 5580 15914
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 3252 13258 3280 13806
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 13530 3372 13670
rect 4816 13530 4844 13806
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2792 11762 2820 12310
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11762 2912 12038
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2792 10810 2820 11698
rect 3068 11218 3096 13126
rect 3884 12368 3936 12374
rect 3882 12336 3884 12345
rect 3936 12336 3938 12345
rect 3882 12271 3938 12280
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3160 11354 3188 11834
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3896 11286 3924 12038
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10810 3280 11086
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2516 9466 2544 10066
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9722 2636 9998
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2516 9450 2636 9466
rect 2516 9444 2648 9450
rect 2516 9438 2596 9444
rect 2596 9386 2648 9392
rect 2608 8974 2636 9386
rect 2700 9178 2728 10066
rect 3252 9722 3280 10542
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10130 3372 10406
rect 3514 10296 3570 10305
rect 3514 10231 3570 10240
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 8430 2636 8910
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2596 7948 2648 7954
rect 2700 7936 2728 8774
rect 2648 7908 2728 7936
rect 2596 7890 2648 7896
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2136 5092 2188 5098
rect 2136 5034 2188 5040
rect 2148 4826 2176 5034
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2424 4826 2452 4966
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2240 4078 2268 4490
rect 2228 4072 2280 4078
rect 2042 4040 2098 4049
rect 2228 4014 2280 4020
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2042 3975 2098 3984
rect 2240 3738 2268 4014
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2516 2774 2544 4014
rect 2424 2746 2544 2774
rect 2424 800 2452 2746
rect 2608 2310 2636 7890
rect 2792 7886 2820 8978
rect 3160 8974 3188 9658
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2884 8090 2912 8910
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2792 5273 2820 6802
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 6390 3004 6734
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3068 6322 3096 6870
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2872 6248 2924 6254
rect 2924 6208 3004 6236
rect 2872 6190 2924 6196
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2700 2650 2728 4694
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 3194 2820 4626
rect 2884 4282 2912 5607
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 3058 2912 3606
rect 2976 3534 3004 6208
rect 3160 5522 3188 8910
rect 3252 7970 3280 9658
rect 3344 8129 3372 10066
rect 3528 9926 3556 10231
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3436 9518 3464 9862
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 9178 3556 9318
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8634 3556 8978
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3330 8120 3386 8129
rect 3330 8055 3386 8064
rect 3252 7942 3464 7970
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7750 3372 7822
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3344 7546 3372 7686
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3436 6066 3464 7942
rect 3620 6254 3648 11154
rect 3884 10192 3936 10198
rect 3790 10160 3846 10169
rect 3884 10134 3936 10140
rect 3790 10095 3846 10104
rect 3698 10024 3754 10033
rect 3698 9959 3754 9968
rect 3712 8430 3740 9959
rect 3804 9058 3832 10095
rect 3896 9178 3924 10134
rect 3988 9654 4016 13330
rect 4080 12889 4108 13398
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4172 12986 4200 13194
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4252 12912 4304 12918
rect 4066 12880 4122 12889
rect 4252 12854 4304 12860
rect 4066 12815 4122 12824
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 4080 11218 4108 11863
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4080 9518 4108 10542
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3804 9030 3924 9058
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 7177 3740 8366
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3698 7168 3754 7177
rect 3698 7103 3754 7112
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3712 6390 3740 6666
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3252 5914 3280 6054
rect 3436 6038 3648 6066
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3160 5494 3280 5522
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2976 3097 3004 3470
rect 3068 3398 3096 4422
rect 3160 3670 3188 4966
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3252 3398 3280 5494
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3344 4282 3372 5170
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3344 3942 3372 4218
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3330 3632 3386 3641
rect 3528 3602 3556 5646
rect 3330 3567 3332 3576
rect 3384 3567 3386 3576
rect 3516 3596 3568 3602
rect 3332 3538 3384 3544
rect 3516 3538 3568 3544
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2962 3088 3018 3097
rect 2872 3052 2924 3058
rect 2962 3023 3018 3032
rect 3240 3052 3292 3058
rect 2872 2994 2924 3000
rect 3240 2994 3292 3000
rect 3252 2854 3280 2994
rect 3344 2961 3372 3538
rect 3514 3496 3570 3505
rect 3514 3431 3570 3440
rect 3424 2984 3476 2990
rect 3330 2952 3386 2961
rect 3528 2938 3556 3431
rect 3476 2932 3556 2938
rect 3424 2926 3556 2932
rect 3436 2910 3556 2926
rect 3330 2887 3386 2896
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2976 1902 3004 2450
rect 3252 2446 3280 2790
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2964 1896 3016 1902
rect 2964 1838 3016 1844
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 2792 800 2820 1362
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 2976 649 3004 1838
rect 3344 1442 3372 2790
rect 3252 1414 3372 1442
rect 3252 800 3280 1414
rect 3528 1057 3556 2910
rect 3514 1048 3570 1057
rect 3514 983 3570 992
rect 2962 640 3018 649
rect 2962 575 3018 584
rect 3238 0 3294 800
rect 3620 241 3648 6038
rect 3712 5778 3740 6326
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3804 5642 3832 7686
rect 3896 5710 3924 9030
rect 3988 7342 4016 9386
rect 4172 8090 4200 12718
rect 4264 12306 4292 12854
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4356 11898 4384 13262
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4908 12434 4936 14486
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 13258 5120 13738
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5000 12442 5028 12650
rect 4816 12406 4936 12434
rect 4988 12436 5040 12442
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4264 11257 4292 11290
rect 4250 11248 4306 11257
rect 4250 11183 4306 11192
rect 4356 10606 4384 11494
rect 4816 11370 4844 12406
rect 4988 12378 5040 12384
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 11626 4936 12174
rect 5000 11762 5028 12378
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4620 11348 4672 11354
rect 4816 11342 5028 11370
rect 4620 11290 4672 11296
rect 4632 11150 4660 11290
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4816 10198 4844 10746
rect 4908 10470 4936 11154
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9518 4384 9998
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4816 9602 4844 9862
rect 4724 9586 4844 9602
rect 4908 9586 4936 10406
rect 5000 9654 5028 11342
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4712 9580 4844 9586
rect 4764 9574 4844 9580
rect 4896 9580 4948 9586
rect 4712 9522 4764 9528
rect 4896 9522 4948 9528
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4264 8430 4292 9454
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4816 9178 4844 9318
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 7744 4120 7750
rect 4066 7712 4068 7721
rect 4120 7712 4122 7721
rect 4066 7647 4122 7656
rect 4356 7342 4384 8978
rect 4988 8968 5040 8974
rect 5092 8956 5120 10746
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10130 5212 10542
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5040 8928 5120 8956
rect 4988 8910 5040 8916
rect 5276 8906 5304 14758
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8090 4844 8774
rect 5276 8294 5304 8842
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4816 7546 4844 7822
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 3988 6225 4016 7278
rect 4356 6882 4384 7278
rect 4080 6854 4384 6882
rect 4080 6769 4108 6854
rect 4160 6792 4212 6798
rect 4066 6760 4122 6769
rect 4448 6746 4476 7278
rect 4908 7206 4936 7890
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4540 7002 4568 7142
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 5368 6934 5396 15370
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 13938 5488 15098
rect 5828 14958 5856 15438
rect 6932 15026 6960 17818
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5828 14618 5856 14894
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6932 14414 6960 14758
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5552 13682 5580 14282
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 5644 13870 5672 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5460 13654 5580 13682
rect 5460 12442 5488 13654
rect 5644 13394 5672 13806
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5448 12436 5500 12442
rect 5552 12434 5580 12786
rect 5736 12782 5764 13670
rect 6012 13394 6040 13670
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6380 13258 6408 13874
rect 6932 13462 6960 14214
rect 7024 14074 7052 17682
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17338 7420 17614
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15162 7144 15846
rect 7208 15366 7236 16050
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 5724 12776 5776 12782
rect 5776 12724 5856 12730
rect 5724 12718 5856 12724
rect 5736 12702 5856 12718
rect 6012 12714 6040 13126
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5552 12406 5672 12434
rect 5448 12378 5500 12384
rect 5460 10810 5488 12378
rect 5644 12306 5672 12406
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10198 5488 10610
rect 5448 10192 5500 10198
rect 5446 10160 5448 10169
rect 5500 10160 5502 10169
rect 5446 10095 5502 10104
rect 5552 9994 5580 11494
rect 5644 11354 5672 12242
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5736 10810 5764 12582
rect 5828 12374 5856 12702
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6196 12374 6224 13126
rect 6380 12850 6408 13194
rect 6932 12850 6960 13398
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5460 9722 5488 9930
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5540 9376 5592 9382
rect 5460 9324 5540 9330
rect 5460 9318 5592 9324
rect 5460 9302 5580 9318
rect 5460 8362 5488 9302
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5460 6798 5488 8298
rect 5644 8090 5672 10542
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10033 5764 10406
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 8430 5764 8774
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 6792 5500 6798
rect 4160 6734 4212 6740
rect 4066 6695 4122 6704
rect 4172 6322 4200 6734
rect 4356 6718 4476 6746
rect 5170 6760 5226 6769
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3974 6216 4030 6225
rect 3974 6151 4030 6160
rect 4172 5846 4200 6258
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 3712 5166 3740 5199
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 3369 3740 5102
rect 3804 4457 3832 5578
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3896 4486 3924 5102
rect 3988 4865 4016 5306
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3974 4856 4030 4865
rect 3974 4791 4030 4800
rect 4080 4690 4108 5170
rect 4356 5166 4384 6718
rect 5448 6734 5500 6740
rect 5552 6746 5580 7754
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7410 5672 7686
rect 5736 7410 5764 8366
rect 5828 8022 5856 8502
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5170 6695 5226 6704
rect 5184 6662 5212 6695
rect 5172 6656 5224 6662
rect 5092 6604 5172 6610
rect 5092 6598 5224 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5092 6582 5212 6598
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4804 6248 4856 6254
rect 4434 6216 4490 6225
rect 4804 6190 4856 6196
rect 4434 6151 4490 6160
rect 4448 5914 4476 6151
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4448 5681 4476 5850
rect 4434 5672 4490 5681
rect 4434 5607 4490 5616
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3884 4480 3936 4486
rect 3790 4448 3846 4457
rect 3884 4422 3936 4428
rect 3790 4383 3846 4392
rect 4080 3738 4108 4626
rect 4264 4486 4292 5034
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3698 3360 3754 3369
rect 3698 3295 3754 3304
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 800 3740 2790
rect 3804 1426 3832 3402
rect 3896 2582 3924 3538
rect 4172 3482 4200 3674
rect 3988 3454 4200 3482
rect 3988 2990 4016 3454
rect 4264 3380 4292 4422
rect 4356 3534 4384 5102
rect 4712 5024 4764 5030
rect 4710 4992 4712 5001
rect 4764 4992 4766 5001
rect 4710 4927 4766 4936
rect 4712 4684 4764 4690
rect 4816 4672 4844 6190
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4908 5166 4936 5782
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4764 4644 4844 4672
rect 4712 4626 4764 4632
rect 4724 4593 4752 4626
rect 4710 4584 4766 4593
rect 4710 4519 4766 4528
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4448 3602 4476 4014
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4080 3352 4292 3380
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4080 2650 4108 3352
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4816 3194 4844 4422
rect 4908 4282 4936 5102
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5000 4162 5028 5850
rect 4908 4134 5028 4162
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4526 3088 4582 3097
rect 4526 3023 4582 3032
rect 4540 2990 4568 3023
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4908 2774 4936 4134
rect 4816 2746 4936 2774
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3884 2576 3936 2582
rect 3976 2576 4028 2582
rect 3884 2518 3936 2524
rect 3974 2544 3976 2553
rect 4028 2544 4030 2553
rect 3974 2479 4030 2488
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4080 2038 4108 2450
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4068 2032 4120 2038
rect 4066 2000 4068 2009
rect 4120 2000 4122 2009
rect 4066 1935 4122 1944
rect 4160 1828 4212 1834
rect 4160 1770 4212 1776
rect 3792 1420 3844 1426
rect 3792 1362 3844 1368
rect 4172 800 4200 1770
rect 4816 1442 4844 2746
rect 5092 2650 5120 6582
rect 5276 5166 5304 6598
rect 5460 5710 5488 6734
rect 5552 6730 5672 6746
rect 5552 6724 5684 6730
rect 5552 6718 5632 6724
rect 5632 6666 5684 6672
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6304 5764 6598
rect 5644 6276 5764 6304
rect 5644 5896 5672 6276
rect 5724 6180 5776 6186
rect 5828 6168 5856 7958
rect 5920 6905 5948 11562
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 9654 6040 11494
rect 6104 11354 6132 12242
rect 6380 12238 6408 12786
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 10044 6132 11290
rect 6184 10056 6236 10062
rect 6104 10016 6184 10044
rect 6184 9998 6236 10004
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 9110 6040 9318
rect 6104 9110 6132 9454
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 5776 6140 5856 6168
rect 5724 6122 5776 6128
rect 5644 5868 5764 5896
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5170 4856 5226 4865
rect 5170 4791 5226 4800
rect 5184 3738 5212 4791
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3670 5304 5102
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4282 5396 4966
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 3754 5488 5102
rect 5552 4826 5580 5510
rect 5644 5370 5672 5714
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4865 5672 4966
rect 5630 4856 5686 4865
rect 5540 4820 5592 4826
rect 5630 4791 5632 4800
rect 5540 4762 5592 4768
rect 5684 4791 5686 4800
rect 5632 4762 5684 4768
rect 5644 4731 5672 4762
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 3942 5580 4490
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5460 3726 5580 3754
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5354 3360 5410 3369
rect 5354 3295 5410 3304
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 4908 1970 4936 2450
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 4988 1760 5040 1766
rect 4988 1702 5040 1708
rect 4632 1414 4844 1442
rect 4632 800 4660 1414
rect 5000 800 5028 1702
rect 5368 1442 5396 3295
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5460 2802 5488 2994
rect 5552 2922 5580 3726
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5644 2802 5672 4626
rect 5736 4146 5764 5868
rect 5906 5400 5962 5409
rect 5906 5335 5908 5344
rect 5960 5335 5962 5344
rect 5908 5306 5960 5312
rect 6012 5166 6040 8298
rect 6104 5778 6132 8298
rect 6196 7886 6224 8978
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6288 6866 6316 9114
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6196 6390 6224 6802
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6288 6202 6316 6802
rect 6196 6174 6316 6202
rect 6196 5914 6224 6174
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5460 2774 5672 2802
rect 5828 2650 5856 4422
rect 5920 3738 5948 4694
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5920 3058 5948 3674
rect 6012 3602 6040 4082
rect 6104 3738 6132 4694
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6196 3913 6224 4626
rect 6288 4554 6316 6054
rect 6380 5914 6408 8366
rect 6472 6322 6500 8434
rect 6564 7750 6592 11766
rect 6748 11218 6776 12174
rect 6932 11665 6960 12582
rect 7116 11898 7144 14962
rect 7208 14550 7236 15302
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6918 11656 6974 11665
rect 6918 11591 6974 11600
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11354 6868 11494
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7024 10266 7052 10542
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6656 7954 6684 9862
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6274 4176 6330 4185
rect 6274 4111 6330 4120
rect 6182 3904 6238 3913
rect 6182 3839 6238 3848
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 3058 6040 3538
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6104 2938 6132 3674
rect 5920 2910 6132 2938
rect 5920 2854 5948 2910
rect 5908 2848 5960 2854
rect 6092 2848 6144 2854
rect 5908 2790 5960 2796
rect 5998 2816 6054 2825
rect 6092 2790 6144 2796
rect 5998 2751 6054 2760
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6012 1442 6040 2751
rect 6104 2582 6132 2790
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6196 2514 6224 3839
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6196 2106 6224 2246
rect 6184 2100 6236 2106
rect 6184 2042 6236 2048
rect 5368 1414 5488 1442
rect 5460 800 5488 1414
rect 5920 1414 6040 1442
rect 6288 1442 6316 4111
rect 6380 2378 6408 4422
rect 6472 4146 6500 6258
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6472 3398 6500 4082
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3126 6500 3334
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6564 1766 6592 6054
rect 6656 4486 6684 7754
rect 6748 6662 6776 10066
rect 7116 9058 7144 10202
rect 7024 9030 7144 9058
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 6866 6868 7414
rect 6932 7274 6960 8230
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6920 6792 6972 6798
rect 7024 6769 7052 9030
rect 7102 8936 7158 8945
rect 7102 8871 7158 8880
rect 7116 7954 7144 8871
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6920 6734 6972 6740
rect 7010 6760 7066 6769
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6932 6254 6960 6734
rect 7010 6695 7066 6704
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 7116 6118 7144 7890
rect 7208 7886 7236 8230
rect 7300 7970 7328 17002
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16658 7512 16934
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8312 16794 8340 17682
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 15638 7420 16390
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7392 15026 7420 15574
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 12986 7420 13670
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7484 12753 7512 16594
rect 8404 16250 8432 17614
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 14822 7604 15302
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7470 12744 7526 12753
rect 7470 12679 7526 12688
rect 7484 12434 7512 12679
rect 7668 12434 7696 14758
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8312 14414 8340 15438
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8312 14006 8340 14350
rect 8588 14074 8616 19246
rect 10612 18970 10640 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8680 15162 8708 18838
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 9600 18426 9628 18770
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 17134 9168 17682
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9508 17134 9536 17614
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8956 16114 8984 17002
rect 9140 16522 9168 17070
rect 9784 16998 9812 17750
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16590 9812 16934
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8772 15706 8800 15846
rect 8956 15706 8984 16050
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9600 15638 9628 16458
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7760 12986 7788 13670
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13530 8248 13874
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7392 12406 7512 12434
rect 7576 12406 7696 12434
rect 7392 10266 7420 12406
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 10810 7512 11494
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7392 9178 7420 10066
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 8974 7512 9930
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8362 7420 8774
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7300 7942 7512 7970
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7410 7236 7822
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6734 5400 6790 5409
rect 6734 5335 6790 5344
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6748 3942 6776 5335
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6656 2825 6684 3062
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6642 2816 6698 2825
rect 6642 2751 6698 2760
rect 6748 2650 6776 2926
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 6288 1414 6408 1442
rect 5920 800 5948 1414
rect 6380 800 6408 1414
rect 6840 800 6868 5850
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7116 5234 7144 5714
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7010 4992 7066 5001
rect 7010 4927 7066 4936
rect 7024 4468 7052 4927
rect 7116 4622 7144 5170
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7024 4440 7144 4468
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 3398 6960 3946
rect 7024 3738 7052 4218
rect 7116 3942 7144 4440
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3618 7144 3878
rect 7024 3590 7144 3618
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 2446 6960 3334
rect 7024 2922 7052 3590
rect 7104 2984 7156 2990
rect 7102 2952 7104 2961
rect 7156 2952 7158 2961
rect 7012 2916 7064 2922
rect 7102 2887 7158 2896
rect 7012 2858 7064 2864
rect 7010 2816 7066 2825
rect 7010 2751 7066 2760
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7024 2310 7052 2751
rect 7208 2650 7236 5238
rect 7392 5166 7420 7754
rect 7484 5914 7512 7942
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7392 3466 7420 3674
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7194 2544 7250 2553
rect 7194 2479 7250 2488
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7208 800 7236 2479
rect 7300 2446 7328 2994
rect 7392 2582 7420 3402
rect 7484 3126 7512 5714
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7576 2310 7604 12406
rect 7760 10130 7788 12582
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12374 8248 13466
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8220 11286 8248 12038
rect 8312 11694 8340 13942
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8404 13394 8432 13806
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12102 8432 13330
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12782 8616 13262
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 10674 8248 11222
rect 8312 11218 8340 11630
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11354 8524 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8392 11280 8444 11286
rect 8390 11248 8392 11257
rect 8444 11248 8446 11257
rect 8300 11212 8352 11218
rect 8390 11183 8446 11192
rect 8300 11154 8352 11160
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8588 10470 8616 12242
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8482 10160 8538 10169
rect 7748 10124 7800 10130
rect 8482 10095 8538 10104
rect 7748 10066 7800 10072
rect 8496 9926 8524 10095
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 7668 9518 7696 9862
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7668 8430 7696 9454
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 8220 8362 8248 9454
rect 8312 9178 8340 9590
rect 8404 9178 8432 9862
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7760 7342 7788 8298
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7342 7972 7958
rect 8312 7818 8340 8910
rect 8588 8498 8616 10406
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8680 8378 8708 8774
rect 8772 8634 8800 15506
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14618 9168 14758
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9876 14498 9904 18158
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 16794 10088 18022
rect 10244 17882 10272 18226
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10888 16726 10916 17818
rect 11072 17202 11100 18090
rect 11256 17882 11284 18770
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11900 17338 11928 17682
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 21362 17232 21418 17241
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 13636 17196 13688 17202
rect 21362 17167 21364 17176
rect 13636 17138 13688 17144
rect 21416 17167 21418 17176
rect 21364 17138 21416 17144
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11716 16130 11744 16390
rect 11624 16102 11744 16130
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15026 9996 15506
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 14618 9996 14962
rect 10152 14822 10180 15982
rect 11624 15502 11652 16102
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10428 14550 10456 14962
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10416 14544 10468 14550
rect 9588 14476 9640 14482
rect 9876 14470 9996 14498
rect 10416 14486 10468 14492
rect 9588 14418 9640 14424
rect 9600 13870 9628 14418
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8956 13530 8984 13670
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 12986 9076 13670
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9232 12850 9260 13738
rect 9876 13530 9904 13806
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8588 8350 8708 8378
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4162 7696 4966
rect 7760 4826 7788 5782
rect 8220 5778 8248 6802
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 5370 7972 5646
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7668 4134 7788 4162
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7668 800 7696 4014
rect 7760 2825 7788 4134
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3738 8248 5510
rect 8312 5370 8340 6054
rect 8404 5710 8432 6394
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8404 5234 8432 5510
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8496 5098 8524 6666
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8392 4684 8444 4690
rect 8588 4672 8616 8350
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8680 5409 8708 6394
rect 8666 5400 8722 5409
rect 8666 5335 8722 5344
rect 8444 4644 8616 4672
rect 8392 4626 8444 4632
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3058 7972 3334
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7746 2816 7802 2825
rect 7746 2751 7802 2760
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 1442 8248 2858
rect 8312 2854 8340 3878
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8312 2446 8340 2790
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8404 1834 8432 4626
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 2990 8524 3878
rect 8576 3528 8628 3534
rect 8680 3516 8708 5335
rect 8772 4690 8800 6598
rect 8864 4826 8892 12650
rect 8956 10062 8984 12786
rect 9218 12744 9274 12753
rect 9218 12679 9274 12688
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10266 9076 10406
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 8945 8984 9522
rect 9140 9160 9168 11018
rect 9232 10130 9260 12679
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 11694 9904 12582
rect 9968 11898 9996 14470
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11218 9812 11494
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9324 9654 9352 10610
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10266 9444 10406
rect 9508 10266 9536 10678
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9588 10192 9640 10198
rect 9586 10160 9588 10169
rect 9640 10160 9642 10169
rect 9586 10095 9642 10104
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9324 9450 9352 9590
rect 9600 9450 9628 9998
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9048 9132 9168 9160
rect 8942 8936 8998 8945
rect 8942 8871 8998 8880
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8628 3488 8708 3516
rect 8576 3470 8628 3476
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2650 8524 2790
rect 8772 2774 8800 4626
rect 8956 3369 8984 7890
rect 9048 7426 9076 9132
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9140 8634 9168 8978
rect 9324 8974 9352 9386
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9232 8430 9260 8774
rect 9416 8498 9444 9046
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9508 7954 9536 8570
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9048 7398 9352 7426
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9232 6254 9260 7210
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 4078 9076 6054
rect 9140 5778 9168 6190
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9324 5030 9352 7398
rect 9416 7342 9444 7822
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9600 7206 9628 9386
rect 9692 9178 9720 10406
rect 9784 10266 9812 10678
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9876 10010 9904 10474
rect 9784 9982 9904 10010
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9692 6866 9720 7890
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9402 6216 9458 6225
rect 9402 6151 9404 6160
rect 9456 6151 9458 6160
rect 9404 6122 9456 6128
rect 9692 5930 9720 6666
rect 9600 5902 9720 5930
rect 9600 5114 9628 5902
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9692 5234 9720 5782
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9600 5086 9720 5114
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4554 9352 4966
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9416 4486 9444 4626
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8942 3360 8998 3369
rect 8942 3295 8998 3304
rect 8588 2746 8800 2774
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8392 1828 8444 1834
rect 8392 1770 8444 1776
rect 8128 1414 8248 1442
rect 8128 800 8156 1414
rect 8588 800 8616 2746
rect 9048 800 9076 3606
rect 9416 800 9444 4422
rect 9600 4078 9628 4558
rect 9692 4185 9720 5086
rect 9784 4826 9812 9982
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9876 5098 9904 9862
rect 9968 9450 9996 9862
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10060 6730 10088 13398
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10244 12850 10272 13330
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9968 4622 9996 5714
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4214 9812 4490
rect 9772 4208 9824 4214
rect 9678 4176 9734 4185
rect 9772 4150 9824 4156
rect 9678 4111 9734 4120
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9772 4072 9824 4078
rect 9968 4060 9996 4558
rect 9824 4032 9996 4060
rect 9772 4014 9824 4020
rect 9678 3768 9734 3777
rect 9678 3703 9680 3712
rect 9732 3703 9734 3712
rect 9680 3674 9732 3680
rect 9692 3534 9720 3674
rect 10060 3602 10088 5102
rect 10152 4826 10180 12582
rect 10244 12442 10272 12786
rect 10232 12436 10284 12442
rect 10796 12434 10824 14758
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 14074 11008 14486
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10796 12406 11008 12434
rect 10232 12378 10284 12384
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11762 10640 12242
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 10810 10456 11494
rect 10612 11354 10640 11698
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10612 10674 10640 11154
rect 10796 11082 10824 11630
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10428 10470 10456 10610
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9784 3194 9812 3538
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9770 3088 9826 3097
rect 9770 3023 9826 3032
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2514 9720 2858
rect 9784 2530 9812 3023
rect 9876 2650 9904 3334
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9680 2508 9732 2514
rect 9784 2502 9904 2530
rect 9680 2450 9732 2456
rect 9876 800 9904 2502
rect 9968 2106 9996 3334
rect 10152 3074 10180 3946
rect 10244 3738 10272 10406
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10520 9450 10548 9930
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10520 8974 10548 9386
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6322 10364 6802
rect 10428 6798 10456 8434
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10520 7954 10548 8230
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7274 10548 7890
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10520 6798 10548 7210
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10428 5778 10456 6122
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10336 4758 10364 5034
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10060 3046 10180 3074
rect 10060 2854 10088 3046
rect 10244 2922 10272 3470
rect 10428 3097 10456 4626
rect 10520 4622 10548 6326
rect 10612 5273 10640 9862
rect 10796 9042 10824 11018
rect 10888 9654 10916 11630
rect 10980 10742 11008 12406
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10980 10044 11008 10678
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10198 11100 10406
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10980 10016 11100 10044
rect 11072 9926 11100 10016
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 7206 10824 8978
rect 10888 8430 10916 9590
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10704 5846 10732 7142
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10796 5794 10824 6258
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5914 10916 6054
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10796 5766 10916 5794
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10598 5264 10654 5273
rect 10796 5234 10824 5510
rect 10598 5199 10654 5208
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10796 4758 10824 5170
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10508 4616 10560 4622
rect 10560 4576 10640 4604
rect 10508 4558 10560 4564
rect 10612 4010 10640 4576
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10414 3088 10470 3097
rect 10612 3058 10640 3946
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10414 3023 10470 3032
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10692 2984 10744 2990
rect 10690 2952 10692 2961
rect 10744 2952 10746 2961
rect 10232 2916 10284 2922
rect 10690 2887 10746 2896
rect 10232 2858 10284 2864
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10140 2848 10192 2854
rect 10692 2848 10744 2854
rect 10140 2790 10192 2796
rect 10690 2816 10692 2825
rect 10744 2816 10746 2825
rect 10060 2446 10088 2790
rect 10152 2650 10180 2790
rect 10690 2751 10746 2760
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 10336 800 10364 1906
rect 10796 800 10824 3674
rect 10888 2990 10916 5766
rect 10980 4078 11008 9318
rect 11072 6390 11100 9862
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5846 11100 6054
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5166 11100 5646
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11164 4826 11192 14826
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11256 12306 11284 13330
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11256 11898 11284 12242
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 11256 8974 11284 9386
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11440 8906 11468 9318
rect 11716 9178 11744 12038
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 6934 11284 7686
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 7410 11744 8230
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5778 11284 6326
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11072 4282 11100 4626
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11072 3924 11100 4218
rect 10980 3896 11100 3924
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10876 2848 10928 2854
rect 10980 2825 11008 3896
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10876 2790 10928 2796
rect 10966 2816 11022 2825
rect 10888 2553 10916 2790
rect 10966 2751 11022 2760
rect 11072 2582 11100 3062
rect 11164 2650 11192 3538
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2576 11112 2582
rect 10874 2544 10930 2553
rect 11060 2518 11112 2524
rect 11256 2514 11284 5306
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11716 4162 11744 6054
rect 11808 5370 11836 15846
rect 12176 13394 12204 16526
rect 12268 16114 12296 17002
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12360 15706 12388 16934
rect 13648 16794 13676 17138
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10606 12020 10950
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 12084 9926 12112 11834
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11900 9518 11928 9862
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11900 7478 11928 8502
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11992 8090 12020 8434
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7546 12020 7890
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11992 7410 12020 7482
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12084 7342 12112 8910
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11900 5778 11928 7210
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6322 12020 6598
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11624 4134 11744 4162
rect 11808 4146 11836 4422
rect 11796 4140 11848 4146
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11532 3466 11560 3946
rect 11624 3670 11652 4134
rect 11796 4082 11848 4088
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 10874 2479 10930 2488
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11348 2360 11376 3062
rect 11256 2332 11376 2360
rect 11256 800 11284 2332
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 800 11744 3946
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 2990 11836 3334
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11900 2854 11928 5714
rect 11992 5710 12020 6258
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12084 5386 12112 7278
rect 11992 5358 12112 5386
rect 11992 4690 12020 5358
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12084 5166 12112 5238
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12084 3738 12112 5102
rect 12176 4554 12204 9046
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6186 12296 6598
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12268 4690 12296 5782
rect 12360 5370 12388 15438
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 7546 12480 8298
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 12084 800 12112 3538
rect 12268 1970 12296 4626
rect 12544 4486 12572 16730
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 19168 11694 19196 12650
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 12912 8430 12940 10474
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 9178 13032 9318
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13096 8634 13124 9454
rect 13280 9382 13308 10066
rect 13556 9722 13584 10134
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 8974 13308 9318
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 13096 6866 13124 8570
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7410 13308 7686
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13372 6866 13400 8502
rect 13556 8430 13584 8774
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6254 13308 6598
rect 13556 6458 13584 7210
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13372 5914 13400 6394
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12636 5166 12664 5646
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12912 5166 12940 5510
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12636 4010 12664 5102
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4758 13124 4966
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13280 4690 13308 5714
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13188 4554 13216 4626
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 2990 12388 3470
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12820 2854 12848 3878
rect 13188 3126 13216 4490
rect 13280 4026 13308 4626
rect 13372 4622 13400 4966
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13280 3998 13400 4026
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3670 13308 3878
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13280 3058 13308 3606
rect 13372 3602 13400 3998
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13556 2990 13584 3334
rect 13648 3126 13676 10474
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 17590 10160 17646 10169
rect 17590 10095 17646 10104
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14568 9178 14596 9386
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8090 14136 8774
rect 15304 8498 15332 8978
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14108 6118 14136 8026
rect 14752 7886 14780 8298
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15396 8090 15424 8230
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 14924 8016 14976 8022
rect 14922 7984 14924 7993
rect 14976 7984 14978 7993
rect 15580 7954 15608 8774
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15764 7954 15792 8230
rect 14922 7919 14978 7928
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14200 6186 14228 6938
rect 14752 6934 14780 7142
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13924 5914 13952 6054
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13740 4826 13768 4966
rect 14108 4826 14136 6054
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14108 4282 14136 4762
rect 14384 4690 14412 6598
rect 14568 5778 14596 6598
rect 14936 6322 14964 6802
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6458 15056 6734
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15580 6118 15608 7890
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13910 4040 13966 4049
rect 13910 3975 13912 3984
rect 13964 3975 13966 3984
rect 13912 3946 13964 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3777 13860 3878
rect 13818 3768 13874 3777
rect 14016 3738 14044 4082
rect 14568 4078 14596 5510
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 13818 3703 13874 3712
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 14292 3058 14320 3878
rect 14660 3194 14688 5102
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14752 4690 14780 4966
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14752 2990 14780 4422
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15396 3602 15424 4966
rect 15580 4690 15608 6054
rect 15856 5778 15884 9658
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 6662 16620 7890
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16592 6322 16620 6598
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5914 16436 6054
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 4758 15700 5170
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15580 4570 15608 4626
rect 15476 4548 15528 4554
rect 15580 4542 15700 4570
rect 15476 4490 15528 4496
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12728 2582 12756 2790
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 12256 1964 12308 1970
rect 12256 1906 12308 1912
rect 12544 800 12572 2314
rect 13004 800 13032 2314
rect 13464 800 13492 2314
rect 13740 2310 13768 2926
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13832 2582 13860 2790
rect 14200 2582 14228 2790
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13924 800 13952 2314
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14292 800 14320 2246
rect 14844 1170 14872 2314
rect 14752 1142 14872 1170
rect 14752 800 14780 1142
rect 15212 800 15240 2858
rect 15488 2582 15516 4490
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 3670 15608 4422
rect 15672 4078 15700 4542
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15672 3738 15700 4014
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15764 3505 15792 5510
rect 15856 5166 15884 5714
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15948 3738 15976 3946
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15750 3496 15806 3505
rect 15750 3431 15806 3440
rect 15948 3058 15976 3674
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15672 800 15700 2858
rect 16040 2582 16068 3878
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 16132 800 16160 3402
rect 16224 2854 16252 4422
rect 16408 4282 16436 4694
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16500 800 16528 2858
rect 16592 1970 16620 4966
rect 16684 2961 16712 5646
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 2990 16804 3470
rect 16960 3058 16988 6802
rect 17132 6316 17184 6322
rect 17236 6304 17264 6802
rect 17184 6276 17264 6304
rect 17132 6258 17184 6264
rect 17144 5710 17172 6258
rect 17604 6254 17632 10095
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17696 7342 17724 7822
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17696 6798 17724 7278
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17512 5914 17540 6054
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 5370 17172 5646
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 17236 4826 17264 5034
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17236 4214 17264 4762
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17420 4146 17448 5238
rect 17696 5166 17724 6734
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17512 4078 17540 4558
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17328 2990 17356 3334
rect 17604 3194 17632 4014
rect 17880 3602 17908 7686
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4690 18552 5102
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17972 2990 18000 3878
rect 16764 2984 16816 2990
rect 16670 2952 16726 2961
rect 16764 2926 16816 2932
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16670 2887 16726 2896
rect 16684 2106 16712 2887
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17972 2582 18000 2790
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 16960 800 16988 2314
rect 17512 1170 17540 2314
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17420 1142 17540 1170
rect 17420 800 17448 1142
rect 17880 800 17908 2246
rect 18064 2038 18092 4422
rect 18156 3641 18184 4422
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18616 4078 18644 6394
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18142 3632 18198 3641
rect 18708 3602 18736 8502
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18142 3567 18198 3576
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18156 2582 18184 3334
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3074 18644 3334
rect 18524 3046 18644 3074
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18524 2514 18552 3046
rect 18800 2990 18828 3878
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18616 2582 18644 2790
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18052 2032 18104 2038
rect 18052 1974 18104 1980
rect 18616 1170 18644 2382
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18340 1142 18644 1170
rect 18340 800 18368 1142
rect 18708 800 18736 2314
rect 19076 1902 19104 3878
rect 19260 3602 19288 4150
rect 19352 3670 19380 11494
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 19064 1896 19116 1902
rect 19064 1838 19116 1844
rect 19168 800 19196 2858
rect 19260 2582 19288 3402
rect 19444 2990 19472 10406
rect 19904 2990 19932 11018
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3584 20576 4014
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20364 3556 20576 3584
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19628 800 19656 2858
rect 20088 800 20116 3402
rect 20364 2650 20392 3556
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20548 800 20576 3402
rect 20640 2582 20668 3674
rect 20732 2990 20760 3946
rect 20824 3670 20852 12038
rect 21362 5808 21418 5817
rect 21362 5743 21364 5752
rect 21416 5743 21418 5752
rect 21364 5714 21416 5720
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 4758 21220 5510
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20916 800 20944 3946
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3602 21404 3878
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21376 2514 21404 3334
rect 21364 2508 21416 2514
rect 21364 2450 21416 2456
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 21192 2106 21220 2246
rect 21180 2100 21232 2106
rect 21180 2042 21232 2048
rect 21376 800 21404 2450
rect 21836 800 21864 4082
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22296 800 22324 2314
rect 22756 800 22784 2926
rect 3606 232 3662 241
rect 3606 167 3662 176
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 2870 22616 2926 22672
rect 2778 21256 2834 21312
rect 2226 20712 2282 20768
rect 2134 20324 2190 20360
rect 2134 20304 2136 20324
rect 2136 20304 2188 20324
rect 2188 20304 2190 20324
rect 4066 22208 4122 22264
rect 3238 21664 3294 21720
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 1582 19796 1584 19816
rect 1584 19796 1636 19816
rect 1636 19796 1638 19816
rect 1582 19760 1638 19796
rect 1582 19352 1638 19408
rect 1582 18844 1584 18864
rect 1584 18844 1636 18864
rect 1636 18844 1638 18864
rect 1582 18808 1638 18844
rect 2226 18420 2282 18456
rect 2226 18400 2228 18420
rect 2228 18400 2280 18420
rect 2280 18400 2282 18420
rect 1674 18028 1676 18048
rect 1676 18028 1728 18048
rect 1728 18028 1730 18048
rect 1674 17992 1730 18028
rect 1674 17484 1676 17504
rect 1676 17484 1728 17504
rect 1728 17484 1730 17504
rect 1674 17448 1730 17484
rect 1582 17060 1638 17096
rect 1582 17040 1584 17060
rect 1584 17040 1636 17060
rect 1636 17040 1638 17060
rect 1582 16496 1638 16552
rect 1582 16124 1584 16144
rect 1584 16124 1636 16144
rect 1636 16124 1638 16144
rect 1582 16088 1638 16124
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 1582 15580 1584 15600
rect 1584 15580 1636 15600
rect 1636 15580 1638 15600
rect 1582 15544 1638 15580
rect 1674 15156 1730 15192
rect 1674 15136 1676 15156
rect 1676 15136 1728 15156
rect 1728 15136 1730 15156
rect 2226 14612 2282 14648
rect 2226 14592 2228 14612
rect 2228 14592 2280 14612
rect 2280 14592 2282 14612
rect 1674 14220 1676 14240
rect 1676 14220 1728 14240
rect 1728 14220 1730 14240
rect 1674 14184 1730 14220
rect 1582 13812 1584 13832
rect 1584 13812 1636 13832
rect 1636 13812 1638 13832
rect 1582 13776 1638 13812
rect 1582 13252 1638 13288
rect 1582 13232 1584 13252
rect 1584 13232 1636 13252
rect 1636 13232 1638 13252
rect 1490 11328 1546 11384
rect 1398 10376 1454 10432
rect 2226 11600 2282 11656
rect 1582 10920 1638 10976
rect 1858 9968 1914 10024
rect 1398 9424 1454 9480
rect 1398 9036 1454 9072
rect 1398 9016 1400 9036
rect 1400 9016 1452 9036
rect 1452 9016 1454 9036
rect 1398 8608 1454 8664
rect 1398 5752 1454 5808
rect 1858 6840 1914 6896
rect 1950 4528 2006 4584
rect 1674 1536 1730 1592
rect 2134 7928 2190 7984
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 3882 12316 3884 12336
rect 3884 12316 3936 12336
rect 3936 12316 3938 12336
rect 3882 12280 3938 12316
rect 3514 10240 3570 10296
rect 2042 3984 2098 4040
rect 2870 5616 2926 5672
rect 2778 5208 2834 5264
rect 3330 8064 3386 8120
rect 3790 10104 3846 10160
rect 3698 9968 3754 10024
rect 4066 12824 4122 12880
rect 4066 11872 4122 11928
rect 3698 7112 3754 7168
rect 3330 3596 3386 3632
rect 3330 3576 3332 3596
rect 3332 3576 3384 3596
rect 3384 3576 3386 3596
rect 2962 3032 3018 3088
rect 3514 3440 3570 3496
rect 3330 2896 3386 2952
rect 3514 992 3570 1048
rect 2962 584 3018 640
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4250 11192 4306 11248
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4066 7692 4068 7712
rect 4068 7692 4120 7712
rect 4120 7692 4122 7712
rect 4066 7656 4122 7692
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4066 6704 4122 6760
rect 5446 10140 5448 10160
rect 5448 10140 5500 10160
rect 5500 10140 5502 10160
rect 5446 10104 5502 10140
rect 5722 9968 5778 10024
rect 3974 6160 4030 6216
rect 3698 5208 3754 5264
rect 3974 4800 4030 4856
rect 5170 6704 5226 6760
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4434 6160 4490 6216
rect 4434 5616 4490 5672
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 3790 4392 3846 4448
rect 3698 3304 3754 3360
rect 4710 4972 4712 4992
rect 4712 4972 4764 4992
rect 4764 4972 4766 4992
rect 4710 4936 4766 4972
rect 4710 4528 4766 4584
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4526 3032 4582 3088
rect 3974 2524 3976 2544
rect 3976 2524 4028 2544
rect 4028 2524 4030 2544
rect 3974 2488 4030 2524
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 4066 1980 4068 2000
rect 4068 1980 4120 2000
rect 4120 1980 4122 2000
rect 4066 1944 4122 1980
rect 5906 6840 5962 6896
rect 5170 4800 5226 4856
rect 5630 4820 5686 4856
rect 5630 4800 5632 4820
rect 5632 4800 5684 4820
rect 5684 4800 5686 4820
rect 5354 3304 5410 3360
rect 5906 5364 5962 5400
rect 5906 5344 5908 5364
rect 5908 5344 5960 5364
rect 5960 5344 5962 5364
rect 6918 11600 6974 11656
rect 6274 4120 6330 4176
rect 6182 3848 6238 3904
rect 5998 2760 6054 2816
rect 7102 8880 7158 8936
rect 7010 6704 7066 6760
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7470 12688 7526 12744
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 6734 5344 6790 5400
rect 6642 2760 6698 2816
rect 7010 4936 7066 4992
rect 7102 2932 7104 2952
rect 7104 2932 7156 2952
rect 7156 2932 7158 2952
rect 7102 2896 7158 2932
rect 7010 2760 7066 2816
rect 7194 2488 7250 2544
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 8390 11228 8392 11248
rect 8392 11228 8444 11248
rect 8444 11228 8446 11248
rect 8390 11192 8446 11228
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8482 10104 8538 10160
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 21362 17196 21418 17232
rect 21362 17176 21364 17196
rect 21364 17176 21416 17196
rect 21416 17176 21418 17196
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8666 5344 8722 5400
rect 7746 2760 7802 2816
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9218 12688 9274 12744
rect 9586 10140 9588 10160
rect 9588 10140 9640 10160
rect 9640 10140 9642 10160
rect 9586 10104 9642 10140
rect 8942 8880 8998 8936
rect 9402 6180 9458 6216
rect 9402 6160 9404 6180
rect 9404 6160 9456 6180
rect 9456 6160 9458 6180
rect 8942 3304 8998 3360
rect 9678 4120 9734 4176
rect 9678 3732 9734 3768
rect 9678 3712 9680 3732
rect 9680 3712 9732 3732
rect 9732 3712 9734 3732
rect 9770 3032 9826 3088
rect 10598 5208 10654 5264
rect 10414 3032 10470 3088
rect 10690 2932 10692 2952
rect 10692 2932 10744 2952
rect 10744 2932 10746 2952
rect 10690 2896 10746 2932
rect 10690 2796 10692 2816
rect 10692 2796 10744 2816
rect 10744 2796 10746 2816
rect 10690 2760 10746 2796
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 10966 2760 11022 2816
rect 10874 2488 10930 2544
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 17590 10104 17646 10160
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14922 7964 14924 7984
rect 14924 7964 14976 7984
rect 14976 7964 14978 7984
rect 14922 7928 14978 7964
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 13910 4004 13966 4040
rect 13910 3984 13912 4004
rect 13912 3984 13964 4004
rect 13964 3984 13966 4004
rect 13818 3712 13874 3768
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15750 3440 15806 3496
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 16670 2896 16726 2952
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18142 3576 18198 3632
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 21362 5772 21418 5808
rect 21362 5752 21364 5772
rect 21364 5752 21416 5772
rect 21416 5752 21418 5772
rect 3606 176 3662 232
<< metal3 >>
rect 0 22674 800 22704
rect 2865 22674 2931 22677
rect 0 22672 2931 22674
rect 0 22616 2870 22672
rect 2926 22616 2931 22672
rect 0 22614 2931 22616
rect 0 22584 800 22614
rect 2865 22611 2931 22614
rect 0 22266 800 22296
rect 4061 22266 4127 22269
rect 0 22264 4127 22266
rect 0 22208 4066 22264
rect 4122 22208 4127 22264
rect 0 22206 4127 22208
rect 0 22176 800 22206
rect 4061 22203 4127 22206
rect 0 21722 800 21752
rect 3233 21722 3299 21725
rect 0 21720 3299 21722
rect 0 21664 3238 21720
rect 3294 21664 3299 21720
rect 0 21662 3299 21664
rect 0 21632 800 21662
rect 3233 21659 3299 21662
rect 0 21314 800 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 800 21254
rect 2773 21251 2839 21254
rect 0 20770 800 20800
rect 2221 20770 2287 20773
rect 0 20768 2287 20770
rect 0 20712 2226 20768
rect 2282 20712 2287 20768
rect 0 20710 2287 20712
rect 0 20680 800 20710
rect 2221 20707 2287 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 2129 20362 2195 20365
rect 0 20360 2195 20362
rect 0 20304 2134 20360
rect 2190 20304 2195 20360
rect 0 20302 2195 20304
rect 0 20272 800 20302
rect 2129 20299 2195 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 800 19758
rect 1577 19755 1643 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 2221 18458 2287 18461
rect 0 18456 2287 18458
rect 0 18400 2226 18456
rect 2282 18400 2287 18456
rect 0 18398 2287 18400
rect 0 18368 800 18398
rect 2221 18395 2287 18398
rect 0 18050 800 18080
rect 1669 18050 1735 18053
rect 0 18048 1735 18050
rect 0 17992 1674 18048
rect 1730 17992 1735 18048
rect 0 17990 1735 17992
rect 0 17960 800 17990
rect 1669 17987 1735 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 0 17506 800 17536
rect 1669 17506 1735 17509
rect 0 17504 1735 17506
rect 0 17448 1674 17504
rect 1730 17448 1735 17504
rect 0 17446 1735 17448
rect 0 17416 800 17446
rect 1669 17443 1735 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 21357 17234 21423 17237
rect 22200 17234 23000 17264
rect 21357 17232 23000 17234
rect 21357 17176 21362 17232
rect 21418 17176 23000 17232
rect 21357 17174 23000 17176
rect 21357 17171 21423 17174
rect 22200 17144 23000 17174
rect 0 17098 800 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 800 17038
rect 1577 17035 1643 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 800 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 800 16494
rect 1577 16491 1643 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 1577 15602 1643 15605
rect 0 15600 1643 15602
rect 0 15544 1582 15600
rect 1638 15544 1643 15600
rect 0 15542 1643 15544
rect 0 15512 800 15542
rect 1577 15539 1643 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 800 15134
rect 1669 15131 1735 15134
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 2221 14650 2287 14653
rect 0 14648 2287 14650
rect 0 14592 2226 14648
rect 2282 14592 2287 14648
rect 0 14590 2287 14592
rect 0 14560 800 14590
rect 2221 14587 2287 14590
rect 0 14242 800 14272
rect 1669 14242 1735 14245
rect 0 14240 1735 14242
rect 0 14184 1674 14240
rect 1730 14184 1735 14240
rect 0 14182 1735 14184
rect 0 14152 800 14182
rect 1669 14179 1735 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 4061 12882 4127 12885
rect 0 12880 4127 12882
rect 0 12824 4066 12880
rect 4122 12824 4127 12880
rect 0 12822 4127 12824
rect 0 12792 800 12822
rect 4061 12819 4127 12822
rect 7465 12746 7531 12749
rect 9213 12746 9279 12749
rect 7465 12744 9279 12746
rect 7465 12688 7470 12744
rect 7526 12688 9218 12744
rect 9274 12688 9279 12744
rect 7465 12686 9279 12688
rect 7465 12683 7531 12686
rect 9213 12683 9279 12686
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12338 800 12368
rect 3877 12338 3943 12341
rect 0 12336 3943 12338
rect 0 12280 3882 12336
rect 3938 12280 3943 12336
rect 0 12278 3943 12280
rect 0 12248 800 12278
rect 3877 12275 3943 12278
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 4061 11930 4127 11933
rect 0 11928 4127 11930
rect 0 11872 4066 11928
rect 4122 11872 4127 11928
rect 0 11870 4127 11872
rect 0 11840 800 11870
rect 4061 11867 4127 11870
rect 2221 11658 2287 11661
rect 6913 11658 6979 11661
rect 2221 11656 6979 11658
rect 2221 11600 2226 11656
rect 2282 11600 6918 11656
rect 6974 11600 6979 11656
rect 2221 11598 6979 11600
rect 2221 11595 2287 11598
rect 6913 11595 6979 11598
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 4245 11250 4311 11253
rect 8385 11250 8451 11253
rect 4245 11248 8451 11250
rect 4245 11192 4250 11248
rect 4306 11192 8390 11248
rect 8446 11192 8451 11248
rect 4245 11190 8451 11192
rect 4245 11187 4311 11190
rect 8385 11187 8451 11190
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 3509 10298 3575 10301
rect 3509 10296 7666 10298
rect 3509 10240 3514 10296
rect 3570 10240 7666 10296
rect 3509 10238 7666 10240
rect 3509 10235 3575 10238
rect 3785 10162 3851 10165
rect 5441 10162 5507 10165
rect 3785 10160 5507 10162
rect 3785 10104 3790 10160
rect 3846 10104 5446 10160
rect 5502 10104 5507 10160
rect 3785 10102 5507 10104
rect 7606 10162 7666 10238
rect 8477 10162 8543 10165
rect 7606 10160 8543 10162
rect 7606 10104 8482 10160
rect 8538 10104 8543 10160
rect 7606 10102 8543 10104
rect 3785 10099 3851 10102
rect 5441 10099 5507 10102
rect 8477 10099 8543 10102
rect 9581 10162 9647 10165
rect 17585 10162 17651 10165
rect 9581 10160 17651 10162
rect 9581 10104 9586 10160
rect 9642 10104 17590 10160
rect 17646 10104 17651 10160
rect 9581 10102 17651 10104
rect 9581 10099 9647 10102
rect 17585 10099 17651 10102
rect 0 10026 800 10056
rect 1853 10026 1919 10029
rect 0 10024 1919 10026
rect 0 9968 1858 10024
rect 1914 9968 1919 10024
rect 0 9966 1919 9968
rect 0 9936 800 9966
rect 1853 9963 1919 9966
rect 3693 10026 3759 10029
rect 5717 10026 5783 10029
rect 3693 10024 5783 10026
rect 3693 9968 3698 10024
rect 3754 9968 5722 10024
rect 5778 9968 5783 10024
rect 3693 9966 5783 9968
rect 3693 9963 3759 9966
rect 5717 9963 5783 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 7097 8938 7163 8941
rect 8937 8938 9003 8941
rect 7097 8936 9003 8938
rect 7097 8880 7102 8936
rect 7158 8880 8942 8936
rect 8998 8880 9003 8936
rect 7097 8878 9003 8880
rect 7097 8875 7163 8878
rect 8937 8875 9003 8878
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 1393 8666 1459 8669
rect 0 8664 1459 8666
rect 0 8608 1398 8664
rect 1454 8608 1459 8664
rect 0 8606 1459 8608
rect 0 8576 800 8606
rect 1393 8603 1459 8606
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 3325 8122 3391 8125
rect 0 8120 3391 8122
rect 0 8064 3330 8120
rect 3386 8064 3391 8120
rect 0 8062 3391 8064
rect 0 8032 800 8062
rect 3325 8059 3391 8062
rect 2129 7986 2195 7989
rect 14917 7986 14983 7989
rect 2129 7984 14983 7986
rect 2129 7928 2134 7984
rect 2190 7928 14922 7984
rect 14978 7928 14983 7984
rect 2129 7926 14983 7928
rect 2129 7923 2195 7926
rect 14917 7923 14983 7926
rect 0 7714 800 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 800 7654
rect 4061 7651 4127 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 0 7170 800 7200
rect 3693 7170 3759 7173
rect 0 7168 3759 7170
rect 0 7112 3698 7168
rect 3754 7112 3759 7168
rect 0 7110 3759 7112
rect 0 7080 800 7110
rect 3693 7107 3759 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 1853 6898 1919 6901
rect 5901 6898 5967 6901
rect 1853 6896 5967 6898
rect 1853 6840 1858 6896
rect 1914 6840 5906 6896
rect 5962 6840 5967 6896
rect 1853 6838 5967 6840
rect 1853 6835 1919 6838
rect 5901 6835 5967 6838
rect 0 6762 800 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 800 6702
rect 4061 6699 4127 6702
rect 5165 6762 5231 6765
rect 7005 6762 7071 6765
rect 5165 6760 7071 6762
rect 5165 6704 5170 6760
rect 5226 6704 7010 6760
rect 7066 6704 7071 6760
rect 5165 6702 7071 6704
rect 5165 6699 5231 6702
rect 7005 6699 7071 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 800 6158
rect 3969 6155 4035 6158
rect 4429 6218 4495 6221
rect 9397 6218 9463 6221
rect 4429 6216 9463 6218
rect 4429 6160 4434 6216
rect 4490 6160 9402 6216
rect 9458 6160 9463 6216
rect 4429 6158 9463 6160
rect 4429 6155 4495 6158
rect 9397 6155 9463 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 21357 5810 21423 5813
rect 22200 5810 23000 5840
rect 21357 5808 23000 5810
rect 21357 5752 21362 5808
rect 21418 5752 23000 5808
rect 21357 5750 23000 5752
rect 21357 5747 21423 5750
rect 22200 5720 23000 5750
rect 2865 5674 2931 5677
rect 4429 5674 4495 5677
rect 2865 5672 4495 5674
rect 2865 5616 2870 5672
rect 2926 5616 4434 5672
rect 4490 5616 4495 5672
rect 2865 5614 4495 5616
rect 2865 5611 2931 5614
rect 4429 5611 4495 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 5901 5402 5967 5405
rect 6729 5402 6795 5405
rect 8661 5402 8727 5405
rect 5901 5400 8727 5402
rect 5901 5344 5906 5400
rect 5962 5344 6734 5400
rect 6790 5344 8666 5400
rect 8722 5344 8727 5400
rect 5901 5342 8727 5344
rect 5901 5339 5967 5342
rect 6729 5339 6795 5342
rect 8661 5339 8727 5342
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 3693 5266 3759 5269
rect 10593 5266 10659 5269
rect 3693 5264 10659 5266
rect 3693 5208 3698 5264
rect 3754 5208 10598 5264
rect 10654 5208 10659 5264
rect 3693 5206 10659 5208
rect 3693 5203 3759 5206
rect 10593 5203 10659 5206
rect 4705 4994 4771 4997
rect 7005 4994 7071 4997
rect 4705 4992 7071 4994
rect 4705 4936 4710 4992
rect 4766 4936 7010 4992
rect 7066 4936 7071 4992
rect 4705 4934 7071 4936
rect 4705 4931 4771 4934
rect 7005 4931 7071 4934
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 800 4798
rect 3969 4795 4035 4798
rect 5165 4858 5231 4861
rect 5625 4858 5691 4861
rect 5165 4856 5691 4858
rect 5165 4800 5170 4856
rect 5226 4800 5630 4856
rect 5686 4800 5691 4856
rect 5165 4798 5691 4800
rect 5165 4795 5231 4798
rect 5625 4795 5691 4798
rect 1945 4586 2011 4589
rect 4705 4586 4771 4589
rect 1945 4584 4771 4586
rect 1945 4528 1950 4584
rect 2006 4528 4710 4584
rect 4766 4528 4771 4584
rect 1945 4526 4771 4528
rect 1945 4523 2011 4526
rect 4705 4523 4771 4526
rect 0 4450 800 4480
rect 3785 4450 3851 4453
rect 0 4448 3851 4450
rect 0 4392 3790 4448
rect 3846 4392 3851 4448
rect 0 4390 3851 4392
rect 0 4360 800 4390
rect 3785 4387 3851 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 6269 4178 6335 4181
rect 9673 4178 9739 4181
rect 6269 4176 9739 4178
rect 6269 4120 6274 4176
rect 6330 4120 9678 4176
rect 9734 4120 9739 4176
rect 6269 4118 9739 4120
rect 6269 4115 6335 4118
rect 9673 4115 9739 4118
rect 2037 4042 2103 4045
rect 13905 4042 13971 4045
rect 2037 4040 13971 4042
rect 2037 3984 2042 4040
rect 2098 3984 13910 4040
rect 13966 3984 13971 4040
rect 2037 3982 13971 3984
rect 2037 3979 2103 3982
rect 13905 3979 13971 3982
rect 0 3906 800 3936
rect 6177 3906 6243 3909
rect 0 3904 6243 3906
rect 0 3848 6182 3904
rect 6238 3848 6243 3904
rect 0 3846 6243 3848
rect 0 3816 800 3846
rect 6177 3843 6243 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 9673 3770 9739 3773
rect 13813 3770 13879 3773
rect 9673 3768 13879 3770
rect 9673 3712 9678 3768
rect 9734 3712 13818 3768
rect 13874 3712 13879 3768
rect 9673 3710 13879 3712
rect 9673 3707 9739 3710
rect 13813 3707 13879 3710
rect 3325 3634 3391 3637
rect 18137 3634 18203 3637
rect 3325 3632 18203 3634
rect 3325 3576 3330 3632
rect 3386 3576 18142 3632
rect 18198 3576 18203 3632
rect 3325 3574 18203 3576
rect 3325 3571 3391 3574
rect 18137 3571 18203 3574
rect 0 3498 800 3528
rect 3509 3498 3575 3501
rect 15745 3498 15811 3501
rect 0 3438 2790 3498
rect 0 3408 800 3438
rect 2730 3362 2790 3438
rect 3509 3496 15811 3498
rect 3509 3440 3514 3496
rect 3570 3440 15750 3496
rect 15806 3440 15811 3496
rect 3509 3438 15811 3440
rect 3509 3435 3575 3438
rect 15745 3435 15811 3438
rect 3693 3362 3759 3365
rect 2730 3360 3759 3362
rect 2730 3304 3698 3360
rect 3754 3304 3759 3360
rect 2730 3302 3759 3304
rect 3693 3299 3759 3302
rect 5349 3362 5415 3365
rect 8937 3362 9003 3365
rect 5349 3360 9003 3362
rect 5349 3304 5354 3360
rect 5410 3304 8942 3360
rect 8998 3304 9003 3360
rect 5349 3302 9003 3304
rect 5349 3299 5415 3302
rect 8937 3299 9003 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 2957 3090 3023 3093
rect 4521 3090 4587 3093
rect 2957 3088 4587 3090
rect 2957 3032 2962 3088
rect 3018 3032 4526 3088
rect 4582 3032 4587 3088
rect 2957 3030 4587 3032
rect 2957 3027 3023 3030
rect 4521 3027 4587 3030
rect 9765 3090 9831 3093
rect 10409 3090 10475 3093
rect 9765 3088 10475 3090
rect 9765 3032 9770 3088
rect 9826 3032 10414 3088
rect 10470 3032 10475 3088
rect 9765 3030 10475 3032
rect 9765 3027 9831 3030
rect 10409 3027 10475 3030
rect 0 2954 800 2984
rect 3325 2954 3391 2957
rect 0 2952 3391 2954
rect 0 2896 3330 2952
rect 3386 2896 3391 2952
rect 0 2894 3391 2896
rect 0 2864 800 2894
rect 3325 2891 3391 2894
rect 7097 2954 7163 2957
rect 10685 2954 10751 2957
rect 16665 2954 16731 2957
rect 7097 2952 16731 2954
rect 7097 2896 7102 2952
rect 7158 2896 10690 2952
rect 10746 2896 16670 2952
rect 16726 2896 16731 2952
rect 7097 2894 16731 2896
rect 7097 2891 7163 2894
rect 10685 2891 10751 2894
rect 16665 2891 16731 2894
rect 5993 2818 6059 2821
rect 6637 2818 6703 2821
rect 5993 2816 6703 2818
rect 5993 2760 5998 2816
rect 6054 2760 6642 2816
rect 6698 2760 6703 2816
rect 5993 2758 6703 2760
rect 5993 2755 6059 2758
rect 6637 2755 6703 2758
rect 7005 2818 7071 2821
rect 7741 2818 7807 2821
rect 7005 2816 7807 2818
rect 7005 2760 7010 2816
rect 7066 2760 7746 2816
rect 7802 2760 7807 2816
rect 7005 2758 7807 2760
rect 7005 2755 7071 2758
rect 7741 2755 7807 2758
rect 10685 2818 10751 2821
rect 10961 2818 11027 2821
rect 10685 2816 11027 2818
rect 10685 2760 10690 2816
rect 10746 2760 10966 2816
rect 11022 2760 11027 2816
rect 10685 2758 11027 2760
rect 10685 2755 10751 2758
rect 10961 2755 11027 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 3969 2546 4035 2549
rect 0 2544 4035 2546
rect 0 2488 3974 2544
rect 4030 2488 4035 2544
rect 0 2486 4035 2488
rect 0 2456 800 2486
rect 3969 2483 4035 2486
rect 7189 2546 7255 2549
rect 10869 2546 10935 2549
rect 7189 2544 10935 2546
rect 7189 2488 7194 2544
rect 7250 2488 10874 2544
rect 10930 2488 10935 2544
rect 7189 2486 10935 2488
rect 7189 2483 7255 2486
rect 10869 2483 10935 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 4061 2002 4127 2005
rect 0 2000 4127 2002
rect 0 1944 4066 2000
rect 4122 1944 4127 2000
rect 0 1942 4127 1944
rect 0 1912 800 1942
rect 4061 1939 4127 1942
rect 0 1594 800 1624
rect 1669 1594 1735 1597
rect 0 1592 1735 1594
rect 0 1536 1674 1592
rect 1730 1536 1735 1592
rect 0 1534 1735 1536
rect 0 1504 800 1534
rect 1669 1531 1735 1534
rect 0 1050 800 1080
rect 3509 1050 3575 1053
rect 0 1048 3575 1050
rect 0 992 3514 1048
rect 3570 992 3575 1048
rect 0 990 3575 992
rect 0 960 800 990
rect 3509 987 3575 990
rect 0 642 800 672
rect 2957 642 3023 645
rect 0 640 3023 642
rect 0 584 2962 640
rect 3018 584 3023 640
rect 0 582 3023 584
rect 0 552 800 582
rect 2957 579 3023 582
rect 0 234 800 264
rect 3601 234 3667 237
rect 0 232 3667 234
rect 0 176 3606 232
rect 3662 176 3667 232
rect 0 174 3667 176
rect 0 144 800 174
rect 3601 171 3667 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1624635492
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1624635492
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2944 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2668 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_20
timestamp 1624635492
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 4600 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1624635492
transform -1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1624635492
transform -1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1624635492
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1624635492
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_38
timestamp 1624635492
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1624635492
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5336 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 6256 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform -1 0 6164 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1624635492
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6716 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10120 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8924 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1624635492
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74
timestamp 1624635492
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1624635492
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1624635492
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10304 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9476 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 10764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1624635492
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1624635492
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1624635492
transform 1 0 11500 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_109
timestamp 1624635492
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1624635492
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1624635492
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1624635492
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11592 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1624635492
transform 1 0 12144 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1624635492
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform -1 0 12328 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 12144 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 12880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13340 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_128
timestamp 1624635492
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1624635492
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1624635492
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1624635492
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 13800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp 1624635492
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1624635492
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140
timestamp 1624635492
transform 1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1624635492
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_152
timestamp 1624635492
transform 1 0 15088 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 15088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15916 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1624635492
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1624635492
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_158
timestamp 1624635492
transform 1 0 15640 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 16192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1624635492
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1624635492
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1624635492
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1624635492
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_183
timestamp 1624635492
transform 1 0 17940 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform 1 0 18124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1624635492
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform 1 0 18584 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_193
timestamp 1624635492
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1624635492
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 19504 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1624635492
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1624635492
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_206
timestamp 1624635492
transform 1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform -1 0 20332 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21436 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform -1 0 21436 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1624635492
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1624635492
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1624635492
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1624635492
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 2944 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1624635492
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1624635492
transform -1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1624635492
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1624635492
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6164 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_53
timestamp 1624635492
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1624635492
transform 1 0 7636 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1624635492
transform 1 0 10672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 9292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1624635492
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_89
timestamp 1624635492
transform 1 0 9292 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1624635492
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1624635492
transform -1 0 12420 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12604 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1624635492
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp 1624635492
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1624635492
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 16560 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1624635492
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1624635492
transform 1 0 16744 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform -1 0 17940 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 18400 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_168
timestamp 1624635492
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1624635492
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_178
timestamp 1624635492
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1624635492
transform 1 0 17940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1624635492
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform 1 0 18584 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1624635492
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 19044 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_198
timestamp 1624635492
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1624635492
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform 1 0 21160 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 20976 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1624635492
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_216
timestamp 1624635492
transform 1 0 20976 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 1932 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1624635492
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1624635492
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5244 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1624635492
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_54
timestamp 1624635492
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9752 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1624635492
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1624635492
transform 1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11408 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1624635492
transform 1 0 10212 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11868 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1624635492
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14352 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1624635492
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1624635492
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14996 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1624635492
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18400 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17940 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1624635492
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1624635492
transform 1 0 17940 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1624635492
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1624635492
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1624635492
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_201
timestamp 1624635492
transform 1 0 19596 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1624635492
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1624635492
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 20700 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 21252 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1624635492
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1624635492
transform 1 0 21252 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2208 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_12
timestamp 1624635492
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform -1 0 4784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1624635492
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1624635492
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_40
timestamp 1624635492
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform 1 0 6164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1624635492
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1624635492
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1624635492
transform -1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform -1 0 8832 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1624635492
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1624635492
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1624635492
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1624635492
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10488 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1624635492
transform -1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624635492
transform -1 0 10120 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1624635492
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1624635492
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1624635492
transform 1 0 10120 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1624635492
transform -1 0 12420 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1624635492
transform -1 0 12880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 1624635492
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1624635492
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1624635492
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_128
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp 1624635492
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_139
timestamp 1624635492
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform -1 0 15640 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 15180 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1624635492
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1624635492
transform 1 0 15180 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1624635492
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1624635492
transform 1 0 17480 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 18124 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1624635492
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1624635492
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_185
timestamp 1624635492
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 21436 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1624635492
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 18860 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1624635492
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1624635492
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1624635492
transform -1 0 3220 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1624635492
transform 1 0 1564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1624635492
transform 1 0 1932 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_13
timestamp 1624635492
transform 1 0 2300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1624635492
transform 1 0 3404 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 3864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 4784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1624635492
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1624635492
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_33
timestamp 1624635492
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1624635492
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform 1 0 5244 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 6624 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1624635492
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1624635492
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1624635492
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1624635492
transform 1 0 6624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1624635492
transform -1 0 8832 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1624635492
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1624635492
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_88
timestamp 1624635492
transform 1 0 9200 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1624635492
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1624635492
transform -1 0 12144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 12604 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_109
timestamp 1624635492
transform 1 0 11132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1624635492
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1624635492
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp 1624635492
transform 1 0 12604 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1624635492
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1624635492
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1624635492
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_143
timestamp 1624635492
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16284 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1624635492
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_153
timestamp 1624635492
transform 1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1624635492
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18584 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1624635492
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 18584 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1624635492
transform 1 0 19688 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 20792 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1624635492
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 2852 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_5
timestamp 1624635492
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_16
timestamp 1624635492
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1624635492
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp 1624635492
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1624635492
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1624635492
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6072 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_51
timestamp 1624635492
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1624635492
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624635492
transform 1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1624635492
transform -1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1624635492
transform 1 0 6624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1624635492
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 6624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5980 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8464 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8464 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1624635492
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_80
timestamp 1624635492
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1624635492
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9384 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10948 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1624635492
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1624635492
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1624635492
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1624635492
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1624635492
transform -1 0 11776 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1624635492
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_117
timestamp 1624635492
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_116
timestamp 1624635492
transform 1 0 11776 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12880 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12144 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1624635492
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1624635492
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform 1 0 13064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1624635492
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1624635492
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14628 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp 1624635492
transform 1 0 15088 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 1624635492
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_153
timestamp 1624635492
transform 1 0 15180 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1624635492
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 15180 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 15640 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1624635492
transform -1 0 15088 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1624635492
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_165
timestamp 1624635492
transform 1 0 16284 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_161
timestamp 1624635492
transform 1 0 15916 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1624635492
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16652 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16376 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1624635492
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1624635492
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1624635492
transform -1 0 17664 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_183
timestamp 1624635492
transform 1 0 17940 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_184
timestamp 1624635492
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_180
timestamp 1624635492
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 18400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_187
timestamp 1624635492
transform 1 0 18308 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_188
timestamp 1624635492
transform 1 0 18400 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_199
timestamp 1624635492
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624635492
transform 1 0 21160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1624635492
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_216
timestamp 1624635492
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1624635492
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1624635492
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 1748 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_5
timestamp 1624635492
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1624635492
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5520 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1624635492
transform -1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1624635492
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1624635492
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1624635492
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_58
timestamp 1624635492
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1624635492
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1624635492
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1624635492
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1624635492
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_92
timestamp 1624635492
transform 1 0 9568 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1624635492
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1624635492
transform -1 0 9568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1624635492
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1624635492
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1624635492
transform -1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10580 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 1624635492
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1624635492
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1624635492
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1624635492
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1624635492
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1624635492
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17572 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14536 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp 1624635492
transform 1 0 15364 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_160
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_179
timestamp 1624635492
transform 1 0 17572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_191
timestamp 1624635492
transform 1 0 18676 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_199
timestamp 1624635492
transform 1 0 19412 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1624635492
transform 1 0 20700 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1624635492
transform 1 0 21436 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1748 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_5
timestamp 1624635492
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1624635492
transform -1 0 3680 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624635492
transform -1 0 4140 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1624635492
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1624635492
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_28
timestamp 1624635492
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 1624635492
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1624635492
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6624 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp 1624635492
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1624635492
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1624635492
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1624635492
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12696 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_105
timestamp 1624635492
transform 1 0 10764 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13340 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_126
timestamp 1624635492
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_130
timestamp 1624635492
transform 1 0 13064 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16468 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1624635492
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1624635492
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_174
timestamp 1624635492
transform 1 0 17112 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_186
timestamp 1624635492
transform 1 0 18216 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_198
timestamp 1624635492
transform 1 0 19320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_210
timestamp 1624635492
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1624635492
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1624635492
transform -1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_5
timestamp 1624635492
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1624635492
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 4140 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_33
timestamp 1624635492
transform 1 0 4140 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5336 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform -1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1624635492
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_44
timestamp 1624635492
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1624635492
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1624635492
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8096 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1624635492
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1624635492
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1624635492
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_81
timestamp 1624635492
transform 1 0 8556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10488 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1624635492
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_98
timestamp 1624635492
transform 1 0 10120 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13616 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_118
timestamp 1624635492
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1624635492
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1624635492
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17664 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15364 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1624635492
transform 1 0 15364 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 1624635492
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1624635492
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1624635492
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1624635492
transform 1 0 20700 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1624635492
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 1932 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_6
timestamp 1624635492
transform 1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4324 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624635492
transform -1 0 3864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 1624635492
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1624635492
transform 1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_34
timestamp 1624635492
transform 1 0 4232 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 6624 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_51
timestamp 1624635492
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1624635492
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_60
timestamp 1624635492
transform 1 0 6624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1624635492
transform -1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1624635492
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1624635492
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1624635492
transform 1 0 9384 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1624635492
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1624635492
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12696 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1624635492
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_109
timestamp 1624635492
transform 1 0 11132 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13432 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1624635492
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_131
timestamp 1624635492
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15916 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1624635492
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1624635492
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1624635492
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1624635492
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_177
timestamp 1624635492
transform 1 0 17388 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_189
timestamp 1624635492
transform 1 0 18492 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1624635492
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1624635492
transform 1 0 20700 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1624635492
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1624635492
transform -1 0 2208 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3220 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_6
timestamp 1624635492
transform 1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_12
timestamp 1624635492
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1624635492
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1624635492
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6900 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1624635492
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1624635492
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1624635492
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1624635492
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_83
timestamp 1624635492
transform 1 0 8740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_89
timestamp 1624635492
transform 1 0 9292 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1624635492
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11868 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12880 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1624635492
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1624635492
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1624635492
transform 1 0 13064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1624635492
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1624635492
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1624635492
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16008 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_162
timestamp 1624635492
transform 1 0 16008 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_174
timestamp 1624635492
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_186
timestamp 1624635492
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1624635492
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_213
timestamp 1624635492
transform 1 0 20700 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1624635492
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1624635492
transform -1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1624635492
transform 1 0 1840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1624635492
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1624635492
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1624635492
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1624635492
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform -1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1624635492
transform -1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1624635492
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_32
timestamp 1624635492
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4232 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform -1 0 4416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_47
timestamp 1624635492
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1624635492
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1624635492
transform 1 0 5060 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1624635492
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_58
timestamp 1624635492
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_60
timestamp 1624635492
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1624635492
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8280 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 8464 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1624635492
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1624635492
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1624635492
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1624635492
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9384 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_103
timestamp 1624635492
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 1624635492
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10764 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1624635492
transform 1 0 11316 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1624635492
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1624635492
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1624635492
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13156 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 13708 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1624635492
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1624635492
transform 1 0 13708 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_131
timestamp 1624635492
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1624635492
transform 1 0 14812 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_161
timestamp 1624635492
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1624635492
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1624635492
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1624635492
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1624635492
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1624635492
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1624635492
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1624635492
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1624635492
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1624635492
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1624635492
transform 1 0 20700 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1624635492
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1656 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1624635492
transform -1 0 3588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1624635492
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1624635492
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 6624 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1624635492
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1624635492
transform 1 0 5888 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1624635492
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1624635492
transform 1 0 6624 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7360 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_65
timestamp 1624635492
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1624635492
transform 1 0 8188 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9016 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1624635492
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1624635492
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13708 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1624635492
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1624635492
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1624635492
transform 1 0 13708 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1624635492
transform 1 0 14812 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_161
timestamp 1624635492
transform 1 0 15916 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _106_
timestamp 1624635492
transform 1 0 18216 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1624635492
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1624635492
transform -1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1624635492
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1624635492
transform 1 0 18860 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1624635492
transform 1 0 19964 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1624635492
transform 1 0 21068 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1624635492
transform 1 0 2208 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1624635492
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1624635492
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4600 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1624635492
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_26
timestamp 1624635492
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_35
timestamp 1624635492
transform 1 0 4324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform -1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7084 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1624635492
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_81
timestamp 1624635492
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9476 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_89
timestamp 1624635492
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1624635492
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1624635492
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1624635492
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1624635492
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1624635492
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1624635492
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1624635492
transform 1 0 17664 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _107_
timestamp 1624635492
transform 1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_188
timestamp 1624635492
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_194
timestamp 1624635492
transform 1 0 18952 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_213
timestamp 1624635492
transform 1 0 20700 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2944 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1624635492
transform -1 0 2760 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform -1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1624635492
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_18
timestamp 1624635492
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1624635492
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 6624 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_47
timestamp 1624635492
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1624635492
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1624635492
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_60
timestamp 1624635492
transform 1 0 6624 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8280 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1624635492
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1624635492
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_94
timestamp 1624635492
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 12144 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1624635492
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1624635492
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_120
timestamp 1624635492
transform 1 0 12144 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_132
timestamp 1624635492
transform 1 0 13248 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1624635492
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1624635492
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_168
timestamp 1624635492
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1624635492
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1624635492
transform 1 0 19136 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_199
timestamp 1624635492
transform 1 0 19412 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_211
timestamp 1624635492
transform 1 0 20516 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3312 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1624635492
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1624635492
transform -1 0 4784 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1624635492
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1624635492
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_35
timestamp 1624635492
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1624635492
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6440 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_58
timestamp 1624635492
transform 1 0 6440 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_82
timestamp 1624635492
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11316 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_89
timestamp 1624635492
transform 1 0 9292 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1624635492
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1624635492
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1624635492
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1624635492
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1624635492
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1624635492
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1624635492
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1624635492
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_206
timestamp 1624635492
transform 1 0 20056 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1624635492
transform 1 0 21160 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1624635492
transform 1 0 21528 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1624635492
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_5
timestamp 1624635492
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1624635492
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1624635492
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1624635492
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3036 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 2576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1624635492
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1624635492
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1624635492
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1624635492
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1624635492
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_40
timestamp 1624635492
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_35
timestamp 1624635492
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 5612 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1624635492
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1624635492
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 5796 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4968 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1624635492
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1624635492
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 6440 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform -1 0 7544 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7728 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1624635492
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1624635492
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1624635492
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1624635492
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_85
timestamp 1624635492
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform 1 0 9384 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_101
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11316 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624635492
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1624635492
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1624635492
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1624635492
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1624635492
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1624635492
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1624635492
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1624635492
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1624635492
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_213
timestamp 1624635492
transform 1 0 20700 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1624635492
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1624635492
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1624635492
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5428 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1624635492
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1624635492
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1624635492
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1624635492
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_60
timestamp 1624635492
transform 1 0 6624 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_73
timestamp 1624635492
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1624635492
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9568 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1624635492
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_108
timestamp 1624635492
transform 1 0 11040 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1624635492
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1624635492
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1624635492
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1624635492
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1624635492
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform 1 0 2668 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1624635492
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_20
timestamp 1624635492
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4324 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_25
timestamp 1624635492
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1624635492
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1624635492
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_55
timestamp 1624635492
transform 1 0 6164 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8372 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_79
timestamp 1624635492
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11408 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1624635492
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_112
timestamp 1624635492
transform 1 0 11408 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_124
timestamp 1624635492
transform 1 0 12512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_136
timestamp 1624635492
transform 1 0 13616 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1624635492
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1624635492
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1624635492
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1624635492
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_213
timestamp 1624635492
transform 1 0 20700 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2852 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1624635492
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1624635492
transform 1 0 2392 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_18
timestamp 1624635492
transform 1 0 2760 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform 1 0 3864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6164 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 1624635492
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1624635492
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp 1624635492
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1624635492
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7176 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8740 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_64
timestamp 1624635492
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_75
timestamp 1624635492
transform 1 0 8004 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9752 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1624635492
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_103
timestamp 1624635492
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_107
timestamp 1624635492
transform 1 0 10948 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1624635492
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1624635492
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1624635492
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1624635492
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1624635492
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1624635492
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1624635492
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1624635492
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1624635492
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform 1 0 2576 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1624635492
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_14
timestamp 1624635492
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1624635492
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4140 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1624635492
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624635492
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8004 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5152 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_42
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1624635492
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1624635492
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1624635492
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_79
timestamp 1624635492
transform 1 0 8372 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10764 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624635492
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12236 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_105
timestamp 1624635492
transform 1 0 10764 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1624635492
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1624635492
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_133
timestamp 1624635492
transform 1 0 13340 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1624635492
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1624635492
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1624635492
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1624635492
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1624635492
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1624635492
transform 1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2944 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 1932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1624635492
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1624635492
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1624635492
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1624635492
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1624635492
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 5060 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_46
timestamp 1624635492
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1624635492
transform 1 0 5704 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1624635492
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 7636 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1624635492
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_74
timestamp 1624635492
transform 1 0 7912 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_78
timestamp 1624635492
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_88
timestamp 1624635492
transform 1 0 9200 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_100
timestamp 1624635492
transform 1 0 10304 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform -1 0 12144 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1624635492
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_120
timestamp 1624635492
transform 1 0 12144 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_132
timestamp 1624635492
transform 1 0 13248 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1624635492
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1624635492
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1624635492
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1624635492
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1624635492
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1624635492
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1624635492
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1624635492
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1624635492
transform 1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp 1624635492
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1624635492
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_16
timestamp 1624635492
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5520 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4324 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624635492
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1624635492
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1624635492
transform 1 0 3772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5980 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7452 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_48
timestamp 1624635492
transform 1 0 5520 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_52
timestamp 1624635492
transform 1 0 5888 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_55
timestamp 1624635492
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform -1 0 8464 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9200 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_26_69
timestamp 1624635492
transform 1 0 7452 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_80
timestamp 1624635492
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp 1624635492
transform 1 0 7452 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9384 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10580 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10396 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1624635492
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1624635492
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1624635492
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12236 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1624635492
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_111
timestamp 1624635492
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_137
timestamp 1624635492
transform 1 0 13708 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_126
timestamp 1624635492
transform 1 0 12696 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_138
timestamp 1624635492
transform 1 0 13800 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1624635492
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_150
timestamp 1624635492
transform 1 0 14904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_162
timestamp 1624635492
transform 1 0 16008 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1624635492
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1624635492
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_170
timestamp 1624635492
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1624635492
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1624635492
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1624635492
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1624635492
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1624635492
transform 1 0 20700 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1624635492
transform 1 0 20976 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2852 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 1932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1624635492
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_14
timestamp 1624635492
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_19
timestamp 1624635492
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1624635492
transform 1 0 3312 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_28
timestamp 1624635492
transform 1 0 3680 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5244 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_42
timestamp 1624635492
transform 1 0 4968 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_61
timestamp 1624635492
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6900 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7912 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1624635492
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_83
timestamp 1624635492
transform 1 0 8740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9568 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1624635492
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1624635492
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_113
timestamp 1624635492
transform 1 0 11500 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_125
timestamp 1624635492
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_137
timestamp 1624635492
transform 1 0 13708 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1624635492
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1624635492
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1624635492
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1624635492
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_213
timestamp 1624635492
transform 1 0 20700 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 1932 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1624635492
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_20
timestamp 1624635492
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_25
timestamp 1624635492
transform 1 0 3404 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_37
timestamp 1624635492
transform 1 0 4508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform -1 0 6164 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_49
timestamp 1624635492
transform 1 0 5612 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_55
timestamp 1624635492
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1624635492
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_82
timestamp 1624635492
transform 1 0 8648 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9568 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1624635492
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_101
timestamp 1624635492
transform 1 0 10396 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1624635492
transform 1 0 11500 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1624635492
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1624635492
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1624635492
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1624635492
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1624635492
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1624635492
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1624635492
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform 1 0 2116 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform 1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 1932 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1624635492
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1624635492
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1624635492
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1624635492
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1624635492
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1624635492
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_40
timestamp 1624635492
transform 1 0 4784 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_52
timestamp 1624635492
transform 1 0 5888 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_64
timestamp 1624635492
transform 1 0 6992 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1624635492
transform 1 0 8096 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp 1624635492
transform -1 0 10856 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1624635492
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1624635492
transform 1 0 10212 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1624635492
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_118
timestamp 1624635492
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_130
timestamp 1624635492
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1624635492
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1624635492
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1624635492
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1624635492
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_213
timestamp 1624635492
transform 1 0 20700 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 2392 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1624635492
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1624635492
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1624635492
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 3312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_24
timestamp 1624635492
transform 1 0 3312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1624635492
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1624635492
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_53
timestamp 1624635492
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1624635492
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1624635492
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1624635492
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1624635492
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1624635492
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1624635492
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1624635492
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1624635492
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1624635492
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1624635492
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1624635492
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_220
timestamp 1624635492
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_9
timestamp 1624635492
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1624635492
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_20
timestamp 1624635492
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1624635492
transform 1 0 3312 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_28
timestamp 1624635492
transform 1 0 3680 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1624635492
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1624635492
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1624635492
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1624635492
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1624635492
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1624635492
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1624635492
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1624635492
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1624635492
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1624635492
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1624635492
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_213
timestamp 1624635492
transform 1 0 20700 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1624635492
transform 1 0 1564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1624635492
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 4416 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1624635492
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1624635492
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_36
timestamp 1624635492
transform 1 0 4416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1624635492
transform 1 0 5520 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_56
timestamp 1624635492
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_59
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_71
timestamp 1624635492
transform 1 0 7636 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_83
timestamp 1624635492
transform 1 0 8740 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1624635492
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1624635492
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1624635492
transform 1 0 12972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_146
timestamp 1624635492
transform 1 0 14536 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_158
timestamp 1624635492
transform 1 0 15640 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_170
timestamp 1624635492
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1624635492
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1624635492
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_216
timestamp 1624635492
transform 1 0 20976 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1624635492
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 bottom_right_grid_pin_1_
port 10 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 11 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 12 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 13 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 14 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 15 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 16 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 17 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 18 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 19 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 20 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 21 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 22 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 24 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 25 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 26 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 27 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 28 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 29 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 30 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 31 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 32 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 33 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 34 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 35 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 36 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 37 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 38 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 39 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 40 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 41 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 42 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 43 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 44 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 45 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 46 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 47 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 48 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 49 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 50 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 51 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 52 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[0]
port 53 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[10]
port 54 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[11]
port 55 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[12]
port 56 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[13]
port 57 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[14]
port 58 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[15]
port 59 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[16]
port 60 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[17]
port 61 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_in[18]
port 62 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[19]
port 63 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[1]
port 64 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[2]
port 65 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[3]
port 66 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[4]
port 67 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[5]
port 68 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[6]
port 69 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[7]
port 70 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[8]
port 71 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[9]
port 72 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[0]
port 73 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[10]
port 74 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[11]
port 75 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[12]
port 76 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 chany_bottom_out[13]
port 77 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 chany_bottom_out[14]
port 78 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[15]
port 79 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 chany_bottom_out[16]
port 80 nsew signal tristate
rlabel metal2 s 20074 0 20130 800 6 chany_bottom_out[17]
port 81 nsew signal tristate
rlabel metal2 s 20534 0 20590 800 6 chany_bottom_out[18]
port 82 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[19]
port 83 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_out[1]
port 84 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_out[2]
port 85 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_out[3]
port 86 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 87 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[5]
port 88 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 89 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 90 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[8]
port 91 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 92 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 93 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 94 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 95 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 96 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 97 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 98 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 99 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 100 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 101 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 102 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 103 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 104 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 105 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 106 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 107 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
