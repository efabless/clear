magic
tech sky130A
magscale 1 2
timestamp 1656242771
<< viali >>
rect 3157 20553 3191 20587
rect 3985 20553 4019 20587
rect 4629 20553 4663 20587
rect 9689 20553 9723 20587
rect 10701 20553 10735 20587
rect 13369 20553 13403 20587
rect 14289 20553 14323 20587
rect 15393 20553 15427 20587
rect 16865 20553 16899 20587
rect 17969 20553 18003 20587
rect 2237 20417 2271 20451
rect 2789 20417 2823 20451
rect 3341 20417 3375 20451
rect 3801 20417 3835 20451
rect 4445 20417 4479 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 5825 20417 5859 20451
rect 6745 20417 6779 20451
rect 7481 20417 7515 20451
rect 7941 20417 7975 20451
rect 8401 20417 8435 20451
rect 9045 20417 9079 20451
rect 9505 20417 9539 20451
rect 10057 20417 10091 20451
rect 10517 20417 10551 20451
rect 11161 20417 11195 20451
rect 11805 20417 11839 20451
rect 12449 20417 12483 20451
rect 12909 20417 12943 20451
rect 13185 20417 13219 20451
rect 14105 20417 14139 20451
rect 14657 20417 14691 20451
rect 15209 20417 15243 20451
rect 15761 20417 15795 20451
rect 16681 20417 16715 20451
rect 17233 20417 17267 20451
rect 17785 20417 17819 20451
rect 18337 20417 18371 20451
rect 20545 20417 20579 20451
rect 1961 20349 1995 20383
rect 6837 20349 6871 20383
rect 7021 20349 7055 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 21189 20349 21223 20383
rect 6377 20281 6411 20315
rect 14841 20281 14875 20315
rect 15945 20281 15979 20315
rect 17417 20281 17451 20315
rect 2605 20213 2639 20247
rect 5089 20213 5123 20247
rect 5549 20213 5583 20247
rect 6009 20213 6043 20247
rect 7665 20213 7699 20247
rect 8125 20213 8159 20247
rect 8585 20213 8619 20247
rect 9229 20213 9263 20247
rect 10241 20213 10275 20247
rect 10977 20213 11011 20247
rect 11989 20213 12023 20247
rect 12265 20213 12299 20247
rect 12725 20213 12759 20247
rect 18521 20213 18555 20247
rect 10609 20009 10643 20043
rect 10977 20009 11011 20043
rect 11713 20009 11747 20043
rect 12173 20009 12207 20043
rect 12633 20009 12667 20043
rect 12909 20009 12943 20043
rect 15669 20009 15703 20043
rect 16313 20009 16347 20043
rect 19441 20009 19475 20043
rect 6101 19941 6135 19975
rect 9229 19941 9263 19975
rect 9689 19941 9723 19975
rect 10149 19941 10183 19975
rect 5549 19873 5583 19907
rect 6469 19873 6503 19907
rect 8125 19873 8159 19907
rect 18613 19873 18647 19907
rect 21373 19873 21407 19907
rect 1961 19805 1995 19839
rect 2237 19805 2271 19839
rect 2513 19805 2547 19839
rect 3249 19805 3283 19839
rect 4169 19805 4203 19839
rect 4445 19805 4479 19839
rect 4905 19805 4939 19839
rect 8033 19805 8067 19839
rect 9045 19805 9079 19839
rect 9505 19805 9539 19839
rect 9965 19805 9999 19839
rect 10425 19805 10459 19839
rect 11253 19805 11287 19839
rect 15485 19805 15519 19839
rect 16129 19805 16163 19839
rect 16681 19805 16715 19839
rect 19257 19805 19291 19839
rect 5641 19737 5675 19771
rect 5733 19737 5767 19771
rect 13369 19737 13403 19771
rect 13737 19737 13771 19771
rect 14197 19737 14231 19771
rect 14565 19737 14599 19771
rect 18346 19737 18380 19771
rect 21128 19737 21162 19771
rect 2697 19669 2731 19703
rect 3433 19669 3467 19703
rect 3985 19669 4019 19703
rect 4629 19669 4663 19703
rect 5089 19669 5123 19703
rect 6653 19669 6687 19703
rect 6745 19669 6779 19703
rect 7113 19669 7147 19703
rect 7573 19669 7607 19703
rect 7941 19669 7975 19703
rect 11437 19669 11471 19703
rect 15209 19669 15243 19703
rect 16865 19669 16899 19703
rect 17233 19669 17267 19703
rect 19993 19669 20027 19703
rect 2513 19465 2547 19499
rect 3617 19465 3651 19499
rect 6837 19465 6871 19499
rect 7481 19465 7515 19499
rect 8677 19465 8711 19499
rect 9137 19465 9171 19499
rect 9597 19465 9631 19499
rect 10057 19465 10091 19499
rect 10517 19465 10551 19499
rect 10793 19465 10827 19499
rect 14105 19465 14139 19499
rect 18061 19465 18095 19499
rect 19073 19465 19107 19499
rect 7389 19397 7423 19431
rect 1685 19329 1719 19363
rect 1961 19329 1995 19363
rect 2697 19329 2731 19363
rect 2973 19329 3007 19363
rect 3433 19329 3467 19363
rect 4169 19329 4203 19363
rect 4813 19329 4847 19363
rect 5549 19329 5583 19363
rect 5825 19329 5859 19363
rect 6653 19329 6687 19363
rect 8493 19329 8527 19363
rect 8953 19329 8987 19363
rect 9413 19329 9447 19363
rect 9873 19329 9907 19363
rect 10333 19329 10367 19363
rect 13562 19329 13596 19363
rect 13829 19329 13863 19363
rect 15218 19329 15252 19363
rect 16937 19329 16971 19363
rect 18337 19329 18371 19363
rect 18889 19329 18923 19363
rect 20830 19329 20864 19363
rect 21097 19329 21131 19363
rect 7297 19261 7331 19295
rect 8217 19261 8251 19295
rect 11621 19261 11655 19295
rect 15485 19261 15519 19295
rect 16681 19261 16715 19295
rect 2145 19193 2179 19227
rect 4629 19193 4663 19227
rect 6009 19193 6043 19227
rect 18521 19193 18555 19227
rect 1501 19125 1535 19159
rect 3157 19125 3191 19159
rect 4353 19125 4387 19159
rect 5365 19125 5399 19159
rect 7849 19125 7883 19159
rect 11989 19125 12023 19159
rect 12449 19125 12483 19159
rect 15761 19125 15795 19159
rect 16129 19125 16163 19159
rect 19717 19125 19751 19159
rect 2513 18921 2547 18955
rect 3801 18921 3835 18955
rect 5365 18921 5399 18955
rect 7389 18921 7423 18955
rect 9781 18921 9815 18955
rect 10333 18921 10367 18955
rect 18797 18921 18831 18955
rect 21097 18921 21131 18955
rect 2145 18853 2179 18887
rect 7849 18853 7883 18887
rect 11069 18853 11103 18887
rect 6193 18785 6227 18819
rect 6837 18785 6871 18819
rect 8493 18785 8527 18819
rect 13737 18785 13771 18819
rect 17509 18785 17543 18819
rect 1685 18717 1719 18751
rect 1961 18717 1995 18751
rect 2697 18717 2731 18751
rect 3065 18717 3099 18751
rect 3985 18717 4019 18751
rect 4445 18717 4479 18751
rect 4905 18717 4939 18751
rect 5181 18717 5215 18751
rect 5733 18717 5767 18751
rect 9045 18717 9079 18751
rect 9965 18717 9999 18751
rect 10701 18717 10735 18751
rect 11437 18717 11471 18751
rect 15485 18717 15519 18751
rect 15761 18717 15795 18751
rect 18061 18717 18095 18751
rect 18613 18717 18647 18751
rect 19257 18717 19291 18751
rect 20913 18717 20947 18751
rect 6929 18649 6963 18683
rect 8309 18649 8343 18683
rect 13470 18649 13504 18683
rect 15218 18649 15252 18683
rect 17242 18649 17276 18683
rect 19524 18649 19558 18683
rect 1501 18581 1535 18615
rect 3249 18581 3283 18615
rect 4261 18581 4295 18615
rect 4721 18581 4755 18615
rect 7021 18581 7055 18615
rect 8217 18581 8251 18615
rect 9229 18581 9263 18615
rect 11989 18581 12023 18615
rect 12357 18581 12391 18615
rect 14105 18581 14139 18615
rect 16129 18581 16163 18615
rect 18245 18581 18279 18615
rect 20637 18581 20671 18615
rect 1961 18377 1995 18411
rect 2605 18377 2639 18411
rect 3525 18377 3559 18411
rect 5641 18377 5675 18411
rect 7573 18377 7607 18411
rect 8033 18377 8067 18411
rect 8309 18377 8343 18411
rect 9597 18377 9631 18411
rect 16681 18377 16715 18411
rect 21373 18377 21407 18411
rect 7665 18309 7699 18343
rect 10885 18309 10919 18343
rect 12992 18309 13026 18343
rect 15516 18309 15550 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2421 18241 2455 18275
rect 2881 18241 2915 18275
rect 3341 18241 3375 18275
rect 4077 18241 4111 18275
rect 5181 18241 5215 18275
rect 5457 18241 5491 18275
rect 8769 18241 8803 18275
rect 9413 18241 9447 18275
rect 10793 18241 10827 18275
rect 11529 18241 11563 18275
rect 15761 18241 15795 18275
rect 17794 18241 17828 18275
rect 19450 18241 19484 18275
rect 19717 18241 19751 18275
rect 19993 18241 20027 18275
rect 20249 18241 20283 18275
rect 4537 18173 4571 18207
rect 7481 18173 7515 18207
rect 9965 18173 9999 18207
rect 10977 18173 11011 18207
rect 12725 18173 12759 18207
rect 18061 18173 18095 18207
rect 3893 18105 3927 18139
rect 5917 18105 5951 18139
rect 8953 18105 8987 18139
rect 14381 18105 14415 18139
rect 16037 18105 16071 18139
rect 1501 18037 1535 18071
rect 3065 18037 3099 18071
rect 4997 18037 5031 18071
rect 6377 18037 6411 18071
rect 6837 18037 6871 18071
rect 10425 18037 10459 18071
rect 11989 18037 12023 18071
rect 12449 18037 12483 18071
rect 14105 18037 14139 18071
rect 18337 18037 18371 18071
rect 2513 17833 2547 17867
rect 4077 17833 4111 17867
rect 5457 17833 5491 17867
rect 10793 17833 10827 17867
rect 12081 17833 12115 17867
rect 17877 17833 17911 17867
rect 18245 17833 18279 17867
rect 18889 17833 18923 17867
rect 11069 17765 11103 17799
rect 19625 17765 19659 17799
rect 4721 17697 4755 17731
rect 6101 17697 6135 17731
rect 8033 17697 8067 17731
rect 9597 17697 9631 17731
rect 10057 17697 10091 17731
rect 1685 17629 1719 17663
rect 1961 17629 1995 17663
rect 2697 17629 2731 17663
rect 4445 17629 4479 17663
rect 9413 17629 9447 17663
rect 10609 17629 10643 17663
rect 13737 17629 13771 17663
rect 15485 17629 15519 17663
rect 15853 17629 15887 17663
rect 16129 17629 16163 17663
rect 19441 17629 19475 17663
rect 21373 17629 21407 17663
rect 5825 17561 5859 17595
rect 6469 17561 6503 17595
rect 8217 17561 8251 17595
rect 13470 17561 13504 17595
rect 15218 17561 15252 17595
rect 16374 17561 16408 17595
rect 21106 17561 21140 17595
rect 1501 17493 1535 17527
rect 2145 17493 2179 17527
rect 3433 17493 3467 17527
rect 4537 17493 4571 17527
rect 5089 17493 5123 17527
rect 5917 17493 5951 17527
rect 7205 17493 7239 17527
rect 8125 17493 8159 17527
rect 8585 17493 8619 17527
rect 8953 17493 8987 17527
rect 9321 17493 9355 17527
rect 11713 17493 11747 17527
rect 12357 17493 12391 17527
rect 14105 17493 14139 17527
rect 17509 17493 17543 17527
rect 19993 17493 20027 17527
rect 1961 17289 1995 17323
rect 2789 17289 2823 17323
rect 3249 17289 3283 17323
rect 3617 17289 3651 17323
rect 4537 17289 4571 17323
rect 4997 17289 5031 17323
rect 6377 17289 6411 17323
rect 6837 17289 6871 17323
rect 7573 17289 7607 17323
rect 8033 17289 8067 17323
rect 9137 17289 9171 17323
rect 9873 17289 9907 17323
rect 11069 17289 11103 17323
rect 11621 17289 11655 17323
rect 11989 17289 12023 17323
rect 14013 17289 14047 17323
rect 14381 17289 14415 17323
rect 14749 17289 14783 17323
rect 19349 17289 19383 17323
rect 2513 17221 2547 17255
rect 7941 17221 7975 17255
rect 9413 17221 9447 17255
rect 13378 17221 13412 17255
rect 17325 17221 17359 17255
rect 21106 17221 21140 17255
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2973 17153 3007 17187
rect 4905 17153 4939 17187
rect 5825 17153 5859 17187
rect 6745 17153 6779 17187
rect 8953 17153 8987 17187
rect 10333 17153 10367 17187
rect 13638 17153 13672 17187
rect 17601 17153 17635 17187
rect 17868 17153 17902 17187
rect 21373 17153 21407 17187
rect 3709 17085 3743 17119
rect 3801 17085 3835 17119
rect 5181 17085 5215 17119
rect 7021 17085 7055 17119
rect 8217 17085 8251 17119
rect 8677 17085 8711 17119
rect 6009 17017 6043 17051
rect 10609 17017 10643 17051
rect 12265 17017 12299 17051
rect 1501 16949 1535 16983
rect 15301 16949 15335 16983
rect 15669 16949 15703 16983
rect 16313 16949 16347 16983
rect 16957 16949 16991 16983
rect 18981 16949 19015 16983
rect 19717 16949 19751 16983
rect 19993 16949 20027 16983
rect 2421 16745 2455 16779
rect 3249 16745 3283 16779
rect 4169 16745 4203 16779
rect 2973 16677 3007 16711
rect 12081 16677 12115 16711
rect 4629 16609 4663 16643
rect 4813 16609 4847 16643
rect 7205 16609 7239 16643
rect 7941 16609 7975 16643
rect 8953 16609 8987 16643
rect 10977 16609 11011 16643
rect 11069 16609 11103 16643
rect 12357 16609 12391 16643
rect 15761 16609 15795 16643
rect 18889 16609 18923 16643
rect 19441 16609 19475 16643
rect 1685 16541 1719 16575
rect 2145 16541 2179 16575
rect 2605 16541 2639 16575
rect 3433 16541 3467 16575
rect 8217 16541 8251 16575
rect 9781 16541 9815 16575
rect 10057 16541 10091 16575
rect 14105 16541 14139 16575
rect 19697 16541 19731 16575
rect 21097 16541 21131 16575
rect 4537 16473 4571 16507
rect 5181 16473 5215 16507
rect 6285 16473 6319 16507
rect 6929 16473 6963 16507
rect 12602 16473 12636 16507
rect 14350 16473 14384 16507
rect 16028 16473 16062 16507
rect 18622 16473 18656 16507
rect 1501 16405 1535 16439
rect 1961 16405 1995 16439
rect 3893 16405 3927 16439
rect 5733 16405 5767 16439
rect 6561 16405 6595 16439
rect 7021 16405 7055 16439
rect 8125 16405 8159 16439
rect 8585 16405 8619 16439
rect 9597 16405 9631 16439
rect 10241 16405 10275 16439
rect 10517 16405 10551 16439
rect 10885 16405 10919 16439
rect 11713 16405 11747 16439
rect 13737 16405 13771 16439
rect 15485 16405 15519 16439
rect 17141 16405 17175 16439
rect 17509 16405 17543 16439
rect 20821 16405 20855 16439
rect 21281 16405 21315 16439
rect 2789 16201 2823 16235
rect 3341 16201 3375 16235
rect 3801 16201 3835 16235
rect 5549 16201 5583 16235
rect 6377 16201 6411 16235
rect 7389 16201 7423 16235
rect 7941 16201 7975 16235
rect 8309 16201 8343 16235
rect 9045 16201 9079 16235
rect 10149 16201 10183 16235
rect 10885 16201 10919 16235
rect 11897 16201 11931 16235
rect 15301 16201 15335 16235
rect 16313 16201 16347 16235
rect 20729 16201 20763 16235
rect 14320 16133 14354 16167
rect 19318 16133 19352 16167
rect 1685 16065 1719 16099
rect 2237 16065 2271 16099
rect 2973 16065 3007 16099
rect 3709 16065 3743 16099
rect 4537 16065 4571 16099
rect 5457 16065 5491 16099
rect 6745 16065 6779 16099
rect 7573 16065 7607 16099
rect 8401 16065 8435 16099
rect 9321 16065 9355 16099
rect 10333 16065 10367 16099
rect 12909 16065 12943 16099
rect 14565 16065 14599 16099
rect 17794 16065 17828 16099
rect 18061 16065 18095 16099
rect 18429 16065 18463 16099
rect 19073 16065 19107 16099
rect 3985 15997 4019 16031
rect 5641 15997 5675 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 8585 15997 8619 16031
rect 11989 15997 12023 16031
rect 12173 15997 12207 16031
rect 18705 15997 18739 16031
rect 2053 15929 2087 15963
rect 4353 15929 4387 15963
rect 21189 15929 21223 15963
rect 1501 15861 1535 15895
rect 5089 15861 5123 15895
rect 9689 15861 9723 15895
rect 11529 15861 11563 15895
rect 13185 15861 13219 15895
rect 14841 15861 14875 15895
rect 15577 15861 15611 15895
rect 16681 15861 16715 15895
rect 20453 15861 20487 15895
rect 1961 15657 1995 15691
rect 2881 15657 2915 15691
rect 7389 15657 7423 15691
rect 8585 15657 8619 15691
rect 10241 15657 10275 15691
rect 13001 15657 13035 15691
rect 2421 15589 2455 15623
rect 15485 15589 15519 15623
rect 18521 15589 18555 15623
rect 18889 15589 18923 15623
rect 4813 15521 4847 15555
rect 6285 15521 6319 15555
rect 6837 15521 6871 15555
rect 8033 15521 8067 15555
rect 11253 15521 11287 15555
rect 11437 15521 11471 15555
rect 21373 15521 21407 15555
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 2605 15453 2639 15487
rect 3065 15453 3099 15487
rect 4997 15453 5031 15487
rect 6929 15453 6963 15487
rect 10425 15453 10459 15487
rect 13369 15453 13403 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 15853 15453 15887 15487
rect 16497 15453 16531 15487
rect 16773 15453 16807 15487
rect 4169 15385 4203 15419
rect 4905 15385 4939 15419
rect 6009 15385 6043 15419
rect 8217 15385 8251 15419
rect 8953 15385 8987 15419
rect 9413 15385 9447 15419
rect 11161 15385 11195 15419
rect 11805 15385 11839 15419
rect 14372 15385 14406 15419
rect 17018 15385 17052 15419
rect 21106 15385 21140 15419
rect 1501 15317 1535 15351
rect 3433 15317 3467 15351
rect 5365 15317 5399 15351
rect 5641 15317 5675 15351
rect 6101 15317 6135 15351
rect 7021 15317 7055 15351
rect 8125 15317 8159 15351
rect 9781 15317 9815 15351
rect 10793 15317 10827 15351
rect 18153 15317 18187 15351
rect 19349 15317 19383 15351
rect 19717 15317 19751 15351
rect 19993 15317 20027 15351
rect 1961 15113 1995 15147
rect 2605 15113 2639 15147
rect 2973 15113 3007 15147
rect 3985 15113 4019 15147
rect 5549 15113 5583 15147
rect 6009 15113 6043 15147
rect 7849 15113 7883 15147
rect 10333 15113 10367 15147
rect 10793 15113 10827 15147
rect 14565 15113 14599 15147
rect 4537 15045 4571 15079
rect 8309 15045 8343 15079
rect 16068 15045 16102 15079
rect 18521 15045 18555 15079
rect 19717 15045 19751 15079
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 2421 14977 2455 15011
rect 3617 14977 3651 15011
rect 4629 14977 4663 15011
rect 5641 14977 5675 15011
rect 7205 14977 7239 15011
rect 8217 14977 8251 15011
rect 9229 14977 9263 15011
rect 9873 14977 9907 15011
rect 10517 14977 10551 15011
rect 10977 14977 11011 15011
rect 13452 14977 13486 15011
rect 16313 14977 16347 15011
rect 17978 14977 18012 15011
rect 18245 14977 18279 15011
rect 18889 14977 18923 15011
rect 21106 14977 21140 15011
rect 21373 14977 21407 15011
rect 3433 14909 3467 14943
rect 3525 14909 3559 14943
rect 4445 14909 4479 14943
rect 5365 14909 5399 14943
rect 6929 14909 6963 14943
rect 7113 14909 7147 14943
rect 8401 14909 8435 14943
rect 9321 14909 9355 14943
rect 9505 14909 9539 14943
rect 13185 14909 13219 14943
rect 4997 14841 5031 14875
rect 1501 14773 1535 14807
rect 6377 14773 6411 14807
rect 7573 14773 7607 14807
rect 8861 14773 8895 14807
rect 14933 14773 14967 14807
rect 16865 14773 16899 14807
rect 19349 14773 19383 14807
rect 19993 14773 20027 14807
rect 2513 14569 2547 14603
rect 3985 14569 4019 14603
rect 5365 14569 5399 14603
rect 5825 14569 5859 14603
rect 6561 14569 6595 14603
rect 6837 14569 6871 14603
rect 7297 14569 7331 14603
rect 7665 14569 7699 14603
rect 8309 14569 8343 14603
rect 8953 14569 8987 14603
rect 11253 14569 11287 14603
rect 16221 14569 16255 14603
rect 16589 14569 16623 14603
rect 18245 14569 18279 14603
rect 19349 14569 19383 14603
rect 3433 14501 3467 14535
rect 5089 14501 5123 14535
rect 15853 14501 15887 14535
rect 19901 14501 19935 14535
rect 4445 14433 4479 14467
rect 4629 14433 4663 14467
rect 6193 14433 6227 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 10701 14433 10735 14467
rect 17969 14433 18003 14467
rect 21281 14433 21315 14467
rect 1685 14365 1719 14399
rect 2237 14365 2271 14399
rect 2697 14365 2731 14399
rect 4353 14365 4387 14399
rect 8125 14365 8159 14399
rect 13737 14365 13771 14399
rect 14105 14365 14139 14399
rect 14473 14365 14507 14399
rect 21014 14365 21048 14399
rect 14718 14297 14752 14331
rect 17702 14297 17736 14331
rect 1501 14229 1535 14263
rect 2053 14229 2087 14263
rect 2973 14229 3007 14263
rect 9321 14229 9355 14263
rect 10793 14229 10827 14263
rect 10885 14229 10919 14263
rect 11529 14229 11563 14263
rect 18889 14229 18923 14263
rect 2421 14025 2455 14059
rect 3065 14025 3099 14059
rect 3525 14025 3559 14059
rect 4629 14025 4663 14059
rect 5641 14025 5675 14059
rect 7205 14025 7239 14059
rect 8033 14025 8067 14059
rect 8401 14025 8435 14059
rect 9137 14025 9171 14059
rect 9505 14025 9539 14059
rect 9873 14025 9907 14059
rect 15209 14025 15243 14059
rect 16681 14025 16715 14059
rect 17049 14025 17083 14059
rect 17417 14025 17451 14059
rect 20729 14025 20763 14059
rect 21189 14025 21223 14059
rect 5181 13957 5215 13991
rect 1685 13889 1719 13923
rect 3433 13889 3467 13923
rect 5273 13889 5307 13923
rect 6837 13889 6871 13923
rect 7481 13889 7515 13923
rect 8493 13889 8527 13923
rect 10241 13889 10275 13923
rect 10885 13889 10919 13923
rect 13297 13889 13331 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 14085 13889 14119 13923
rect 15945 13889 15979 13923
rect 18530 13889 18564 13923
rect 18797 13889 18831 13923
rect 20197 13889 20231 13923
rect 20453 13889 20487 13923
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 3709 13821 3743 13855
rect 5089 13821 5123 13855
rect 6009 13821 6043 13855
rect 6653 13821 6687 13855
rect 6745 13821 6779 13855
rect 8677 13821 8711 13855
rect 10333 13821 10367 13855
rect 10517 13821 10551 13855
rect 16313 13821 16347 13855
rect 2789 13753 2823 13787
rect 4077 13753 4111 13787
rect 19073 13753 19107 13787
rect 1501 13685 1535 13719
rect 12173 13685 12207 13719
rect 15577 13685 15611 13719
rect 2697 13481 2731 13515
rect 3985 13481 4019 13515
rect 6377 13481 6411 13515
rect 7849 13481 7883 13515
rect 21189 13481 21223 13515
rect 2421 13413 2455 13447
rect 5825 13413 5859 13447
rect 9045 13413 9079 13447
rect 15485 13413 15519 13447
rect 18889 13413 18923 13447
rect 3157 13345 3191 13379
rect 3341 13345 3375 13379
rect 4537 13345 4571 13379
rect 5273 13345 5307 13379
rect 6929 13345 6963 13379
rect 8401 13345 8435 13379
rect 11345 13345 11379 13379
rect 11529 13345 11563 13379
rect 15853 13345 15887 13379
rect 16405 13345 16439 13379
rect 16865 13345 16899 13379
rect 17233 13345 17267 13379
rect 17509 13345 17543 13379
rect 20913 13345 20947 13379
rect 1409 13277 1443 13311
rect 1869 13277 1903 13311
rect 3065 13277 3099 13311
rect 5365 13277 5399 13311
rect 12173 13277 12207 13311
rect 14105 13277 14139 13311
rect 17765 13277 17799 13311
rect 21373 13277 21407 13311
rect 4445 13209 4479 13243
rect 5457 13209 5491 13243
rect 6745 13209 6779 13243
rect 7389 13209 7423 13243
rect 8309 13209 8343 13243
rect 10517 13209 10551 13243
rect 11253 13209 11287 13243
rect 12418 13209 12452 13243
rect 14372 13209 14406 13243
rect 20668 13209 20702 13243
rect 1593 13141 1627 13175
rect 4353 13141 4387 13175
rect 6837 13141 6871 13175
rect 8217 13141 8251 13175
rect 10885 13141 10919 13175
rect 13553 13141 13587 13175
rect 19533 13141 19567 13175
rect 1961 12937 1995 12971
rect 3065 12937 3099 12971
rect 5273 12937 5307 12971
rect 5733 12937 5767 12971
rect 7113 12937 7147 12971
rect 8125 12937 8159 12971
rect 8677 12937 8711 12971
rect 9137 12937 9171 12971
rect 11529 12937 11563 12971
rect 12817 12937 12851 12971
rect 16681 12937 16715 12971
rect 18429 12937 18463 12971
rect 18981 12937 19015 12971
rect 19349 12937 19383 12971
rect 19809 12937 19843 12971
rect 6653 12869 6687 12903
rect 9689 12869 9723 12903
rect 14228 12869 14262 12903
rect 1777 12801 1811 12835
rect 2237 12801 2271 12835
rect 2697 12801 2731 12835
rect 5365 12801 5399 12835
rect 6745 12801 6779 12835
rect 8033 12801 8067 12835
rect 9045 12801 9079 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 14473 12801 14507 12835
rect 17794 12801 17828 12835
rect 18061 12801 18095 12835
rect 20922 12801 20956 12835
rect 21189 12801 21223 12835
rect 3525 12733 3559 12767
rect 4353 12733 4387 12767
rect 5181 12733 5215 12767
rect 6561 12733 6595 12767
rect 8217 12733 8251 12767
rect 9321 12733 9355 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 1409 12665 1443 12699
rect 2421 12665 2455 12699
rect 3985 12597 4019 12631
rect 7665 12597 7699 12631
rect 13093 12597 13127 12631
rect 14841 12597 14875 12631
rect 2145 12393 2179 12427
rect 3433 12393 3467 12427
rect 4537 12393 4571 12427
rect 9689 12393 9723 12427
rect 12081 12393 12115 12427
rect 18889 12393 18923 12427
rect 19257 12393 19291 12427
rect 5549 12325 5583 12359
rect 7297 12325 7331 12359
rect 14565 12325 14599 12359
rect 16773 12325 16807 12359
rect 2789 12257 2823 12291
rect 2973 12257 3007 12291
rect 3893 12257 3927 12291
rect 4077 12257 4111 12291
rect 4997 12257 5031 12291
rect 5089 12257 5123 12291
rect 6285 12257 6319 12291
rect 6745 12257 6779 12291
rect 8401 12257 8435 12291
rect 9137 12257 9171 12291
rect 11529 12257 11563 12291
rect 17141 12257 17175 12291
rect 21373 12257 21407 12291
rect 1409 12189 1443 12223
rect 2329 12189 2363 12223
rect 3065 12189 3099 12223
rect 4169 12189 4203 12223
rect 11621 12189 11655 12223
rect 13481 12189 13515 12223
rect 13737 12189 13771 12223
rect 14197 12189 14231 12223
rect 15025 12189 15059 12223
rect 6837 12121 6871 12155
rect 9321 12121 9355 12155
rect 9965 12121 9999 12155
rect 15292 12121 15326 12155
rect 17386 12121 17420 12155
rect 21106 12121 21140 12155
rect 1593 12053 1627 12087
rect 5181 12053 5215 12087
rect 6929 12053 6963 12087
rect 9229 12053 9263 12087
rect 11069 12053 11103 12087
rect 11713 12053 11747 12087
rect 12357 12053 12391 12087
rect 16405 12053 16439 12087
rect 18521 12053 18555 12087
rect 19625 12053 19659 12087
rect 19993 12053 20027 12087
rect 1961 11849 1995 11883
rect 2789 11849 2823 11883
rect 4261 11849 4295 11883
rect 6377 11849 6411 11883
rect 10425 11849 10459 11883
rect 10885 11849 10919 11883
rect 13829 11849 13863 11883
rect 14197 11849 14231 11883
rect 15945 11849 15979 11883
rect 17693 11849 17727 11883
rect 19625 11849 19659 11883
rect 21281 11849 21315 11883
rect 20738 11781 20772 11815
rect 1409 11713 1443 11747
rect 2145 11713 2179 11747
rect 4721 11713 4755 11747
rect 5365 11713 5399 11747
rect 6561 11713 6595 11747
rect 10057 11713 10091 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 13205 11713 13239 11747
rect 13461 11713 13495 11747
rect 14821 11713 14855 11747
rect 16313 11713 16347 11747
rect 16681 11713 16715 11747
rect 17233 11713 17267 11747
rect 18806 11713 18840 11747
rect 19073 11713 19107 11747
rect 21005 11713 21039 11747
rect 2421 11645 2455 11679
rect 3617 11645 3651 11679
rect 5457 11645 5491 11679
rect 5549 11645 5583 11679
rect 11069 11645 11103 11679
rect 14565 11645 14599 11679
rect 1593 11577 1627 11611
rect 3157 11509 3191 11543
rect 4997 11509 5031 11543
rect 12081 11509 12115 11543
rect 1961 11305 1995 11339
rect 2605 11305 2639 11339
rect 3801 11305 3835 11339
rect 5549 11305 5583 11339
rect 6745 11305 6779 11339
rect 8953 11305 8987 11339
rect 15485 11305 15519 11339
rect 17417 11305 17451 11339
rect 21005 11305 21039 11339
rect 21373 11305 21407 11339
rect 1593 11237 1627 11271
rect 12357 11237 12391 11271
rect 15761 11237 15795 11271
rect 4905 11169 4939 11203
rect 6193 11169 6227 11203
rect 9505 11169 9539 11203
rect 10701 11169 10735 11203
rect 10885 11169 10919 11203
rect 17141 11169 17175 11203
rect 18797 11169 18831 11203
rect 1409 11101 1443 11135
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2881 11101 2915 11135
rect 3985 11101 4019 11135
rect 6285 11101 6319 11135
rect 7021 11101 7055 11135
rect 9413 11101 9447 11135
rect 10609 11101 10643 11135
rect 13481 11101 13515 11135
rect 13737 11101 13771 11135
rect 14105 11101 14139 11135
rect 19625 11101 19659 11135
rect 19881 11101 19915 11135
rect 5089 11033 5123 11067
rect 5181 11033 5215 11067
rect 6377 11033 6411 11067
rect 8585 11033 8619 11067
rect 9321 11033 9355 11067
rect 14350 11033 14384 11067
rect 16874 11033 16908 11067
rect 18530 11033 18564 11067
rect 19257 11033 19291 11067
rect 10241 10965 10275 10999
rect 2513 10761 2547 10795
rect 3157 10761 3191 10795
rect 3617 10761 3651 10795
rect 5365 10761 5399 10795
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 7757 10761 7791 10795
rect 9873 10761 9907 10795
rect 10333 10761 10367 10795
rect 13001 10761 13035 10795
rect 14657 10761 14691 10795
rect 18337 10761 18371 10795
rect 19993 10761 20027 10795
rect 8769 10693 8803 10727
rect 12725 10693 12759 10727
rect 16948 10693 16982 10727
rect 19450 10693 19484 10727
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 3341 10625 3375 10659
rect 3801 10625 3835 10659
rect 5549 10625 5583 10659
rect 6009 10625 6043 10659
rect 7849 10625 7883 10659
rect 10241 10625 10275 10659
rect 10885 10625 10919 10659
rect 14114 10625 14148 10659
rect 14381 10625 14415 10659
rect 15770 10625 15804 10659
rect 16037 10625 16071 10659
rect 16681 10625 16715 10659
rect 19717 10625 19751 10659
rect 21106 10625 21140 10659
rect 21373 10625 21407 10659
rect 2237 10557 2271 10591
rect 6561 10557 6595 10591
rect 6653 10557 6687 10591
rect 8033 10557 8067 10591
rect 9321 10557 9355 10591
rect 10517 10557 10551 10591
rect 1593 10489 1627 10523
rect 7389 10489 7423 10523
rect 5825 10421 5859 10455
rect 18061 10421 18095 10455
rect 1961 10217 1995 10251
rect 4169 10217 4203 10251
rect 5733 10217 5767 10251
rect 6837 10217 6871 10251
rect 7849 10217 7883 10251
rect 9689 10217 9723 10251
rect 10701 10217 10735 10251
rect 14105 10217 14139 10251
rect 19349 10217 19383 10251
rect 21373 10217 21407 10251
rect 2421 10149 2455 10183
rect 12357 10149 12391 10183
rect 2789 10081 2823 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 5273 10081 5307 10115
rect 7297 10081 7331 10115
rect 7481 10081 7515 10115
rect 8493 10081 8527 10115
rect 9137 10081 9171 10115
rect 13737 10081 13771 10115
rect 1409 10013 1443 10047
rect 2145 10013 2179 10047
rect 7205 10013 7239 10047
rect 9321 10013 9355 10047
rect 13470 10013 13504 10047
rect 15229 10013 15263 10047
rect 15485 10013 15519 10047
rect 16874 10013 16908 10047
rect 17141 10013 17175 10047
rect 17417 10013 17451 10047
rect 17673 10013 17707 10047
rect 19993 10013 20027 10047
rect 4537 9945 4571 9979
rect 20238 9945 20272 9979
rect 1593 9877 1627 9911
rect 6561 9877 6595 9911
rect 8217 9877 8251 9911
rect 8309 9877 8343 9911
rect 9229 9877 9263 9911
rect 10333 9877 10367 9911
rect 15761 9877 15795 9911
rect 18797 9877 18831 9911
rect 1593 9673 1627 9707
rect 6745 9673 6779 9707
rect 9413 9673 9447 9707
rect 9781 9673 9815 9707
rect 10425 9673 10459 9707
rect 10793 9673 10827 9707
rect 10885 9673 10919 9707
rect 17049 9673 17083 9707
rect 20269 9673 20303 9707
rect 21005 9673 21039 9707
rect 21373 9673 21407 9707
rect 7113 9605 7147 9639
rect 7205 9605 7239 9639
rect 9873 9605 9907 9639
rect 14718 9605 14752 9639
rect 16221 9605 16255 9639
rect 16773 9605 16807 9639
rect 17509 9605 17543 9639
rect 18245 9605 18279 9639
rect 18981 9605 19015 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 4721 9537 4755 9571
rect 5917 9537 5951 9571
rect 8769 9537 8803 9571
rect 13286 9537 13320 9571
rect 13553 9537 13587 9571
rect 13921 9537 13955 9571
rect 14473 9537 14507 9571
rect 19809 9537 19843 9571
rect 7297 9469 7331 9503
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 10057 9469 10091 9503
rect 10977 9469 11011 9503
rect 19533 9469 19567 9503
rect 2237 9401 2271 9435
rect 5733 9401 5767 9435
rect 8401 9401 8435 9435
rect 12173 9401 12207 9435
rect 15853 9401 15887 9435
rect 20545 9401 20579 9435
rect 4537 9333 4571 9367
rect 6469 9333 6503 9367
rect 7849 9333 7883 9367
rect 11529 9333 11563 9367
rect 18613 9333 18647 9367
rect 2053 9129 2087 9163
rect 4537 9129 4571 9163
rect 7297 9129 7331 9163
rect 9597 9129 9631 9163
rect 10609 9129 10643 9163
rect 13737 9129 13771 9163
rect 16037 9129 16071 9163
rect 19349 9129 19383 9163
rect 20453 9129 20487 9163
rect 20821 9129 20855 9163
rect 21189 9129 21223 9163
rect 2513 9061 2547 9095
rect 19809 9061 19843 9095
rect 2881 8993 2915 9027
rect 5181 8993 5215 9027
rect 6193 8993 6227 9027
rect 10241 8993 10275 9027
rect 11253 8993 11287 9027
rect 12081 8993 12115 9027
rect 12265 8993 12299 9027
rect 1409 8925 1443 8959
rect 2237 8925 2271 8959
rect 4997 8925 5031 8959
rect 4905 8857 4939 8891
rect 5917 8857 5951 8891
rect 6561 8857 6595 8891
rect 9321 8857 9355 8891
rect 9965 8857 9999 8891
rect 10977 8857 11011 8891
rect 1593 8789 1627 8823
rect 5549 8789 5583 8823
rect 6009 8789 6043 8823
rect 8585 8789 8619 8823
rect 10057 8789 10091 8823
rect 11069 8789 11103 8823
rect 11621 8789 11655 8823
rect 11989 8789 12023 8823
rect 2053 8585 2087 8619
rect 5457 8585 5491 8619
rect 6837 8585 6871 8619
rect 7389 8585 7423 8619
rect 9045 8585 9079 8619
rect 9413 8585 9447 8619
rect 10425 8585 10459 8619
rect 10885 8585 10919 8619
rect 12449 8585 12483 8619
rect 21005 8585 21039 8619
rect 21373 8585 21407 8619
rect 2697 8517 2731 8551
rect 7757 8517 7791 8551
rect 10149 8517 10183 8551
rect 12909 8517 12943 8551
rect 1409 8449 1443 8483
rect 1869 8449 1903 8483
rect 2329 8449 2363 8483
rect 6745 8449 6779 8483
rect 7849 8449 7883 8483
rect 9505 8449 9539 8483
rect 10793 8449 10827 8483
rect 12817 8449 12851 8483
rect 7021 8381 7055 8415
rect 8033 8381 8067 8415
rect 8769 8381 8803 8415
rect 9689 8381 9723 8415
rect 10977 8381 11011 8415
rect 13093 8381 13127 8415
rect 1593 8313 1627 8347
rect 11529 8313 11563 8347
rect 6377 8245 6411 8279
rect 12081 8245 12115 8279
rect 2053 8041 2087 8075
rect 6009 8041 6043 8075
rect 7297 8041 7331 8075
rect 8953 8041 8987 8075
rect 10057 8041 10091 8075
rect 12265 8041 12299 8075
rect 1593 7973 1627 8007
rect 8401 7973 8435 8007
rect 2697 7905 2731 7939
rect 6469 7905 6503 7939
rect 6653 7905 6687 7939
rect 7757 7905 7791 7939
rect 7941 7905 7975 7939
rect 9597 7905 9631 7939
rect 12725 7905 12759 7939
rect 12817 7905 12851 7939
rect 1409 7837 1443 7871
rect 1869 7837 1903 7871
rect 2329 7837 2363 7871
rect 9321 7837 9355 7871
rect 12633 7837 12667 7871
rect 10425 7769 10459 7803
rect 6377 7701 6411 7735
rect 7665 7701 7699 7735
rect 9413 7701 9447 7735
rect 11897 7701 11931 7735
rect 1593 7497 1627 7531
rect 6653 7497 6687 7531
rect 7021 7497 7055 7531
rect 8033 7497 8067 7531
rect 8401 7497 8435 7531
rect 9505 7497 9539 7531
rect 8861 7429 8895 7463
rect 1409 7361 1443 7395
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 7389 7361 7423 7395
rect 8769 7361 8803 7395
rect 7481 7293 7515 7327
rect 7573 7293 7607 7327
rect 9045 7293 9079 7327
rect 2053 7225 2087 7259
rect 5917 7157 5951 7191
rect 9965 7157 9999 7191
rect 1869 6953 1903 6987
rect 8033 6953 8067 6987
rect 9045 6953 9079 6987
rect 10333 6953 10367 6987
rect 5365 6817 5399 6851
rect 7665 6817 7699 6851
rect 8493 6817 8527 6851
rect 9505 6817 9539 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 11437 6817 11471 6851
rect 1409 6749 1443 6783
rect 2237 6749 2271 6783
rect 5733 6749 5767 6783
rect 5917 6749 5951 6783
rect 7481 6749 7515 6783
rect 5181 6681 5215 6715
rect 6285 6681 6319 6715
rect 6469 6681 6503 6715
rect 1593 6613 1627 6647
rect 7021 6613 7055 6647
rect 7389 6613 7423 6647
rect 9413 6613 9447 6647
rect 10701 6613 10735 6647
rect 10793 6613 10827 6647
rect 1593 6409 1627 6443
rect 7849 6409 7883 6443
rect 9137 6409 9171 6443
rect 9597 6409 9631 6443
rect 10241 6409 10275 6443
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 8769 6273 8803 6307
rect 9505 6273 9539 6307
rect 9781 6205 9815 6239
rect 8401 6137 8435 6171
rect 2053 6069 2087 6103
rect 6653 6069 6687 6103
rect 7021 6069 7055 6103
rect 1869 5865 1903 5899
rect 1593 5797 1627 5831
rect 1409 5661 1443 5695
rect 2237 5661 2271 5695
rect 10977 5253 11011 5287
rect 11161 5253 11195 5287
rect 1961 5185 1995 5219
rect 2237 5117 2271 5151
rect 2513 5117 2547 5151
rect 1961 4641 1995 4675
rect 2237 4573 2271 4607
rect 2513 4573 2547 4607
rect 1501 4097 1535 4131
rect 2053 4097 2087 4131
rect 2513 4097 2547 4131
rect 1685 4029 1719 4063
rect 2237 3961 2271 3995
rect 1961 3689 1995 3723
rect 1685 3621 1719 3655
rect 1501 3417 1535 3451
rect 2329 3417 2363 3451
rect 2145 3145 2179 3179
rect 1685 3077 1719 3111
rect 1501 3009 1535 3043
rect 2053 3009 2087 3043
rect 2513 3009 2547 3043
rect 2881 2941 2915 2975
rect 2789 2533 2823 2567
rect 1961 2465 1995 2499
rect 2237 2397 2271 2431
rect 3801 2397 3835 2431
rect 11805 2397 11839 2431
rect 2605 2329 2639 2363
rect 3065 2329 3099 2363
rect 11621 2261 11655 2295
<< metal1 >>
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8662 20788 8668 20800
rect 8536 20760 8668 20788
rect 8536 20748 8542 20760
rect 8662 20748 8668 20760
rect 8720 20748 8726 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 18966 20788 18972 20800
rect 9732 20760 18972 20788
rect 9732 20748 9738 20760
rect 18966 20748 18972 20760
rect 19024 20748 19030 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 3142 20584 3148 20596
rect 3103 20556 3148 20584
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 3970 20584 3976 20596
rect 3931 20556 3976 20584
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 5626 20584 5632 20596
rect 4663 20556 5632 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 7098 20584 7104 20596
rect 5736 20556 7104 20584
rect 5736 20516 5764 20556
rect 7098 20544 7104 20556
rect 7156 20584 7162 20596
rect 7374 20584 7380 20596
rect 7156 20556 7380 20584
rect 7156 20544 7162 20556
rect 7374 20544 7380 20556
rect 7432 20544 7438 20596
rect 9398 20584 9404 20596
rect 8404 20556 9404 20584
rect 7282 20516 7288 20528
rect 4908 20488 5764 20516
rect 5828 20488 7288 20516
rect 198 20408 204 20460
rect 256 20448 262 20460
rect 1302 20448 1308 20460
rect 256 20420 1308 20448
rect 256 20408 262 20420
rect 1302 20408 1308 20420
rect 1360 20448 1366 20460
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 1360 20420 2237 20448
rect 1360 20408 1366 20420
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20417 2835 20451
rect 3326 20448 3332 20460
rect 3287 20420 3332 20448
rect 2777 20411 2835 20417
rect 1949 20383 2007 20389
rect 1949 20349 1961 20383
rect 1995 20380 2007 20383
rect 2682 20380 2688 20392
rect 1995 20352 2688 20380
rect 1995 20349 2007 20352
rect 1949 20343 2007 20349
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 2792 20380 2820 20411
rect 3326 20408 3332 20420
rect 3384 20408 3390 20460
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20448 3847 20451
rect 3878 20448 3884 20460
rect 3835 20420 3884 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4522 20448 4528 20460
rect 4479 20420 4528 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4522 20408 4528 20420
rect 4580 20448 4586 20460
rect 4908 20457 4936 20488
rect 4893 20451 4951 20457
rect 4580 20420 4844 20448
rect 4580 20408 4586 20420
rect 4706 20380 4712 20392
rect 2792 20352 4712 20380
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 4816 20380 4844 20420
rect 4893 20417 4905 20451
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 5442 20448 5448 20460
rect 5399 20420 5448 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 5828 20457 5856 20488
rect 7282 20476 7288 20488
rect 7340 20516 7346 20528
rect 8018 20516 8024 20528
rect 7340 20488 8024 20516
rect 7340 20476 7346 20488
rect 8018 20476 8024 20488
rect 8076 20476 8082 20528
rect 8404 20460 8432 20556
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 9674 20544 9680 20596
rect 9732 20584 9738 20596
rect 10689 20587 10747 20593
rect 9732 20556 9777 20584
rect 9732 20544 9738 20556
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 11054 20584 11060 20596
rect 10735 20556 11060 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 13136 20556 13369 20584
rect 13136 20544 13142 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 13357 20547 13415 20553
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13872 20556 14289 20584
rect 13872 20544 13878 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 14516 20556 15393 20584
rect 14516 20544 14522 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 15896 20556 16865 20584
rect 15896 20544 15902 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 17034 20544 17040 20596
rect 17092 20584 17098 20596
rect 17957 20587 18015 20593
rect 17957 20584 17969 20587
rect 17092 20556 17969 20584
rect 17092 20544 17098 20556
rect 17957 20553 17969 20556
rect 18003 20553 18015 20587
rect 17957 20547 18015 20553
rect 9858 20516 9864 20528
rect 9048 20488 9864 20516
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 6546 20448 6552 20460
rect 5813 20411 5871 20417
rect 6012 20420 6552 20448
rect 6012 20380 6040 20420
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 6730 20448 6736 20460
rect 6691 20420 6736 20448
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 7929 20451 7987 20457
rect 7515 20420 7880 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 4816 20352 6040 20380
rect 6086 20340 6092 20392
rect 6144 20380 6150 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6144 20352 6837 20380
rect 6144 20340 6150 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7742 20380 7748 20392
rect 7055 20352 7748 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7742 20340 7748 20352
rect 7800 20340 7806 20392
rect 4798 20272 4804 20324
rect 4856 20312 4862 20324
rect 6365 20315 6423 20321
rect 6365 20312 6377 20315
rect 4856 20284 6377 20312
rect 4856 20272 4862 20284
rect 6365 20281 6377 20284
rect 6411 20281 6423 20315
rect 7852 20312 7880 20420
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 8202 20448 8208 20460
rect 7975 20420 8208 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8386 20448 8392 20460
rect 8347 20420 8392 20448
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8570 20408 8576 20460
rect 8628 20448 8634 20460
rect 9048 20457 9076 20488
rect 9858 20476 9864 20488
rect 9916 20476 9922 20528
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 10008 20488 13216 20516
rect 10008 20476 10014 20488
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 8628 20420 9045 20448
rect 8628 20408 8634 20420
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 9493 20451 9551 20457
rect 9493 20417 9505 20451
rect 9539 20448 9551 20451
rect 9582 20448 9588 20460
rect 9539 20420 9588 20448
rect 9539 20417 9551 20420
rect 9493 20411 9551 20417
rect 9582 20408 9588 20420
rect 9640 20408 9646 20460
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10318 20448 10324 20460
rect 10091 20420 10324 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 10778 20448 10784 20460
rect 10551 20420 10784 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11238 20448 11244 20460
rect 11195 20420 11244 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11756 20420 11805 20448
rect 11756 20408 11762 20420
rect 11793 20417 11805 20420
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 12216 20420 12449 20448
rect 12216 20408 12222 20420
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 12437 20411 12495 20417
rect 12618 20408 12624 20460
rect 12676 20448 12682 20460
rect 13188 20457 13216 20488
rect 14366 20476 14372 20528
rect 14424 20516 14430 20528
rect 14424 20488 15792 20516
rect 14424 20476 14430 20488
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12676 20420 12909 20448
rect 12676 20408 12682 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 13320 20420 14105 20448
rect 13320 20408 13326 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14093 20411 14151 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15194 20448 15200 20460
rect 15155 20420 15200 20448
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15764 20457 15792 20488
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 8018 20340 8024 20392
rect 8076 20380 8082 20392
rect 16684 20380 16712 20411
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 16816 20420 17233 20448
rect 16816 20408 16822 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 17770 20448 17776 20460
rect 17731 20420 17776 20448
rect 17221 20411 17279 20417
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 17862 20408 17868 20460
rect 17920 20448 17926 20460
rect 18325 20451 18383 20457
rect 18325 20448 18337 20451
rect 17920 20420 18337 20448
rect 17920 20408 17926 20420
rect 18325 20417 18337 20420
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20714 20448 20720 20460
rect 20579 20420 20720 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20714 20408 20720 20420
rect 20772 20448 20778 20460
rect 22278 20448 22284 20460
rect 20772 20420 22284 20448
rect 20772 20408 20778 20420
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 8076 20352 9628 20380
rect 8076 20340 8082 20352
rect 8662 20312 8668 20324
rect 7852 20284 8668 20312
rect 6365 20275 6423 20281
rect 8662 20272 8668 20284
rect 8720 20312 8726 20324
rect 8720 20284 9168 20312
rect 8720 20272 8726 20284
rect 9140 20256 9168 20284
rect 2593 20247 2651 20253
rect 2593 20213 2605 20247
rect 2639 20244 2651 20247
rect 2774 20244 2780 20256
rect 2639 20216 2780 20244
rect 2639 20213 2651 20216
rect 2593 20207 2651 20213
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 5074 20244 5080 20256
rect 5035 20216 5080 20244
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5534 20244 5540 20256
rect 5495 20216 5540 20244
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 5994 20244 6000 20256
rect 5955 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 6822 20244 6828 20256
rect 6236 20216 6828 20244
rect 6236 20204 6242 20216
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7653 20247 7711 20253
rect 7653 20213 7665 20247
rect 7699 20244 7711 20247
rect 7742 20244 7748 20256
rect 7699 20216 7748 20244
rect 7699 20213 7711 20216
rect 7653 20207 7711 20213
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8294 20244 8300 20256
rect 8159 20216 8300 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8536 20216 8585 20244
rect 8536 20204 8542 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9122 20204 9128 20256
rect 9180 20204 9186 20256
rect 9217 20247 9275 20253
rect 9217 20213 9229 20247
rect 9263 20244 9275 20247
rect 9306 20244 9312 20256
rect 9263 20216 9312 20244
rect 9263 20213 9275 20216
rect 9217 20207 9275 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9600 20244 9628 20352
rect 13924 20352 16712 20380
rect 10594 20272 10600 20324
rect 10652 20312 10658 20324
rect 13924 20312 13952 20352
rect 17586 20340 17592 20392
rect 17644 20380 17650 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 17644 20352 19257 20380
rect 17644 20340 17650 20352
rect 19245 20349 19257 20352
rect 19291 20349 19303 20383
rect 19245 20343 19303 20349
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19794 20380 19800 20392
rect 19567 20352 19800 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21358 20380 21364 20392
rect 21223 20352 21364 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 10652 20284 13952 20312
rect 10652 20272 10658 20284
rect 13998 20272 14004 20324
rect 14056 20312 14062 20324
rect 14829 20315 14887 20321
rect 14829 20312 14841 20315
rect 14056 20284 14841 20312
rect 14056 20272 14062 20284
rect 14829 20281 14841 20284
rect 14875 20281 14887 20315
rect 14829 20275 14887 20281
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 15933 20315 15991 20321
rect 15933 20312 15945 20315
rect 14976 20284 15945 20312
rect 14976 20272 14982 20284
rect 15933 20281 15945 20284
rect 15979 20281 15991 20315
rect 15933 20275 15991 20281
rect 16298 20272 16304 20324
rect 16356 20312 16362 20324
rect 17405 20315 17463 20321
rect 17405 20312 17417 20315
rect 16356 20284 17417 20312
rect 16356 20272 16362 20284
rect 17405 20281 17417 20284
rect 17451 20281 17463 20315
rect 17405 20275 17463 20281
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 21266 20312 21272 20324
rect 17552 20284 21272 20312
rect 17552 20272 17558 20284
rect 21266 20272 21272 20284
rect 21324 20272 21330 20324
rect 9766 20244 9772 20256
rect 9600 20216 9772 20244
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 10229 20247 10287 20253
rect 10229 20213 10241 20247
rect 10275 20244 10287 20247
rect 10686 20244 10692 20256
rect 10275 20216 10692 20244
rect 10275 20213 10287 20216
rect 10229 20207 10287 20213
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 10962 20244 10968 20256
rect 10923 20216 10968 20244
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 11977 20247 12035 20253
rect 11977 20213 11989 20247
rect 12023 20244 12035 20247
rect 12066 20244 12072 20256
rect 12023 20216 12072 20244
rect 12023 20213 12035 20216
rect 11977 20207 12035 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 12250 20244 12256 20256
rect 12211 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12710 20244 12716 20256
rect 12671 20216 12716 20244
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 17276 20216 18521 20244
rect 17276 20204 17282 20216
rect 18509 20213 18521 20216
rect 18555 20213 18567 20247
rect 18509 20207 18567 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 8018 20040 8024 20052
rect 2746 20012 8024 20040
rect 2746 19916 2774 20012
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 8662 20000 8668 20052
rect 8720 20040 8726 20052
rect 9950 20040 9956 20052
rect 8720 20012 9956 20040
rect 8720 20000 8726 20012
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 10594 20040 10600 20052
rect 10555 20012 10600 20040
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 10965 20043 11023 20049
rect 10965 20009 10977 20043
rect 11011 20040 11023 20043
rect 11238 20040 11244 20052
rect 11011 20012 11244 20040
rect 11011 20009 11023 20012
rect 10965 20003 11023 20009
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11698 20040 11704 20052
rect 11659 20012 11704 20040
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 12158 20040 12164 20052
rect 12119 20012 12164 20040
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 12618 20040 12624 20052
rect 12579 20012 12624 20040
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 12894 20040 12900 20052
rect 12855 20012 12900 20040
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15436 20012 15669 20040
rect 15436 20000 15442 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 17494 20040 17500 20052
rect 16347 20012 17500 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 19429 20043 19487 20049
rect 19429 20040 19441 20043
rect 18288 20012 19441 20040
rect 18288 20000 18294 20012
rect 19429 20009 19441 20012
rect 19475 20009 19487 20043
rect 19429 20003 19487 20009
rect 6086 19932 6092 19984
rect 6144 19972 6150 19984
rect 6144 19944 6189 19972
rect 6144 19932 6150 19944
rect 6362 19932 6368 19984
rect 6420 19972 6426 19984
rect 6914 19972 6920 19984
rect 6420 19944 6920 19972
rect 6420 19932 6426 19944
rect 6914 19932 6920 19944
rect 6972 19932 6978 19984
rect 9217 19975 9275 19981
rect 9217 19941 9229 19975
rect 9263 19972 9275 19975
rect 9398 19972 9404 19984
rect 9263 19944 9404 19972
rect 9263 19941 9275 19944
rect 9217 19935 9275 19941
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 9674 19972 9680 19984
rect 9635 19944 9680 19972
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 10137 19975 10195 19981
rect 10137 19941 10149 19975
rect 10183 19941 10195 19975
rect 10137 19935 10195 19941
rect 658 19864 664 19916
rect 716 19904 722 19916
rect 1210 19904 1216 19916
rect 716 19876 1216 19904
rect 716 19864 722 19876
rect 1210 19864 1216 19876
rect 1268 19904 1274 19916
rect 1268 19876 2084 19904
rect 1268 19864 1274 19876
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19805 2007 19839
rect 2056 19836 2084 19876
rect 2682 19864 2688 19916
rect 2740 19876 2774 19916
rect 5258 19904 5264 19916
rect 4448 19876 5264 19904
rect 2740 19864 2746 19876
rect 4448 19848 4476 19876
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 6457 19907 6515 19913
rect 5583 19876 6408 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 2225 19839 2283 19845
rect 2225 19836 2237 19839
rect 2056 19808 2237 19836
rect 1949 19799 2007 19805
rect 2225 19805 2237 19808
rect 2271 19805 2283 19839
rect 2498 19836 2504 19848
rect 2459 19808 2504 19836
rect 2225 19799 2283 19805
rect 1964 19768 1992 19799
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3510 19836 3516 19848
rect 3283 19808 3516 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19805 4215 19839
rect 4430 19836 4436 19848
rect 4391 19808 4436 19836
rect 4157 19799 4215 19805
rect 2406 19768 2412 19780
rect 1964 19740 2412 19768
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 4172 19768 4200 19799
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 4614 19836 4620 19848
rect 4540 19808 4620 19836
rect 4540 19768 4568 19808
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 6178 19836 6184 19848
rect 4939 19808 6184 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 6380 19836 6408 19876
rect 6457 19873 6469 19907
rect 6503 19904 6515 19907
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 6503 19876 8125 19904
rect 6503 19873 6515 19876
rect 6457 19867 6515 19873
rect 8113 19873 8125 19876
rect 8159 19904 8171 19907
rect 10042 19904 10048 19916
rect 8159 19876 10048 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10152 19904 10180 19935
rect 10410 19932 10416 19984
rect 10468 19972 10474 19984
rect 16758 19972 16764 19984
rect 10468 19944 16764 19972
rect 10468 19932 10474 19944
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 18601 19907 18659 19913
rect 10152 19876 12434 19904
rect 8018 19836 8024 19848
rect 6380 19808 7880 19836
rect 7979 19808 8024 19836
rect 5629 19771 5687 19777
rect 5629 19768 5641 19771
rect 4172 19740 4568 19768
rect 4632 19740 5641 19768
rect 2685 19703 2743 19709
rect 2685 19669 2697 19703
rect 2731 19700 2743 19703
rect 2774 19700 2780 19712
rect 2731 19672 2780 19700
rect 2731 19669 2743 19672
rect 2685 19663 2743 19669
rect 2774 19660 2780 19672
rect 2832 19660 2838 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 3970 19700 3976 19712
rect 3931 19672 3976 19700
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 4632 19709 4660 19740
rect 5629 19737 5641 19740
rect 5675 19737 5687 19771
rect 5629 19731 5687 19737
rect 5721 19771 5779 19777
rect 5721 19737 5733 19771
rect 5767 19768 5779 19771
rect 6362 19768 6368 19780
rect 5767 19740 6368 19768
rect 5767 19737 5779 19740
rect 5721 19731 5779 19737
rect 6362 19728 6368 19740
rect 6420 19728 6426 19780
rect 6546 19728 6552 19780
rect 6604 19768 6610 19780
rect 7852 19768 7880 19808
rect 8018 19796 8024 19808
rect 8076 19796 8082 19848
rect 9033 19839 9091 19845
rect 9033 19805 9045 19839
rect 9079 19836 9091 19839
rect 9122 19836 9128 19848
rect 9079 19808 9128 19836
rect 9079 19805 9091 19808
rect 9033 19799 9091 19805
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 9490 19836 9496 19848
rect 9451 19808 9496 19836
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19836 10011 19839
rect 10134 19836 10140 19848
rect 9999 19808 10140 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 10226 19796 10232 19848
rect 10284 19836 10290 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10284 19808 10425 19836
rect 10284 19796 10290 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 10413 19799 10471 19805
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 12406 19836 12434 19876
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 19978 19904 19984 19916
rect 18647 19876 19984 19904
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 21358 19904 21364 19916
rect 21319 19876 21364 19904
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 12406 19808 15485 19836
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 15896 19808 16129 19836
rect 15896 19796 15902 19808
rect 16117 19805 16129 19808
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 6604 19740 6776 19768
rect 7852 19740 9352 19768
rect 6604 19728 6610 19740
rect 4617 19703 4675 19709
rect 4617 19669 4629 19703
rect 4663 19669 4675 19703
rect 4617 19663 4675 19669
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5350 19700 5356 19712
rect 5123 19672 5356 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5810 19660 5816 19712
rect 5868 19700 5874 19712
rect 6748 19709 6776 19740
rect 6641 19703 6699 19709
rect 6641 19700 6653 19703
rect 5868 19672 6653 19700
rect 5868 19660 5874 19672
rect 6641 19669 6653 19672
rect 6687 19669 6699 19703
rect 6641 19663 6699 19669
rect 6733 19703 6791 19709
rect 6733 19669 6745 19703
rect 6779 19669 6791 19703
rect 6733 19663 6791 19669
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 7466 19700 7472 19712
rect 7147 19672 7472 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 7926 19700 7932 19712
rect 7616 19672 7661 19700
rect 7887 19672 7932 19700
rect 7616 19660 7622 19672
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 9324 19700 9352 19740
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 13357 19771 13415 19777
rect 9456 19740 13308 19768
rect 9456 19728 9462 19740
rect 10502 19700 10508 19712
rect 9324 19672 10508 19700
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19700 11483 19703
rect 11882 19700 11888 19712
rect 11471 19672 11888 19700
rect 11471 19669 11483 19672
rect 11425 19663 11483 19669
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 13280 19700 13308 19740
rect 13357 19737 13369 19771
rect 13403 19768 13415 19771
rect 13722 19768 13728 19780
rect 13403 19740 13728 19768
rect 13403 19737 13415 19740
rect 13357 19731 13415 19737
rect 13722 19728 13728 19740
rect 13780 19768 13786 19780
rect 14185 19771 14243 19777
rect 14185 19768 14197 19771
rect 13780 19740 14197 19768
rect 13780 19728 13786 19740
rect 14185 19737 14197 19740
rect 14231 19768 14243 19771
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 14231 19740 14565 19768
rect 14231 19737 14243 19740
rect 14185 19731 14243 19737
rect 14553 19737 14565 19740
rect 14599 19768 14611 19771
rect 14599 19740 15516 19768
rect 14599 19737 14611 19740
rect 14553 19731 14611 19737
rect 15488 19712 15516 19740
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16684 19768 16712 19799
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19024 19808 19257 19836
rect 19024 19796 19030 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 15804 19740 16712 19768
rect 16868 19740 18276 19768
rect 15804 19728 15810 19740
rect 14366 19700 14372 19712
rect 13280 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 15194 19700 15200 19712
rect 15155 19672 15200 19700
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 15470 19660 15476 19712
rect 15528 19660 15534 19712
rect 16868 19709 16896 19740
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 17221 19703 17279 19709
rect 17221 19669 17233 19703
rect 17267 19700 17279 19703
rect 17310 19700 17316 19712
rect 17267 19672 17316 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 18248 19700 18276 19740
rect 18322 19728 18328 19780
rect 18380 19777 18386 19780
rect 18380 19768 18392 19777
rect 21116 19771 21174 19777
rect 18380 19740 18425 19768
rect 18380 19731 18392 19740
rect 21116 19737 21128 19771
rect 21162 19768 21174 19771
rect 21266 19768 21272 19780
rect 21162 19740 21272 19768
rect 21162 19737 21174 19740
rect 21116 19731 21174 19737
rect 18380 19728 18386 19731
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 19886 19700 19892 19712
rect 18248 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 19981 19703 20039 19709
rect 19981 19669 19993 19703
rect 20027 19700 20039 19703
rect 20070 19700 20076 19712
rect 20027 19672 20076 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2498 19496 2504 19508
rect 2459 19468 2504 19496
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 3605 19499 3663 19505
rect 3605 19465 3617 19499
rect 3651 19496 3663 19499
rect 4982 19496 4988 19508
rect 3651 19468 4988 19496
rect 3651 19465 3663 19468
rect 3605 19459 3663 19465
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 5408 19468 6040 19496
rect 5408 19456 5414 19468
rect 4522 19388 4528 19440
rect 4580 19428 4586 19440
rect 5902 19428 5908 19440
rect 4580 19400 5908 19428
rect 4580 19388 4586 19400
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 6012 19428 6040 19468
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6638 19496 6644 19508
rect 6144 19468 6644 19496
rect 6144 19456 6150 19468
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 6825 19499 6883 19505
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 7466 19496 7472 19508
rect 6871 19468 7328 19496
rect 7427 19468 7472 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 6362 19428 6368 19440
rect 6012 19400 6368 19428
rect 6362 19388 6368 19400
rect 6420 19388 6426 19440
rect 6454 19388 6460 19440
rect 6512 19428 6518 19440
rect 6914 19428 6920 19440
rect 6512 19400 6920 19428
rect 6512 19388 6518 19400
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 1946 19360 1952 19372
rect 1907 19332 1952 19360
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2866 19360 2872 19372
rect 2731 19332 2872 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 3234 19360 3240 19372
rect 3007 19332 3240 19360
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3418 19360 3424 19372
rect 3379 19332 3424 19360
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19360 4215 19363
rect 4338 19360 4344 19372
rect 4203 19332 4344 19360
rect 4203 19329 4215 19332
rect 4157 19323 4215 19329
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 4798 19360 4804 19372
rect 4759 19332 4804 19360
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 5537 19363 5595 19369
rect 5537 19329 5549 19363
rect 5583 19360 5595 19363
rect 5718 19360 5724 19372
rect 5583 19332 5724 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 5718 19320 5724 19332
rect 5776 19320 5782 19372
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 6638 19360 6644 19372
rect 5859 19332 6500 19360
rect 6599 19332 6644 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 1118 19252 1124 19304
rect 1176 19292 1182 19304
rect 4522 19292 4528 19304
rect 1176 19264 4528 19292
rect 1176 19252 1182 19264
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 6086 19292 6092 19304
rect 6012 19264 6092 19292
rect 2130 19224 2136 19236
rect 2091 19196 2136 19224
rect 2130 19184 2136 19196
rect 2188 19184 2194 19236
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 6012 19233 6040 19264
rect 6086 19252 6092 19264
rect 6144 19252 6150 19304
rect 6472 19292 6500 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7300 19360 7328 19468
rect 7466 19456 7472 19468
rect 7524 19456 7530 19508
rect 8662 19496 8668 19508
rect 8623 19468 8668 19496
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 9398 19496 9404 19508
rect 9171 19468 9404 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 9858 19496 9864 19508
rect 9631 19468 9864 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 10045 19499 10103 19505
rect 10045 19465 10057 19499
rect 10091 19496 10103 19499
rect 10410 19496 10416 19508
rect 10091 19468 10416 19496
rect 10091 19465 10103 19468
rect 10045 19459 10103 19465
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19465 10563 19499
rect 10778 19496 10784 19508
rect 10739 19468 10784 19496
rect 10505 19459 10563 19465
rect 7377 19431 7435 19437
rect 7377 19397 7389 19431
rect 7423 19428 7435 19431
rect 7558 19428 7564 19440
rect 7423 19400 7564 19428
rect 7423 19397 7435 19400
rect 7377 19391 7435 19397
rect 7558 19388 7564 19400
rect 7616 19388 7622 19440
rect 9674 19428 9680 19440
rect 7668 19400 9680 19428
rect 7668 19360 7696 19400
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 10520 19428 10548 19459
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 13872 19468 14105 19496
rect 13872 19456 13878 19468
rect 14093 19465 14105 19468
rect 14139 19465 14151 19499
rect 14093 19459 14151 19465
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15746 19496 15752 19508
rect 15252 19468 15752 19496
rect 15252 19456 15258 19468
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 18049 19499 18107 19505
rect 18049 19496 18061 19499
rect 17460 19468 18061 19496
rect 17460 19456 17466 19468
rect 18049 19465 18061 19468
rect 18095 19465 18107 19499
rect 18049 19459 18107 19465
rect 18598 19456 18604 19508
rect 18656 19496 18662 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 18656 19468 19073 19496
rect 18656 19456 18662 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 14642 19428 14648 19440
rect 10520 19400 14648 19428
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 20036 19400 21128 19428
rect 20036 19388 20042 19400
rect 8478 19360 8484 19372
rect 7300 19332 7696 19360
rect 8439 19332 8484 19360
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19360 8999 19363
rect 9401 19363 9459 19369
rect 8987 19332 9352 19360
rect 8987 19329 8999 19332
rect 8941 19323 8999 19329
rect 9324 19304 9352 19332
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9858 19360 9864 19372
rect 9447 19332 9628 19360
rect 9819 19332 9864 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 7098 19292 7104 19304
rect 6472 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19292 7343 19295
rect 7558 19292 7564 19304
rect 7331 19264 7564 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 7558 19252 7564 19264
rect 7616 19292 7622 19304
rect 8110 19292 8116 19304
rect 7616 19264 8116 19292
rect 7616 19252 7622 19264
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19292 8263 19295
rect 8570 19292 8576 19304
rect 8251 19264 8576 19292
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 4617 19227 4675 19233
rect 4617 19224 4629 19227
rect 4212 19196 4629 19224
rect 4212 19184 4218 19196
rect 4617 19193 4629 19196
rect 4663 19193 4675 19227
rect 4617 19187 4675 19193
rect 5997 19227 6055 19233
rect 5997 19193 6009 19227
rect 6043 19193 6055 19227
rect 5997 19187 6055 19193
rect 7374 19184 7380 19236
rect 7432 19224 7438 19236
rect 8662 19224 8668 19236
rect 7432 19196 8668 19224
rect 7432 19184 7438 19196
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 9600 19224 9628 19332
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10336 19292 10364 19323
rect 13538 19320 13544 19372
rect 13596 19369 13602 19372
rect 13596 19360 13608 19369
rect 13596 19332 13641 19360
rect 13596 19323 13608 19332
rect 13596 19320 13602 19323
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13780 19332 13829 19360
rect 13780 19320 13786 19332
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 15206 19363 15264 19369
rect 15206 19360 15218 19363
rect 14516 19332 15218 19360
rect 14516 19320 14522 19332
rect 15206 19329 15218 19332
rect 15252 19329 15264 19363
rect 16925 19363 16983 19369
rect 16925 19360 16937 19363
rect 15206 19323 15264 19329
rect 16546 19332 16937 19360
rect 9732 19264 10364 19292
rect 9732 19252 9738 19264
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 11609 19295 11667 19301
rect 11609 19292 11621 19295
rect 10836 19264 11621 19292
rect 10836 19252 10842 19264
rect 11609 19261 11621 19264
rect 11655 19292 11667 19295
rect 12802 19292 12808 19304
rect 11655 19264 12808 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 9766 19224 9772 19236
rect 9600 19196 9772 19224
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 15488 19168 15516 19255
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 16546 19292 16574 19332
rect 16925 19329 16937 19332
rect 16971 19329 16983 19363
rect 16925 19323 16983 19329
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 18012 19332 18337 19360
rect 18012 19320 18018 19332
rect 18325 19329 18337 19332
rect 18371 19329 18383 19363
rect 18874 19360 18880 19372
rect 18835 19332 18880 19360
rect 18325 19323 18383 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 20806 19320 20812 19372
rect 20864 19369 20870 19372
rect 21100 19369 21128 19400
rect 20864 19360 20876 19369
rect 21085 19363 21143 19369
rect 20864 19332 20909 19360
rect 20864 19323 20876 19332
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21358 19360 21364 19372
rect 21131 19332 21364 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 20864 19320 20870 19323
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 16172 19264 16574 19292
rect 16669 19295 16727 19301
rect 16172 19252 16178 19264
rect 16669 19261 16681 19295
rect 16715 19261 16727 19295
rect 16669 19255 16727 19261
rect 16684 19224 16712 19255
rect 15764 19196 16712 19224
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 3142 19156 3148 19168
rect 3103 19128 3148 19156
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 4304 19128 4353 19156
rect 4304 19116 4310 19128
rect 4341 19125 4353 19128
rect 4387 19125 4399 19159
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 4341 19119 4399 19125
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 5442 19116 5448 19168
rect 5500 19156 5506 19168
rect 7650 19156 7656 19168
rect 5500 19128 7656 19156
rect 5500 19116 5506 19128
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 7834 19156 7840 19168
rect 7795 19128 7840 19156
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 11977 19159 12035 19165
rect 11977 19156 11989 19159
rect 9272 19128 11989 19156
rect 9272 19116 9278 19128
rect 11977 19125 11989 19128
rect 12023 19125 12035 19159
rect 11977 19119 12035 19125
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13630 19156 13636 19168
rect 12492 19128 13636 19156
rect 12492 19116 12498 19128
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 15470 19116 15476 19168
rect 15528 19156 15534 19168
rect 15764 19165 15792 19196
rect 17678 19184 17684 19236
rect 17736 19224 17742 19236
rect 18509 19227 18567 19233
rect 18509 19224 18521 19227
rect 17736 19196 18521 19224
rect 17736 19184 17742 19196
rect 18509 19193 18521 19196
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 19536 19196 20208 19224
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 15528 19128 15761 19156
rect 15528 19116 15534 19128
rect 15749 19125 15761 19128
rect 15795 19125 15807 19159
rect 15749 19119 15807 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15896 19128 16129 19156
rect 15896 19116 15902 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 19536 19156 19564 19196
rect 19702 19156 19708 19168
rect 17644 19128 19564 19156
rect 19663 19128 19708 19156
rect 17644 19116 17650 19128
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20180 19156 20208 19196
rect 22738 19156 22744 19168
rect 20180 19128 22744 19156
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 1728 18924 2513 18952
rect 1728 18912 1734 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3384 18924 3801 18952
rect 3384 18912 3390 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 5166 18952 5172 18964
rect 3789 18915 3847 18921
rect 3896 18924 5172 18952
rect 2038 18844 2044 18896
rect 2096 18884 2102 18896
rect 2133 18887 2191 18893
rect 2133 18884 2145 18887
rect 2096 18856 2145 18884
rect 2096 18844 2102 18856
rect 2133 18853 2145 18856
rect 2179 18853 2191 18887
rect 2133 18847 2191 18853
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 3896 18884 3924 18924
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 5353 18955 5411 18961
rect 5353 18921 5365 18955
rect 5399 18952 5411 18955
rect 5534 18952 5540 18964
rect 5399 18924 5540 18952
rect 5399 18921 5411 18924
rect 5353 18915 5411 18921
rect 5534 18912 5540 18924
rect 5592 18952 5598 18964
rect 5810 18952 5816 18964
rect 5592 18924 5816 18952
rect 5592 18912 5598 18924
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18952 7435 18955
rect 7423 18924 8064 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 7837 18887 7895 18893
rect 7837 18884 7849 18887
rect 2280 18856 3924 18884
rect 5276 18856 7849 18884
rect 2280 18844 2286 18856
rect 1578 18776 1584 18828
rect 1636 18816 1642 18828
rect 5276 18816 5304 18856
rect 7837 18853 7849 18856
rect 7883 18853 7895 18887
rect 7837 18847 7895 18853
rect 1636 18788 4384 18816
rect 1636 18776 1642 18788
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1688 18612 1716 18711
rect 1854 18708 1860 18760
rect 1912 18748 1918 18760
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1912 18720 1961 18748
rect 1912 18708 1918 18720
rect 1949 18717 1961 18720
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18717 2743 18751
rect 3050 18748 3056 18760
rect 3011 18720 3056 18748
rect 2685 18711 2743 18717
rect 2700 18680 2728 18711
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 4154 18748 4160 18760
rect 4019 18720 4160 18748
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 4356 18680 4384 18788
rect 4448 18788 5304 18816
rect 6181 18819 6239 18825
rect 4448 18757 4476 18788
rect 6181 18785 6193 18819
rect 6227 18816 6239 18819
rect 6730 18816 6736 18828
rect 6227 18788 6736 18816
rect 6227 18785 6239 18788
rect 6181 18779 6239 18785
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18816 6883 18819
rect 6914 18816 6920 18828
rect 6871 18788 6920 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 8036 18816 8064 18924
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 8444 18924 9352 18952
rect 8444 18912 8450 18924
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 9324 18884 9352 18924
rect 9582 18912 9588 18964
rect 9640 18952 9646 18964
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 9640 18924 9781 18952
rect 9640 18912 9646 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 10318 18952 10324 18964
rect 10279 18924 10324 18952
rect 9769 18915 9827 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 18785 18955 18843 18961
rect 11940 18924 18644 18952
rect 11940 18912 11946 18924
rect 11057 18887 11115 18893
rect 11057 18884 11069 18887
rect 8168 18856 8708 18884
rect 9324 18856 11069 18884
rect 8168 18844 8174 18856
rect 8481 18819 8539 18825
rect 8036 18788 8340 18816
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 4982 18748 4988 18760
rect 4939 18720 4988 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5721 18751 5779 18757
rect 5224 18720 5396 18748
rect 5224 18708 5230 18720
rect 5258 18680 5264 18692
rect 2700 18652 4292 18680
rect 4356 18652 5264 18680
rect 2682 18612 2688 18624
rect 1688 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3237 18615 3295 18621
rect 3237 18581 3249 18615
rect 3283 18612 3295 18615
rect 3786 18612 3792 18624
rect 3283 18584 3792 18612
rect 3283 18581 3295 18584
rect 3237 18575 3295 18581
rect 3786 18572 3792 18584
rect 3844 18612 3850 18624
rect 4062 18612 4068 18624
rect 3844 18584 4068 18612
rect 3844 18572 3850 18584
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 4264 18621 4292 18652
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18581 4307 18615
rect 4706 18612 4712 18624
rect 4667 18584 4712 18612
rect 4249 18575 4307 18581
rect 4706 18572 4712 18584
rect 4764 18572 4770 18624
rect 5368 18612 5396 18720
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 8202 18748 8208 18760
rect 5767 18744 5856 18748
rect 5920 18744 8208 18748
rect 5767 18720 8208 18744
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 5828 18716 5948 18720
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8312 18748 8340 18788
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 8570 18816 8576 18828
rect 8527 18788 8576 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 8680 18816 8708 18856
rect 11057 18853 11069 18856
rect 11103 18853 11115 18887
rect 12618 18884 12624 18896
rect 11057 18847 11115 18853
rect 11440 18856 12624 18884
rect 10778 18816 10784 18828
rect 8680 18788 10784 18816
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 9033 18751 9091 18757
rect 8312 18720 8432 18748
rect 6914 18680 6920 18692
rect 6827 18652 6920 18680
rect 6914 18640 6920 18652
rect 6972 18680 6978 18692
rect 7926 18680 7932 18692
rect 6972 18652 7932 18680
rect 6972 18640 6978 18652
rect 7926 18640 7932 18652
rect 7984 18640 7990 18692
rect 8110 18640 8116 18692
rect 8168 18680 8174 18692
rect 8297 18683 8355 18689
rect 8297 18680 8309 18683
rect 8168 18652 8309 18680
rect 8168 18640 8174 18652
rect 8297 18649 8309 18652
rect 8343 18649 8355 18683
rect 8297 18643 8355 18649
rect 5718 18612 5724 18624
rect 5368 18584 5724 18612
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 6822 18612 6828 18624
rect 5868 18584 6828 18612
rect 5868 18572 5874 18584
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 8202 18612 8208 18624
rect 7064 18584 7109 18612
rect 8163 18584 8208 18612
rect 7064 18572 7070 18584
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8404 18612 8432 18720
rect 9033 18717 9045 18751
rect 9079 18748 9091 18751
rect 9582 18748 9588 18760
rect 9079 18720 9588 18748
rect 9079 18717 9091 18720
rect 9033 18711 9091 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9950 18748 9956 18760
rect 9911 18720 9956 18748
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10318 18748 10324 18760
rect 10100 18720 10324 18748
rect 10100 18708 10106 18720
rect 10318 18708 10324 18720
rect 10376 18748 10382 18760
rect 11440 18757 11468 18856
rect 12618 18844 12624 18856
rect 12676 18844 12682 18896
rect 13722 18816 13728 18828
rect 13683 18788 13728 18816
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 18138 18816 18144 18828
rect 17543 18788 18144 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 10376 18720 10701 18748
rect 10376 18708 10382 18720
rect 10689 18717 10701 18720
rect 10735 18748 10747 18751
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 10735 18720 11437 18748
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 11425 18717 11437 18720
rect 11471 18717 11483 18751
rect 15470 18748 15476 18760
rect 11425 18711 11483 18717
rect 11716 18720 15332 18748
rect 15431 18720 15476 18748
rect 9030 18612 9036 18624
rect 8404 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9217 18615 9275 18621
rect 9217 18581 9229 18615
rect 9263 18612 9275 18615
rect 11716 18612 11744 18720
rect 13446 18640 13452 18692
rect 13504 18689 13510 18692
rect 13504 18680 13516 18689
rect 13504 18652 13549 18680
rect 13504 18643 13516 18652
rect 13504 18640 13510 18643
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 15206 18683 15264 18689
rect 15206 18680 15218 18683
rect 13688 18652 15218 18680
rect 13688 18640 13694 18652
rect 15206 18649 15218 18652
rect 15252 18649 15264 18683
rect 15304 18680 15332 18720
rect 15470 18708 15476 18720
rect 15528 18748 15534 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15528 18720 15761 18748
rect 15528 18708 15534 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 18046 18748 18052 18760
rect 18007 18720 18052 18748
rect 15749 18711 15807 18717
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18616 18757 18644 18924
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 19058 18952 19064 18964
rect 18831 18924 19064 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 19518 18912 19524 18964
rect 19576 18952 19582 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 19576 18924 21097 18952
rect 19576 18912 19582 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21085 18915 21143 18921
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18748 19303 18751
rect 19978 18748 19984 18760
rect 19291 18720 19984 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21174 18748 21180 18760
rect 20947 18720 21180 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 15304 18652 16252 18680
rect 15206 18643 15264 18649
rect 11974 18612 11980 18624
rect 9263 18584 11744 18612
rect 11935 18584 11980 18612
rect 9263 18581 9275 18584
rect 9217 18575 9275 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 12216 18584 12357 18612
rect 12216 18572 12222 18584
rect 12345 18581 12357 18584
rect 12391 18581 12403 18615
rect 12345 18575 12403 18581
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13136 18584 14105 18612
rect 13136 18572 13142 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 14093 18575 14151 18581
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16224 18612 16252 18652
rect 17126 18640 17132 18692
rect 17184 18680 17190 18692
rect 17230 18683 17288 18689
rect 17230 18680 17242 18683
rect 17184 18652 17242 18680
rect 17184 18640 17190 18652
rect 17230 18649 17242 18652
rect 17276 18649 17288 18683
rect 17230 18643 17288 18649
rect 19512 18683 19570 18689
rect 19512 18649 19524 18683
rect 19558 18680 19570 18683
rect 19702 18680 19708 18692
rect 19558 18652 19708 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 17954 18612 17960 18624
rect 16224 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 20438 18612 20444 18624
rect 18279 18584 20444 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 20622 18612 20628 18624
rect 20583 18584 20628 18612
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18377 2651 18411
rect 2593 18371 2651 18377
rect 2608 18340 2636 18371
rect 3234 18368 3240 18420
rect 3292 18408 3298 18420
rect 3513 18411 3571 18417
rect 3292 18380 3464 18408
rect 3292 18368 3298 18380
rect 2608 18312 3372 18340
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2314 18272 2320 18284
rect 2179 18244 2320 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18241 2467 18275
rect 2409 18235 2467 18241
rect 2424 18204 2452 18235
rect 2590 18232 2596 18284
rect 2648 18272 2654 18284
rect 3344 18281 3372 18312
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2648 18244 2881 18272
rect 2648 18232 2654 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 3329 18275 3387 18281
rect 3329 18241 3341 18275
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 3234 18204 3240 18216
rect 2424 18176 3240 18204
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3436 18204 3464 18380
rect 3513 18377 3525 18411
rect 3559 18408 3571 18411
rect 3878 18408 3884 18420
rect 3559 18380 3884 18408
rect 3559 18377 3571 18380
rect 3513 18371 3571 18377
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 4522 18368 4528 18420
rect 4580 18408 4586 18420
rect 5629 18411 5687 18417
rect 4580 18380 5488 18408
rect 4580 18368 4586 18380
rect 4062 18272 4068 18284
rect 4023 18244 4068 18272
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18272 5227 18275
rect 5258 18272 5264 18284
rect 5215 18244 5264 18272
rect 5215 18241 5227 18244
rect 5169 18235 5227 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5460 18281 5488 18380
rect 5629 18377 5641 18411
rect 5675 18408 5687 18411
rect 6914 18408 6920 18420
rect 5675 18380 6920 18408
rect 5675 18377 5687 18380
rect 5629 18371 5687 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 7561 18411 7619 18417
rect 7561 18377 7573 18411
rect 7607 18408 7619 18411
rect 7834 18408 7840 18420
rect 7607 18380 7840 18408
rect 7607 18377 7619 18380
rect 7561 18371 7619 18377
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8021 18411 8079 18417
rect 8021 18377 8033 18411
rect 8067 18408 8079 18411
rect 8067 18380 8156 18408
rect 8067 18377 8079 18380
rect 8021 18371 8079 18377
rect 5902 18300 5908 18352
rect 5960 18340 5966 18352
rect 6178 18340 6184 18352
rect 5960 18312 6184 18340
rect 5960 18300 5966 18312
rect 6178 18300 6184 18312
rect 6236 18300 6242 18352
rect 6822 18300 6828 18352
rect 6880 18340 6886 18352
rect 7190 18340 7196 18352
rect 6880 18312 7196 18340
rect 6880 18300 6886 18312
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 7650 18340 7656 18352
rect 7611 18312 7656 18340
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 5445 18275 5503 18281
rect 5445 18241 5457 18275
rect 5491 18272 5503 18275
rect 5994 18272 6000 18284
rect 5491 18244 6000 18272
rect 5491 18241 5503 18244
rect 5445 18235 5503 18241
rect 5994 18232 6000 18244
rect 6052 18232 6058 18284
rect 8128 18272 8156 18380
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8260 18380 8309 18408
rect 8260 18368 8266 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 9585 18411 9643 18417
rect 9585 18408 9597 18411
rect 9548 18380 9597 18408
rect 9548 18368 9554 18380
rect 9585 18377 9597 18380
rect 9631 18377 9643 18411
rect 9585 18371 9643 18377
rect 12802 18368 12808 18420
rect 12860 18408 12866 18420
rect 12860 18380 13501 18408
rect 12860 18368 12866 18380
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 10873 18343 10931 18349
rect 10873 18340 10885 18343
rect 9088 18312 10885 18340
rect 9088 18300 9094 18312
rect 10873 18309 10885 18312
rect 10919 18309 10931 18343
rect 10873 18303 10931 18309
rect 12980 18343 13038 18349
rect 12980 18309 12992 18343
rect 13026 18340 13038 18343
rect 13078 18340 13084 18352
rect 13026 18312 13084 18340
rect 13026 18309 13038 18312
rect 12980 18303 13038 18309
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 13473 18340 13501 18380
rect 13538 18368 13544 18420
rect 13596 18408 13602 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 13596 18380 16681 18408
rect 13596 18368 13602 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 20070 18408 20076 18420
rect 16669 18371 16727 18377
rect 17052 18380 20076 18408
rect 14826 18340 14832 18352
rect 13473 18312 14832 18340
rect 14826 18300 14832 18312
rect 14884 18300 14890 18352
rect 15504 18343 15562 18349
rect 15504 18309 15516 18343
rect 15550 18340 15562 18343
rect 15654 18340 15660 18352
rect 15550 18312 15660 18340
rect 15550 18309 15562 18312
rect 15504 18303 15562 18309
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 8757 18275 8815 18281
rect 8757 18272 8769 18275
rect 6104 18244 7604 18272
rect 8128 18244 8769 18272
rect 4522 18204 4528 18216
rect 3436 18176 4016 18204
rect 4483 18176 4528 18204
rect 2866 18096 2872 18148
rect 2924 18136 2930 18148
rect 3881 18139 3939 18145
rect 3881 18136 3893 18139
rect 2924 18108 3893 18136
rect 2924 18096 2930 18108
rect 3881 18105 3893 18108
rect 3927 18105 3939 18139
rect 3988 18136 4016 18176
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 6104 18204 6132 18244
rect 4632 18176 6132 18204
rect 4632 18136 4660 18176
rect 6178 18164 6184 18216
rect 6236 18204 6242 18216
rect 7466 18204 7472 18216
rect 6236 18176 7052 18204
rect 7427 18176 7472 18204
rect 6236 18164 6242 18176
rect 3988 18108 4660 18136
rect 3881 18099 3939 18105
rect 5166 18096 5172 18148
rect 5224 18136 5230 18148
rect 5905 18139 5963 18145
rect 5905 18136 5917 18139
rect 5224 18108 5917 18136
rect 5224 18096 5230 18108
rect 5905 18105 5917 18108
rect 5951 18105 5963 18139
rect 7024 18136 7052 18176
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7576 18204 7604 18244
rect 8757 18241 8769 18244
rect 8803 18241 8815 18275
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 8757 18235 8815 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 10781 18275 10839 18281
rect 10781 18241 10793 18275
rect 10827 18272 10839 18275
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 10827 18244 11529 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 15749 18275 15807 18281
rect 11517 18235 11575 18241
rect 11716 18244 15700 18272
rect 9490 18204 9496 18216
rect 7576 18176 9496 18204
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 10042 18204 10048 18216
rect 9999 18176 10048 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 11716 18204 11744 18244
rect 11011 18176 11744 18204
rect 12713 18207 12771 18213
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 12713 18173 12725 18207
rect 12759 18173 12771 18207
rect 15672 18204 15700 18244
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 16206 18272 16212 18284
rect 15795 18244 16212 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 17052 18204 17080 18380
rect 20070 18368 20076 18380
rect 20128 18408 20134 18420
rect 20990 18408 20996 18420
rect 20128 18380 20996 18408
rect 20128 18368 20134 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21358 18408 21364 18420
rect 21319 18380 21364 18408
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 19610 18300 19616 18352
rect 19668 18340 19674 18352
rect 21634 18340 21640 18352
rect 19668 18312 21640 18340
rect 19668 18300 19674 18312
rect 21634 18300 21640 18312
rect 21692 18300 21698 18352
rect 17402 18232 17408 18284
rect 17460 18272 17466 18284
rect 17782 18275 17840 18281
rect 17782 18272 17794 18275
rect 17460 18244 17794 18272
rect 17460 18232 17466 18244
rect 17782 18241 17794 18244
rect 17828 18241 17840 18275
rect 17782 18235 17840 18241
rect 19426 18232 19432 18284
rect 19484 18281 19490 18284
rect 19484 18272 19496 18281
rect 19705 18275 19763 18281
rect 19484 18244 19529 18272
rect 19484 18235 19496 18244
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 19978 18272 19984 18284
rect 19751 18244 19984 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 19484 18232 19490 18235
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20070 18232 20076 18284
rect 20128 18272 20134 18284
rect 20237 18275 20295 18281
rect 20237 18272 20249 18275
rect 20128 18244 20249 18272
rect 20128 18232 20134 18244
rect 20237 18241 20249 18244
rect 20283 18272 20295 18275
rect 20622 18272 20628 18284
rect 20283 18244 20628 18272
rect 20283 18241 20295 18244
rect 20237 18235 20295 18241
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 18046 18204 18052 18216
rect 15672 18176 17080 18204
rect 18007 18176 18052 18204
rect 12713 18167 12771 18173
rect 7834 18136 7840 18148
rect 5905 18099 5963 18105
rect 6012 18108 6960 18136
rect 7024 18108 7840 18136
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 3053 18071 3111 18077
rect 3053 18037 3065 18071
rect 3099 18068 3111 18071
rect 3326 18068 3332 18080
rect 3099 18040 3332 18068
rect 3099 18037 3111 18040
rect 3053 18031 3111 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 4706 18028 4712 18080
rect 4764 18068 4770 18080
rect 4985 18071 5043 18077
rect 4985 18068 4997 18071
rect 4764 18040 4997 18068
rect 4764 18028 4770 18040
rect 4985 18037 4997 18040
rect 5031 18037 5043 18071
rect 4985 18031 5043 18037
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 6012 18068 6040 18108
rect 6362 18068 6368 18080
rect 5500 18040 6040 18068
rect 6323 18040 6368 18068
rect 5500 18028 5506 18040
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6822 18068 6828 18080
rect 6783 18040 6828 18068
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 6932 18068 6960 18108
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 8941 18139 8999 18145
rect 8941 18105 8953 18139
rect 8987 18136 8999 18139
rect 9674 18136 9680 18148
rect 8987 18108 9680 18136
rect 8987 18105 8999 18108
rect 8941 18099 8999 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 11330 18136 11336 18148
rect 9784 18108 11336 18136
rect 9784 18068 9812 18108
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 6932 18040 9812 18068
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 10100 18040 10425 18068
rect 10100 18028 10106 18040
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 10413 18031 10471 18037
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 12023 18040 12449 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12437 18037 12449 18040
rect 12483 18068 12495 18071
rect 12728 18068 12756 18167
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 14369 18139 14427 18145
rect 14369 18136 14381 18139
rect 13648 18108 14381 18136
rect 12894 18068 12900 18080
rect 12483 18040 12900 18068
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 13648 18068 13676 18108
rect 14369 18105 14381 18108
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 16025 18139 16083 18145
rect 16025 18105 16037 18139
rect 16071 18136 16083 18139
rect 16206 18136 16212 18148
rect 16071 18108 16212 18136
rect 16071 18105 16083 18108
rect 16025 18099 16083 18105
rect 16206 18096 16212 18108
rect 16264 18096 16270 18148
rect 13504 18040 13676 18068
rect 14093 18071 14151 18077
rect 13504 18028 13510 18040
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 14182 18068 14188 18080
rect 14139 18040 14188 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 17126 18068 17132 18080
rect 14332 18040 17132 18068
rect 14332 18028 14338 18040
rect 17126 18028 17132 18040
rect 17184 18068 17190 18080
rect 18325 18071 18383 18077
rect 18325 18068 18337 18071
rect 17184 18040 18337 18068
rect 17184 18028 17190 18040
rect 18325 18037 18337 18040
rect 18371 18037 18383 18071
rect 18325 18031 18383 18037
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 1728 17836 2513 17864
rect 1728 17824 1734 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 2501 17827 2559 17833
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3476 17836 4077 17864
rect 3476 17824 3482 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 5445 17867 5503 17873
rect 5445 17864 5457 17867
rect 4212 17836 5457 17864
rect 4212 17824 4218 17836
rect 5445 17833 5457 17836
rect 5491 17833 5503 17867
rect 5445 17827 5503 17833
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10318 17864 10324 17876
rect 9732 17836 10324 17864
rect 9732 17824 9738 17836
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11238 17864 11244 17876
rect 10827 17836 11244 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 17865 17867 17923 17873
rect 12115 17836 17816 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 3878 17756 3884 17808
rect 3936 17756 3942 17808
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 11057 17799 11115 17805
rect 11057 17796 11069 17799
rect 7248 17768 11069 17796
rect 7248 17756 7254 17768
rect 11057 17765 11069 17768
rect 11103 17765 11115 17799
rect 11057 17759 11115 17765
rect 11422 17756 11428 17808
rect 11480 17796 11486 17808
rect 12084 17796 12112 17827
rect 11480 17768 12112 17796
rect 17788 17796 17816 17836
rect 17865 17833 17877 17867
rect 17911 17864 17923 17867
rect 18046 17864 18052 17876
rect 17911 17836 18052 17864
rect 17911 17833 17923 17836
rect 17865 17827 17923 17833
rect 18046 17824 18052 17836
rect 18104 17864 18110 17876
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 18104 17836 18245 17864
rect 18104 17824 18110 17836
rect 18233 17833 18245 17836
rect 18279 17864 18291 17867
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18279 17836 18889 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18877 17833 18889 17836
rect 18923 17864 18935 17867
rect 19978 17864 19984 17876
rect 18923 17836 19984 17864
rect 18923 17833 18935 17836
rect 18877 17827 18935 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 19426 17796 19432 17808
rect 17788 17768 19432 17796
rect 11480 17756 11486 17768
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 19610 17796 19616 17808
rect 19571 17768 19616 17796
rect 19610 17756 19616 17768
rect 19668 17756 19674 17808
rect 3896 17728 3924 17756
rect 4062 17728 4068 17740
rect 3896 17700 4068 17728
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 4890 17728 4896 17740
rect 4755 17700 4896 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17728 6147 17731
rect 6822 17728 6828 17740
rect 6135 17700 6828 17728
rect 6135 17697 6147 17700
rect 6089 17691 6147 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 8202 17728 8208 17740
rect 8067 17700 8208 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9674 17728 9680 17740
rect 9631 17700 9680 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 14182 17728 14188 17740
rect 10091 17700 12434 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 1946 17660 1952 17672
rect 1907 17632 1952 17660
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2685 17663 2743 17669
rect 2685 17629 2697 17663
rect 2731 17660 2743 17663
rect 3878 17660 3884 17672
rect 2731 17632 3884 17660
rect 2731 17629 2743 17632
rect 2685 17623 2743 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4522 17660 4528 17672
rect 4479 17632 4528 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7524 17632 8340 17660
rect 7524 17620 7530 17632
rect 5813 17595 5871 17601
rect 5813 17561 5825 17595
rect 5859 17592 5871 17595
rect 6457 17595 6515 17601
rect 6457 17592 6469 17595
rect 5859 17564 6469 17592
rect 5859 17561 5871 17564
rect 5813 17555 5871 17561
rect 6457 17561 6469 17564
rect 6503 17561 6515 17595
rect 6457 17555 6515 17561
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 8205 17595 8263 17601
rect 8205 17592 8217 17595
rect 7340 17564 8217 17592
rect 7340 17552 7346 17564
rect 8205 17561 8217 17564
rect 8251 17561 8263 17595
rect 8312 17592 8340 17632
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9272 17632 9413 17660
rect 9272 17620 9278 17632
rect 9401 17629 9413 17632
rect 9447 17660 9459 17663
rect 10060 17660 10088 17691
rect 10594 17660 10600 17672
rect 9447 17632 10088 17660
rect 10555 17632 10600 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 12406 17660 12434 17700
rect 13648 17700 14188 17728
rect 13648 17660 13676 17700
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 19702 17728 19708 17740
rect 17184 17700 19708 17728
rect 17184 17688 17190 17700
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 12406 17632 13676 17660
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17660 13783 17663
rect 13998 17660 14004 17672
rect 13771 17632 14004 17660
rect 13771 17629 13783 17632
rect 13725 17623 13783 17629
rect 11422 17592 11428 17604
rect 8312 17564 11428 17592
rect 8205 17555 8263 17561
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 11790 17552 11796 17604
rect 11848 17592 11854 17604
rect 12158 17592 12164 17604
rect 11848 17564 12164 17592
rect 11848 17552 11854 17564
rect 12158 17552 12164 17564
rect 12216 17592 12222 17604
rect 13458 17595 13516 17601
rect 13458 17592 13470 17595
rect 12216 17564 13470 17592
rect 12216 17552 12222 17564
rect 13458 17561 13470 17564
rect 13504 17561 13516 17595
rect 13458 17555 13516 17561
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2130 17524 2136 17536
rect 2091 17496 2136 17524
rect 2130 17484 2136 17496
rect 2188 17484 2194 17536
rect 2406 17484 2412 17536
rect 2464 17524 2470 17536
rect 2682 17524 2688 17536
rect 2464 17496 2688 17524
rect 2464 17484 2470 17496
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3421 17527 3479 17533
rect 3421 17493 3433 17527
rect 3467 17524 3479 17527
rect 3602 17524 3608 17536
rect 3467 17496 3608 17524
rect 3467 17493 3479 17496
rect 3421 17487 3479 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 4580 17496 4625 17524
rect 4580 17484 4586 17496
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 4856 17496 5089 17524
rect 4856 17484 4862 17496
rect 5077 17493 5089 17496
rect 5123 17493 5135 17527
rect 5902 17524 5908 17536
rect 5863 17496 5908 17524
rect 5077 17487 5135 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6822 17524 6828 17536
rect 6420 17496 6828 17524
rect 6420 17484 6426 17496
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 7064 17496 7205 17524
rect 7064 17484 7070 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7984 17496 8125 17524
rect 7984 17484 7990 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8570 17524 8576 17536
rect 8531 17496 8576 17524
rect 8113 17487 8171 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 9088 17496 9321 17524
rect 9088 17484 9094 17496
rect 9309 17493 9321 17496
rect 9355 17493 9367 17527
rect 11698 17524 11704 17536
rect 11659 17496 11704 17524
rect 9309 17487 9367 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 12342 17524 12348 17536
rect 12303 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12894 17484 12900 17536
rect 12952 17524 12958 17536
rect 13740 17524 13768 17623
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 15470 17660 15476 17672
rect 15383 17632 15476 17660
rect 15470 17620 15476 17632
rect 15528 17660 15534 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15528 17632 15853 17660
rect 15528 17620 15534 17632
rect 15841 17629 15853 17632
rect 15887 17660 15899 17663
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15887 17632 16129 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 16117 17629 16129 17632
rect 16163 17660 16175 17663
rect 16206 17660 16212 17672
rect 16163 17632 16212 17660
rect 16163 17629 16175 17632
rect 16117 17623 16175 17629
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 21358 17660 21364 17672
rect 21319 17632 21364 17660
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 14918 17552 14924 17604
rect 14976 17592 14982 17604
rect 15206 17595 15264 17601
rect 15206 17592 15218 17595
rect 14976 17564 15218 17592
rect 14976 17552 14982 17564
rect 15206 17561 15218 17564
rect 15252 17561 15264 17595
rect 15206 17555 15264 17561
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 16362 17595 16420 17601
rect 16362 17592 16374 17595
rect 15620 17564 16374 17592
rect 15620 17552 15626 17564
rect 16362 17561 16374 17564
rect 16408 17561 16420 17595
rect 20806 17592 20812 17604
rect 16362 17555 16420 17561
rect 17512 17564 20812 17592
rect 17512 17536 17540 17564
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 20990 17552 20996 17604
rect 21048 17592 21054 17604
rect 21094 17595 21152 17601
rect 21094 17592 21106 17595
rect 21048 17564 21106 17592
rect 21048 17552 21054 17564
rect 21094 17561 21106 17564
rect 21140 17561 21152 17595
rect 21094 17555 21152 17561
rect 12952 17496 13768 17524
rect 14093 17527 14151 17533
rect 12952 17484 12958 17496
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 14366 17524 14372 17536
rect 14139 17496 14372 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 19334 17524 19340 17536
rect 17736 17496 19340 17524
rect 17736 17484 17742 17496
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 19518 17484 19524 17536
rect 19576 17524 19582 17536
rect 19981 17527 20039 17533
rect 19981 17524 19993 17527
rect 19576 17496 19993 17524
rect 19576 17484 19582 17496
rect 19981 17493 19993 17496
rect 20027 17493 20039 17527
rect 19981 17487 20039 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2314 17280 2320 17332
rect 2372 17320 2378 17332
rect 2777 17323 2835 17329
rect 2777 17320 2789 17323
rect 2372 17292 2789 17320
rect 2372 17280 2378 17292
rect 2777 17289 2789 17292
rect 2823 17289 2835 17323
rect 3234 17320 3240 17332
rect 3195 17292 3240 17320
rect 2777 17283 2835 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 3602 17320 3608 17332
rect 3563 17292 3608 17320
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 4522 17320 4528 17332
rect 4483 17292 4528 17320
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 4890 17280 4896 17332
rect 4948 17280 4954 17332
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5350 17320 5356 17332
rect 5031 17292 5356 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 5960 17292 6377 17320
rect 5960 17280 5966 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6604 17292 6837 17320
rect 6604 17280 6610 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 6825 17283 6883 17289
rect 7561 17323 7619 17329
rect 7561 17289 7573 17323
rect 7607 17320 7619 17323
rect 7650 17320 7656 17332
rect 7607 17292 7656 17320
rect 7607 17289 7619 17292
rect 7561 17283 7619 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 8021 17323 8079 17329
rect 8021 17289 8033 17323
rect 8067 17320 8079 17323
rect 8938 17320 8944 17332
rect 8067 17292 8944 17320
rect 8067 17289 8079 17292
rect 8021 17283 8079 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 9861 17323 9919 17329
rect 9861 17320 9873 17323
rect 9732 17292 9873 17320
rect 9732 17280 9738 17292
rect 9861 17289 9873 17292
rect 9907 17289 9919 17323
rect 9861 17283 9919 17289
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11238 17320 11244 17332
rect 11103 17292 11244 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 11609 17323 11667 17329
rect 11609 17289 11621 17323
rect 11655 17320 11667 17323
rect 11698 17320 11704 17332
rect 11655 17292 11704 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 11698 17280 11704 17292
rect 11756 17320 11762 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 11756 17292 11989 17320
rect 11756 17280 11762 17292
rect 11977 17289 11989 17292
rect 12023 17320 12035 17323
rect 12894 17320 12900 17332
rect 12023 17292 12900 17320
rect 12023 17289 12035 17292
rect 11977 17283 12035 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13814 17320 13820 17332
rect 13320 17292 13820 17320
rect 13320 17280 13326 17292
rect 2501 17255 2559 17261
rect 2501 17221 2513 17255
rect 2547 17252 2559 17255
rect 4908 17252 4936 17280
rect 13381 17261 13409 17292
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 14056 17292 14381 17320
rect 14056 17280 14062 17292
rect 14369 17289 14381 17292
rect 14415 17320 14427 17323
rect 14737 17323 14795 17329
rect 14737 17320 14749 17323
rect 14415 17292 14749 17320
rect 14415 17289 14427 17292
rect 14369 17283 14427 17289
rect 14737 17289 14749 17292
rect 14783 17320 14795 17323
rect 15470 17320 15476 17332
rect 14783 17292 15476 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 16316 17292 18276 17320
rect 2547 17224 4936 17252
rect 7929 17255 7987 17261
rect 2547 17221 2559 17224
rect 2501 17215 2559 17221
rect 7929 17221 7941 17255
rect 7975 17252 7987 17255
rect 9401 17255 9459 17261
rect 9401 17252 9413 17255
rect 7975 17224 9413 17252
rect 7975 17221 7987 17224
rect 7929 17215 7987 17221
rect 9401 17221 9413 17224
rect 9447 17221 9459 17255
rect 9401 17215 9459 17221
rect 13366 17255 13424 17261
rect 13366 17221 13378 17255
rect 13412 17221 13424 17255
rect 13366 17215 13424 17221
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 13964 17224 14136 17252
rect 13964 17212 13970 17224
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 1762 17184 1768 17196
rect 1719 17156 1768 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2866 17184 2872 17196
rect 2179 17156 2872 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 4154 17184 4160 17196
rect 3007 17156 4160 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4522 17144 4528 17196
rect 4580 17184 4586 17196
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4580 17156 4905 17184
rect 4580 17144 4586 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 4893 17147 4951 17153
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 3384 17088 3709 17116
rect 3384 17076 3390 17088
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 3844 17088 3937 17116
rect 3844 17076 3850 17088
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 3804 17048 3832 17076
rect 3016 17020 3832 17048
rect 3016 17008 3022 17020
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 4908 16980 4936 17147
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6822 17184 6828 17196
rect 6779 17156 6828 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8628 17156 8953 17184
rect 8628 17144 8634 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10502 17184 10508 17196
rect 10367 17156 10508 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10502 17144 10508 17156
rect 10560 17184 10566 17196
rect 13626 17187 13684 17193
rect 10560 17156 13584 17184
rect 10560 17144 10566 17156
rect 5166 17116 5172 17128
rect 5127 17088 5172 17116
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 5718 17076 5724 17128
rect 5776 17116 5782 17128
rect 6546 17116 6552 17128
rect 5776 17088 6552 17116
rect 5776 17076 5782 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 7006 17116 7012 17128
rect 6919 17088 7012 17116
rect 7006 17076 7012 17088
rect 7064 17116 7070 17128
rect 7064 17088 7328 17116
rect 7064 17076 7070 17088
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 6638 17048 6644 17060
rect 6043 17020 6644 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 6638 17008 6644 17020
rect 6696 17008 6702 17060
rect 5166 16980 5172 16992
rect 4908 16952 5172 16980
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 7300 16980 7328 17088
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 8205 17119 8263 17125
rect 8205 17116 8217 17119
rect 7616 17088 8217 17116
rect 7616 17076 7622 17088
rect 8205 17085 8217 17088
rect 8251 17116 8263 17119
rect 8665 17119 8723 17125
rect 8665 17116 8677 17119
rect 8251 17088 8677 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8665 17085 8677 17088
rect 8711 17085 8723 17119
rect 13556 17116 13584 17156
rect 13626 17153 13638 17187
rect 13672 17184 13684 17187
rect 13998 17184 14004 17196
rect 13672 17156 14004 17184
rect 13672 17153 13684 17156
rect 13626 17147 13684 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14108 17184 14136 17224
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 16316 17252 16344 17292
rect 14240 17224 16344 17252
rect 14240 17212 14246 17224
rect 16390 17212 16396 17264
rect 16448 17252 16454 17264
rect 17313 17255 17371 17261
rect 17313 17252 17325 17255
rect 16448 17224 17325 17252
rect 16448 17212 16454 17224
rect 17313 17221 17325 17224
rect 17359 17252 17371 17255
rect 18046 17252 18052 17264
rect 17359 17224 18052 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17034 17184 17040 17196
rect 14108 17156 17040 17184
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17604 17193 17632 17224
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 17678 17144 17684 17196
rect 17736 17144 17742 17196
rect 17856 17187 17914 17193
rect 17856 17153 17868 17187
rect 17902 17184 17914 17187
rect 18138 17184 18144 17196
rect 17902 17156 18144 17184
rect 17902 17153 17914 17156
rect 17856 17147 17914 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18248 17184 18276 17292
rect 19058 17280 19064 17332
rect 19116 17320 19122 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 19116 17292 19349 17320
rect 19116 17280 19122 17292
rect 19337 17289 19349 17292
rect 19383 17320 19395 17323
rect 19978 17320 19984 17332
rect 19383 17292 19984 17320
rect 19383 17289 19395 17292
rect 19337 17283 19395 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20990 17212 20996 17264
rect 21048 17252 21054 17264
rect 21094 17255 21152 17261
rect 21094 17252 21106 17255
rect 21048 17224 21106 17252
rect 21048 17212 21054 17224
rect 21094 17221 21106 17224
rect 21140 17221 21152 17255
rect 21094 17215 21152 17221
rect 19794 17184 19800 17196
rect 18248 17156 19800 17184
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 21358 17184 21364 17196
rect 21319 17156 21364 17184
rect 21358 17144 21364 17156
rect 21416 17144 21422 17196
rect 17696 17116 17724 17144
rect 13556 17088 17724 17116
rect 8665 17079 8723 17085
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 7432 17020 10609 17048
rect 7432 17008 7438 17020
rect 10597 17017 10609 17020
rect 10643 17017 10655 17051
rect 10597 17011 10655 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 10836 17020 12265 17048
rect 10836 17008 10842 17020
rect 12253 17017 12265 17020
rect 12299 17017 12311 17051
rect 12253 17011 12311 17017
rect 11238 16980 11244 16992
rect 7300 16952 11244 16980
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12268 16980 12296 17011
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 15194 17048 15200 17060
rect 13780 17020 15200 17048
rect 13780 17008 13786 17020
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 15396 17020 17632 17048
rect 15396 16992 15424 17020
rect 13814 16980 13820 16992
rect 12268 16952 13820 16980
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 15289 16983 15347 16989
rect 15289 16949 15301 16983
rect 15335 16980 15347 16983
rect 15378 16980 15384 16992
rect 15335 16952 15384 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15528 16952 15669 16980
rect 15528 16940 15534 16952
rect 15657 16949 15669 16952
rect 15703 16980 15715 16983
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15703 16952 16313 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 16301 16949 16313 16952
rect 16347 16980 16359 16983
rect 16390 16980 16396 16992
rect 16347 16952 16396 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17604 16980 17632 17020
rect 19334 17008 19340 17060
rect 19392 17048 19398 17060
rect 20346 17048 20352 17060
rect 19392 17020 20352 17048
rect 19392 17008 19398 17020
rect 20346 17008 20352 17020
rect 20404 17008 20410 17060
rect 17954 16980 17960 16992
rect 17604 16952 17960 16980
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18966 16980 18972 16992
rect 18927 16952 18972 16980
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19702 16980 19708 16992
rect 19663 16952 19708 16980
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 19981 16983 20039 16989
rect 19981 16980 19993 16983
rect 19944 16952 19993 16980
rect 19944 16940 19950 16952
rect 19981 16949 19993 16952
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 2409 16779 2467 16785
rect 2409 16776 2421 16779
rect 1728 16748 2421 16776
rect 1728 16736 1734 16748
rect 2409 16745 2421 16748
rect 2455 16745 2467 16779
rect 2409 16739 2467 16745
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 2924 16748 3249 16776
rect 2924 16736 2930 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 4154 16776 4160 16788
rect 4115 16748 4160 16776
rect 3237 16739 3295 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5132 16748 7236 16776
rect 5132 16736 5138 16748
rect 2961 16711 3019 16717
rect 2961 16677 2973 16711
rect 3007 16708 3019 16711
rect 4522 16708 4528 16720
rect 3007 16680 4528 16708
rect 3007 16677 3019 16680
rect 2961 16671 3019 16677
rect 4522 16668 4528 16680
rect 4580 16668 4586 16720
rect 5994 16708 6000 16720
rect 4632 16680 6000 16708
rect 4632 16649 4660 16680
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7208 16708 7236 16748
rect 7834 16736 7840 16788
rect 7892 16776 7898 16788
rect 8754 16776 8760 16788
rect 7892 16748 8760 16776
rect 7892 16736 7898 16748
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 20070 16776 20076 16788
rect 11072 16748 20076 16776
rect 7208 16680 7328 16708
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16609 4675 16643
rect 4798 16640 4804 16652
rect 4759 16612 4804 16640
rect 4617 16603 4675 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 7190 16640 7196 16652
rect 7151 16612 7196 16640
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 1946 16572 1952 16584
rect 1719 16544 1952 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16572 2651 16575
rect 2774 16572 2780 16584
rect 2639 16544 2780 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 2148 16504 2176 16535
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3467 16544 5856 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3234 16504 3240 16516
rect 2148 16476 3240 16504
rect 3234 16464 3240 16476
rect 3292 16464 3298 16516
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16504 4583 16507
rect 5169 16507 5227 16513
rect 5169 16504 5181 16507
rect 4571 16476 5181 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 5169 16473 5181 16476
rect 5215 16473 5227 16507
rect 5169 16467 5227 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1912 16408 1961 16436
rect 1912 16396 1918 16408
rect 1949 16405 1961 16408
rect 1995 16405 2007 16439
rect 1949 16399 2007 16405
rect 3881 16439 3939 16445
rect 3881 16405 3893 16439
rect 3927 16436 3939 16439
rect 4062 16436 4068 16448
rect 3927 16408 4068 16436
rect 3927 16405 3939 16408
rect 3881 16399 3939 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5828 16436 5856 16544
rect 6273 16507 6331 16513
rect 6273 16473 6285 16507
rect 6319 16504 6331 16507
rect 6917 16507 6975 16513
rect 6917 16504 6929 16507
rect 6319 16476 6929 16504
rect 6319 16473 6331 16476
rect 6273 16467 6331 16473
rect 6917 16473 6929 16476
rect 6963 16473 6975 16507
rect 6917 16467 6975 16473
rect 6549 16439 6607 16445
rect 6549 16436 6561 16439
rect 5828 16408 6561 16436
rect 6549 16405 6561 16408
rect 6595 16405 6607 16439
rect 6549 16399 6607 16405
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7098 16436 7104 16448
rect 7055 16408 7104 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 7300 16436 7328 16680
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 7929 16643 7987 16649
rect 7929 16640 7941 16643
rect 7892 16612 7941 16640
rect 7892 16600 7898 16612
rect 7929 16609 7941 16612
rect 7975 16609 7987 16643
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 7929 16603 7987 16609
rect 8036 16612 8953 16640
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 8036 16572 8064 16612
rect 7432 16544 8064 16572
rect 7432 16532 7438 16544
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 8220 16581 8248 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 11072 16649 11100 16748
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 12069 16711 12127 16717
rect 12069 16708 12081 16711
rect 11164 16680 12081 16708
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 9180 16612 10977 16640
rect 9180 16600 9186 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 8205 16535 8263 16541
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 8128 16504 8156 16532
rect 8128 16476 8616 16504
rect 8588 16445 8616 16476
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11164 16504 11192 16680
rect 12069 16677 12081 16680
rect 12115 16708 12127 16711
rect 12158 16708 12164 16720
rect 12115 16680 12164 16708
rect 12115 16677 12127 16680
rect 12069 16671 12127 16677
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12391 16612 12480 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12452 16572 12480 16612
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15528 16612 15761 16640
rect 15528 16600 15534 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16640 18935 16643
rect 19058 16640 19064 16652
rect 18923 16612 19064 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 19058 16600 19064 16612
rect 19116 16640 19122 16652
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 19116 16612 19441 16640
rect 19116 16600 19122 16612
rect 19429 16609 19441 16612
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 12452 16544 14105 16572
rect 14093 16541 14105 16544
rect 14139 16572 14151 16575
rect 15488 16572 15516 16600
rect 19702 16581 19708 16584
rect 19685 16575 19708 16581
rect 19685 16572 19697 16575
rect 14139 16544 15516 16572
rect 15948 16544 19697 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 12590 16507 12648 16513
rect 12590 16504 12602 16507
rect 11020 16476 11192 16504
rect 12406 16476 12602 16504
rect 11020 16464 11026 16476
rect 12406 16448 12434 16476
rect 12590 16473 12602 16476
rect 12636 16473 12648 16507
rect 12590 16467 12648 16473
rect 13814 16464 13820 16516
rect 13872 16504 13878 16516
rect 14338 16507 14396 16513
rect 14338 16504 14350 16507
rect 13872 16476 14350 16504
rect 13872 16464 13878 16476
rect 14338 16473 14350 16476
rect 14384 16473 14396 16507
rect 15948 16504 15976 16544
rect 19685 16541 19697 16544
rect 19760 16572 19766 16584
rect 21082 16572 21088 16584
rect 19760 16544 19833 16572
rect 21043 16544 21088 16572
rect 19685 16535 19708 16541
rect 19702 16532 19708 16535
rect 19760 16532 19766 16544
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 16022 16513 16028 16516
rect 14338 16467 14396 16473
rect 15396 16476 15976 16504
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7300 16408 8125 16436
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 8573 16439 8631 16445
rect 8573 16405 8585 16439
rect 8619 16405 8631 16439
rect 9582 16436 9588 16448
rect 9543 16408 9588 16436
rect 8573 16399 8631 16405
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 10226 16436 10232 16448
rect 10187 16408 10232 16436
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10376 16408 10517 16436
rect 10376 16396 10382 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10870 16436 10876 16448
rect 10831 16408 10876 16436
rect 10505 16399 10563 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11882 16436 11888 16448
rect 11747 16408 11888 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12342 16396 12348 16448
rect 12400 16408 12434 16448
rect 12400 16396 12406 16408
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13596 16408 13737 16436
rect 13596 16396 13602 16408
rect 13725 16405 13737 16408
rect 13771 16436 13783 16439
rect 15396 16436 15424 16476
rect 16016 16467 16028 16513
rect 16080 16504 16086 16516
rect 17218 16504 17224 16516
rect 16080 16476 16116 16504
rect 17131 16476 17224 16504
rect 16022 16464 16028 16467
rect 16080 16464 16086 16476
rect 13771 16408 15424 16436
rect 15473 16439 15531 16445
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 15654 16436 15660 16448
rect 15519 16408 15660 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 17144 16445 17172 16476
rect 17218 16464 17224 16476
rect 17276 16504 17282 16516
rect 17276 16476 18184 16504
rect 17276 16464 17282 16476
rect 17129 16439 17187 16445
rect 17129 16405 17141 16439
rect 17175 16405 17187 16439
rect 17494 16436 17500 16448
rect 17455 16408 17500 16436
rect 17129 16399 17187 16405
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 18156 16436 18184 16476
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 18610 16507 18668 16513
rect 18610 16504 18622 16507
rect 18288 16476 18622 16504
rect 18288 16464 18294 16476
rect 18610 16473 18622 16476
rect 18656 16473 18668 16507
rect 20990 16504 20996 16516
rect 18610 16467 18668 16473
rect 18708 16476 20996 16504
rect 18708 16436 18736 16476
rect 20990 16464 20996 16476
rect 21048 16464 21054 16516
rect 20806 16436 20812 16448
rect 18156 16408 18736 16436
rect 20767 16408 20812 16436
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21269 16439 21327 16445
rect 21269 16436 21281 16439
rect 20956 16408 21281 16436
rect 20956 16396 20962 16408
rect 21269 16405 21281 16408
rect 21315 16405 21327 16439
rect 21269 16399 21327 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 3326 16232 3332 16244
rect 2832 16204 2877 16232
rect 3287 16204 3332 16232
rect 2832 16192 2838 16204
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 3970 16232 3976 16244
rect 3835 16204 3976 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 5534 16232 5540 16244
rect 5495 16204 5540 16232
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 6052 16204 6377 16232
rect 6052 16192 6058 16204
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 6365 16195 6423 16201
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7006 16232 7012 16244
rect 6788 16204 7012 16232
rect 6788 16192 6794 16204
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7377 16235 7435 16241
rect 7377 16232 7389 16235
rect 7248 16204 7389 16232
rect 7248 16192 7254 16204
rect 7377 16201 7389 16204
rect 7423 16201 7435 16235
rect 7926 16232 7932 16244
rect 7887 16204 7932 16232
rect 7377 16195 7435 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8343 16204 9045 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 9033 16201 9045 16204
rect 9079 16232 9091 16235
rect 9214 16232 9220 16244
rect 9079 16204 9220 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10870 16232 10876 16244
rect 10831 16204 10876 16232
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 15289 16235 15347 16241
rect 12406 16204 15240 16232
rect 6822 16164 6828 16176
rect 2976 16136 6828 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2976 16105 3004 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 8018 16124 8024 16176
rect 8076 16164 8082 16176
rect 8076 16136 12112 16164
rect 8076 16124 8082 16136
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3326 16056 3332 16108
rect 3384 16096 3390 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3384 16068 3709 16096
rect 3384 16056 3390 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 4522 16096 4528 16108
rect 4483 16068 4528 16096
rect 3697 16059 3755 16065
rect 4522 16056 4528 16068
rect 4580 16056 4586 16108
rect 5445 16099 5503 16105
rect 5445 16065 5457 16099
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 16028 4031 16031
rect 4062 16028 4068 16040
rect 4019 16000 4068 16028
rect 4019 15997 4031 16000
rect 3973 15991 4031 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 5074 16028 5080 16040
rect 4212 16000 5080 16028
rect 4212 15988 4218 16000
rect 5074 15988 5080 16000
rect 5132 16028 5138 16040
rect 5460 16028 5488 16059
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 5776 16068 6745 16096
rect 5776 16056 5782 16068
rect 6733 16065 6745 16068
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 5132 16000 5488 16028
rect 5629 16031 5687 16037
rect 5132 15988 5138 16000
rect 5629 15997 5641 16031
rect 5675 15997 5687 16031
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 5629 15991 5687 15997
rect 5920 16000 6837 16028
rect 2038 15960 2044 15972
rect 1999 15932 2044 15960
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 3878 15920 3884 15972
rect 3936 15960 3942 15972
rect 4341 15963 4399 15969
rect 4341 15960 4353 15963
rect 3936 15932 4353 15960
rect 3936 15920 3942 15932
rect 4341 15929 4353 15932
rect 4387 15929 4399 15963
rect 4341 15923 4399 15929
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 5644 15960 5672 15991
rect 5500 15932 5672 15960
rect 5500 15920 5506 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 5040 15864 5089 15892
rect 5040 15852 5046 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 5077 15855 5135 15861
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 5920 15892 5948 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 6825 15991 6883 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 5994 15920 6000 15972
rect 6052 15960 6058 15972
rect 7576 15960 7604 16059
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 8168 16068 8401 16096
rect 8168 16056 8174 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 8662 16056 8668 16108
rect 8720 16096 8726 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 8720 16068 9321 16096
rect 8720 16056 8726 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 10318 16096 10324 16108
rect 10279 16068 10324 16096
rect 9309 16059 9367 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 8570 16028 8576 16040
rect 8531 16000 8576 16028
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 6052 15932 7604 15960
rect 6052 15920 6058 15932
rect 7650 15920 7656 15972
rect 7708 15960 7714 15972
rect 11992 15960 12020 15991
rect 7708 15932 12020 15960
rect 12084 15960 12112 16136
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 16028 12219 16031
rect 12406 16028 12434 16204
rect 14308 16167 14366 16173
rect 14308 16133 14320 16167
rect 14354 16164 14366 16167
rect 15102 16164 15108 16176
rect 14354 16136 15108 16164
rect 14354 16133 14366 16136
rect 14308 16127 14366 16133
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 15212 16164 15240 16204
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15470 16232 15476 16244
rect 15335 16204 15476 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 16298 16232 16304 16244
rect 16259 16204 16304 16232
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 20717 16235 20775 16241
rect 20717 16232 20729 16235
rect 20404 16204 20729 16232
rect 20404 16192 20410 16204
rect 20717 16201 20729 16204
rect 20763 16201 20775 16235
rect 20717 16195 20775 16201
rect 17402 16164 17408 16176
rect 15212 16136 17408 16164
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 19306 16167 19364 16173
rect 19306 16164 19318 16167
rect 19024 16136 19318 16164
rect 19024 16124 19030 16136
rect 19306 16133 19318 16136
rect 19352 16133 19364 16167
rect 19306 16127 19364 16133
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 12986 16096 12992 16108
rect 12943 16068 12992 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 15470 16096 15476 16108
rect 14599 16068 15476 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 17494 16096 17500 16108
rect 17052 16068 17500 16096
rect 12207 16000 12434 16028
rect 12207 15997 12219 16000
rect 12161 15991 12219 15997
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 17052 16028 17080 16068
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 17770 16056 17776 16108
rect 17828 16105 17834 16108
rect 17828 16096 17840 16105
rect 18049 16099 18107 16105
rect 17828 16068 18000 16096
rect 17828 16059 17840 16068
rect 17828 16056 17834 16059
rect 15068 16000 17080 16028
rect 17972 16028 18000 16068
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18417 16099 18475 16105
rect 18417 16096 18429 16099
rect 18095 16068 18429 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18417 16065 18429 16068
rect 18463 16096 18475 16099
rect 19058 16096 19064 16108
rect 18463 16068 19064 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19886 16096 19892 16108
rect 19168 16068 19892 16096
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 17972 16000 18705 16028
rect 15068 15988 15074 16000
rect 18693 15997 18705 16000
rect 18739 16028 18751 16031
rect 19168 16028 19196 16068
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 18739 16000 19196 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 13538 15960 13544 15972
rect 12084 15932 13544 15960
rect 7708 15920 7714 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 16022 15960 16028 15972
rect 14752 15932 16028 15960
rect 5684 15864 5948 15892
rect 5684 15852 5690 15864
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 6144 15864 9689 15892
rect 6144 15852 6150 15864
rect 9677 15861 9689 15864
rect 9723 15861 9735 15895
rect 9677 15855 9735 15861
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 10468 15864 11529 15892
rect 10468 15852 10474 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 13170 15892 13176 15904
rect 13131 15864 13176 15892
rect 11517 15855 11575 15861
rect 13170 15852 13176 15864
rect 13228 15892 13234 15904
rect 14752 15892 14780 15932
rect 16022 15920 16028 15932
rect 16080 15920 16086 15972
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 21140 15932 21189 15960
rect 21140 15920 21146 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21177 15923 21235 15929
rect 13228 15864 14780 15892
rect 13228 15852 13234 15864
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 14884 15864 14929 15892
rect 14884 15852 14890 15864
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 15565 15895 15623 15901
rect 15565 15892 15577 15895
rect 15160 15864 15577 15892
rect 15160 15852 15166 15864
rect 15565 15861 15577 15864
rect 15611 15861 15623 15895
rect 15565 15855 15623 15861
rect 15930 15852 15936 15904
rect 15988 15892 15994 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 15988 15864 16681 15892
rect 15988 15852 15994 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20441 15895 20499 15901
rect 20441 15892 20453 15895
rect 20036 15864 20453 15892
rect 20036 15852 20042 15864
rect 20441 15861 20453 15864
rect 20487 15861 20499 15895
rect 20441 15855 20499 15861
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2648 15660 2881 15688
rect 2648 15648 2654 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 2869 15651 2927 15657
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3510 15688 3516 15700
rect 3384 15660 3516 15688
rect 3384 15648 3390 15660
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 6086 15688 6092 15700
rect 4672 15660 6092 15688
rect 4672 15648 4678 15660
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7650 15688 7656 15700
rect 7423 15660 7656 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 8202 15688 8208 15700
rect 7760 15660 8208 15688
rect 1762 15580 1768 15632
rect 1820 15620 1826 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 1820 15592 2421 15620
rect 1820 15580 1826 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 7760 15620 7788 15660
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15688 8631 15691
rect 9398 15688 9404 15700
rect 8619 15660 9404 15688
rect 8619 15657 8631 15660
rect 8573 15651 8631 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 9732 15660 10241 15688
rect 9732 15648 9738 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10229 15651 10287 15657
rect 12989 15691 13047 15697
rect 12989 15657 13001 15691
rect 13035 15688 13047 15691
rect 20714 15688 20720 15700
rect 13035 15660 20720 15688
rect 13035 15657 13047 15660
rect 12989 15651 13047 15657
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 13446 15620 13452 15632
rect 5500 15592 7788 15620
rect 8036 15592 13452 15620
rect 5500 15580 5506 15592
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5626 15552 5632 15564
rect 4847 15524 5632 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 6288 15561 6316 15592
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 7190 15552 7196 15564
rect 6871 15524 7196 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 8036 15561 8064 15592
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 15473 15623 15531 15629
rect 15473 15589 15485 15623
rect 15519 15620 15531 15623
rect 15562 15620 15568 15632
rect 15519 15592 15568 15620
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 18509 15623 18567 15629
rect 18509 15589 18521 15623
rect 18555 15620 18567 15623
rect 18874 15620 18880 15632
rect 18555 15592 18880 15620
rect 18555 15589 18567 15592
rect 18509 15583 18567 15589
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 8352 15524 11253 15552
rect 8352 15512 8358 15524
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 11425 15555 11483 15561
rect 11425 15521 11437 15555
rect 11471 15552 11483 15555
rect 11471 15524 12434 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 1854 15484 1860 15496
rect 1719 15456 1860 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2133 15487 2191 15493
rect 2133 15484 2145 15487
rect 2004 15456 2145 15484
rect 2004 15444 2010 15456
rect 2133 15453 2145 15456
rect 2179 15453 2191 15487
rect 2590 15484 2596 15496
rect 2551 15456 2596 15484
rect 2133 15447 2191 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3418 15484 3424 15496
rect 3099 15456 3424 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5534 15444 5540 15496
rect 5592 15484 5598 15496
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 5592 15456 6929 15484
rect 5592 15444 5598 15456
rect 6917 15453 6929 15456
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 10410 15484 10416 15496
rect 8628 15456 10272 15484
rect 10371 15456 10416 15484
rect 8628 15444 8634 15456
rect 4154 15416 4160 15428
rect 4115 15388 4160 15416
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 4893 15419 4951 15425
rect 4893 15385 4905 15419
rect 4939 15416 4951 15419
rect 5997 15419 6055 15425
rect 4939 15388 5672 15416
rect 4939 15385 4951 15388
rect 4893 15379 4951 15385
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 3421 15351 3479 15357
rect 3421 15317 3433 15351
rect 3467 15348 3479 15351
rect 3510 15348 3516 15360
rect 3467 15320 3516 15348
rect 3467 15317 3479 15320
rect 3421 15311 3479 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15348 5411 15351
rect 5442 15348 5448 15360
rect 5399 15320 5448 15348
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5644 15357 5672 15388
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 6730 15416 6736 15428
rect 6043 15388 6736 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 7834 15416 7840 15428
rect 6840 15388 7840 15416
rect 5629 15351 5687 15357
rect 5629 15317 5641 15351
rect 5675 15317 5687 15351
rect 5629 15311 5687 15317
rect 6089 15351 6147 15357
rect 6089 15317 6101 15351
rect 6135 15348 6147 15351
rect 6840 15348 6868 15388
rect 7834 15376 7840 15388
rect 7892 15416 7898 15428
rect 8128 15416 8156 15444
rect 7892 15388 8156 15416
rect 8205 15419 8263 15425
rect 7892 15376 7898 15388
rect 8205 15385 8217 15419
rect 8251 15416 8263 15419
rect 8662 15416 8668 15428
rect 8251 15388 8668 15416
rect 8251 15385 8263 15388
rect 8205 15379 8263 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 8941 15419 8999 15425
rect 8941 15416 8953 15419
rect 8812 15388 8953 15416
rect 8812 15376 8818 15388
rect 8941 15385 8953 15388
rect 8987 15385 8999 15419
rect 8941 15379 8999 15385
rect 9401 15419 9459 15425
rect 9401 15385 9413 15419
rect 9447 15416 9459 15419
rect 9490 15416 9496 15428
rect 9447 15388 9496 15416
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 10244 15416 10272 15456
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 11149 15419 11207 15425
rect 10244 15388 10916 15416
rect 6135 15320 6868 15348
rect 6135 15317 6147 15320
rect 6089 15311 6147 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 8110 15348 8116 15360
rect 7064 15320 7109 15348
rect 8071 15320 8116 15348
rect 7064 15308 7070 15320
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 10318 15348 10324 15360
rect 9815 15320 10324 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10560 15320 10793 15348
rect 10560 15308 10566 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10888 15348 10916 15388
rect 11149 15385 11161 15419
rect 11195 15416 11207 15419
rect 11793 15419 11851 15425
rect 11793 15416 11805 15419
rect 11195 15388 11805 15416
rect 11195 15385 11207 15388
rect 11149 15379 11207 15385
rect 11793 15385 11805 15388
rect 11839 15385 11851 15419
rect 12406 15416 12434 15524
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13403 15456 13737 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13725 15453 13737 15456
rect 13771 15484 13783 15487
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13771 15456 14105 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14093 15453 14105 15456
rect 14139 15484 14151 15487
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 14139 15456 15853 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 15841 15453 15853 15456
rect 15887 15484 15899 15487
rect 16298 15484 16304 15496
rect 15887 15456 16304 15484
rect 15887 15453 15899 15456
rect 15841 15447 15899 15453
rect 16298 15444 16304 15456
rect 16356 15484 16362 15496
rect 16485 15487 16543 15493
rect 16485 15484 16497 15487
rect 16356 15456 16497 15484
rect 16356 15444 16362 15456
rect 16485 15453 16497 15456
rect 16531 15484 16543 15487
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16531 15456 16773 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 16761 15453 16773 15456
rect 16807 15484 16819 15487
rect 18524 15484 18552 15583
rect 18874 15580 18880 15592
rect 18932 15620 18938 15632
rect 19058 15620 19064 15632
rect 18932 15592 19064 15620
rect 18932 15580 18938 15592
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 21358 15552 21364 15564
rect 21319 15524 21364 15552
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 16807 15456 18552 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 14182 15416 14188 15428
rect 12406 15388 14188 15416
rect 11793 15379 11851 15385
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 14360 15419 14418 15425
rect 14360 15385 14372 15419
rect 14406 15416 14418 15419
rect 15010 15416 15016 15428
rect 14406 15388 15016 15416
rect 14406 15385 14418 15388
rect 14360 15379 14418 15385
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 17006 15419 17064 15425
rect 17006 15416 17018 15419
rect 16448 15388 17018 15416
rect 16448 15376 16454 15388
rect 17006 15385 17018 15388
rect 17052 15385 17064 15419
rect 17006 15379 17064 15385
rect 20806 15376 20812 15428
rect 20864 15416 20870 15428
rect 21082 15416 21088 15428
rect 21140 15425 21146 15428
rect 20864 15388 21088 15416
rect 20864 15376 20870 15388
rect 21082 15376 21088 15388
rect 21140 15416 21152 15425
rect 21140 15388 21185 15416
rect 21140 15379 21152 15388
rect 21140 15376 21146 15379
rect 15562 15348 15568 15360
rect 10888 15320 15568 15348
rect 10781 15311 10839 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 18138 15348 18144 15360
rect 18099 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 18966 15348 18972 15360
rect 18656 15320 18972 15348
rect 18656 15308 18662 15320
rect 18966 15308 18972 15320
rect 19024 15348 19030 15360
rect 19337 15351 19395 15357
rect 19337 15348 19349 15351
rect 19024 15320 19349 15348
rect 19024 15308 19030 15320
rect 19337 15317 19349 15320
rect 19383 15317 19395 15351
rect 19702 15348 19708 15360
rect 19663 15320 19708 15348
rect 19337 15311 19395 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1728 15116 1961 15144
rect 1728 15104 1734 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 2590 15144 2596 15156
rect 2551 15116 2596 15144
rect 1949 15107 2007 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 2958 15144 2964 15156
rect 2919 15116 2964 15144
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 4019 15116 5549 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 5994 15144 6000 15156
rect 5955 15116 6000 15144
rect 5537 15107 5595 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 6914 15144 6920 15156
rect 6788 15116 6920 15144
rect 6788 15104 6794 15116
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7156 15116 7849 15144
rect 7156 15104 7162 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 9916 15116 10333 15144
rect 9916 15104 9922 15116
rect 10321 15113 10333 15116
rect 10367 15113 10379 15147
rect 10321 15107 10379 15113
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 4154 15076 4160 15088
rect 3436 15048 4160 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1762 15008 1768 15020
rect 1719 14980 1768 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2406 15008 2412 15020
rect 2367 14980 2412 15008
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 3436 14949 3464 15048
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 4525 15079 4583 15085
rect 4525 15045 4537 15079
rect 4571 15076 4583 15079
rect 4706 15076 4712 15088
rect 4571 15048 4712 15076
rect 4571 15045 4583 15048
rect 4525 15039 4583 15045
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 5000 15048 7328 15076
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3878 15008 3884 15020
rect 3651 14980 3884 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 3970 14940 3976 14952
rect 3559 14912 3976 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4430 14940 4436 14952
rect 4391 14912 4436 14940
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 2590 14832 2596 14884
rect 2648 14872 2654 14884
rect 4632 14872 4660 14971
rect 5000 14881 5028 15048
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 7190 15008 7196 15020
rect 5675 14980 5948 15008
rect 7151 14980 7196 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5920 14952 5948 14980
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5534 14940 5540 14952
rect 5399 14912 5540 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5902 14900 5908 14952
rect 5960 14900 5966 14952
rect 6914 14940 6920 14952
rect 6875 14912 6920 14940
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7300 14940 7328 15048
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 7800 15048 8309 15076
rect 7800 15036 7806 15048
rect 8297 15045 8309 15048
rect 8343 15045 8355 15079
rect 8297 15039 8355 15045
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 10796 15076 10824 15107
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 14182 15144 14188 15156
rect 10928 15116 14188 15144
rect 10928 15104 10934 15116
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 14550 15144 14556 15156
rect 14463 15116 14556 15144
rect 14550 15104 14556 15116
rect 14608 15144 14614 15156
rect 17494 15144 17500 15156
rect 14608 15116 17500 15144
rect 14608 15104 14614 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 19426 15144 19432 15156
rect 17972 15116 19432 15144
rect 15102 15076 15108 15088
rect 9732 15048 10824 15076
rect 13096 15048 15108 15076
rect 9732 15036 9738 15048
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7708 14980 8217 15008
rect 7708 14968 7714 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9263 14980 9873 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 9861 14971 9919 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11238 15008 11244 15020
rect 11011 14980 11244 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 8294 14940 8300 14952
rect 7300 14912 8300 14940
rect 7101 14903 7159 14909
rect 2648 14844 4660 14872
rect 4985 14875 5043 14881
rect 2648 14832 2654 14844
rect 4985 14841 4997 14875
rect 5031 14841 5043 14875
rect 4985 14835 5043 14841
rect 5442 14832 5448 14884
rect 5500 14872 5506 14884
rect 7116 14872 7144 14903
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14909 8447 14943
rect 9306 14940 9312 14952
rect 9267 14912 9312 14940
rect 8389 14903 8447 14909
rect 5500 14844 7144 14872
rect 7208 14844 7696 14872
rect 5500 14832 5506 14844
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 5316 14776 6377 14804
rect 5316 14764 5322 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6365 14767 6423 14773
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7208 14804 7236 14844
rect 7558 14804 7564 14816
rect 6880 14776 7236 14804
rect 7519 14776 7564 14804
rect 6880 14764 6886 14776
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7668 14804 7696 14844
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8404 14872 8432 14903
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 12986 14940 12992 14952
rect 9493 14903 9551 14909
rect 12406 14912 12992 14940
rect 7984 14844 8432 14872
rect 9508 14872 9536 14903
rect 12406 14872 12434 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 9508 14844 12434 14872
rect 7984 14832 7990 14844
rect 8849 14807 8907 14813
rect 8849 14804 8861 14807
rect 7668 14776 8861 14804
rect 8849 14773 8861 14776
rect 8895 14773 8907 14807
rect 8849 14767 8907 14773
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 13096 14804 13124 15048
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 16056 15079 16114 15085
rect 16056 15045 16068 15079
rect 16102 15076 16114 15079
rect 17972 15076 18000 15116
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19978 15144 19984 15156
rect 19536 15116 19984 15144
rect 18509 15079 18567 15085
rect 18509 15076 18521 15079
rect 16102 15048 18000 15076
rect 18064 15048 18521 15076
rect 16102 15045 16114 15048
rect 16056 15039 16114 15045
rect 13440 15011 13498 15017
rect 13440 14977 13452 15011
rect 13486 15008 13498 15011
rect 14826 15008 14832 15020
rect 13486 14980 14832 15008
rect 13486 14977 13498 14980
rect 13440 14971 13498 14977
rect 14826 14968 14832 14980
rect 14884 15008 14890 15020
rect 15194 15008 15200 15020
rect 14884 14980 15200 15008
rect 14884 14968 14890 14980
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 16298 15008 16304 15020
rect 16259 14980 16304 15008
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 17954 14968 17960 15020
rect 18012 15017 18018 15020
rect 18012 15008 18024 15017
rect 18064 15008 18092 15048
rect 18509 15045 18521 15048
rect 18555 15076 18567 15079
rect 19536 15076 19564 15116
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 18555 15048 19564 15076
rect 18555 15045 18567 15048
rect 18509 15039 18567 15045
rect 19702 15036 19708 15088
rect 19760 15076 19766 15088
rect 19760 15048 21404 15076
rect 19760 15036 19766 15048
rect 21376 15020 21404 15048
rect 18012 14980 18092 15008
rect 18012 14971 18024 14980
rect 18012 14968 18018 14971
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 18874 15008 18880 15020
rect 18288 14980 18880 15008
rect 18288 14968 18294 14980
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 21094 15011 21152 15017
rect 21094 15008 21106 15011
rect 18984 14980 21106 15008
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 9456 14776 13124 14804
rect 13188 14804 13216 14903
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 15010 14940 15016 14952
rect 14332 14912 15016 14940
rect 14332 14900 14338 14912
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 14182 14832 14188 14884
rect 14240 14872 14246 14884
rect 15286 14872 15292 14884
rect 14240 14844 15292 14872
rect 14240 14832 14246 14844
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 13814 14804 13820 14816
rect 13188 14776 13820 14804
rect 9456 14764 9462 14776
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14918 14804 14924 14816
rect 14879 14776 14924 14804
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15010 14764 15016 14816
rect 15068 14804 15074 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15068 14776 16865 14804
rect 15068 14764 15074 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 18984 14804 19012 14980
rect 21094 14977 21106 14980
rect 21140 14977 21152 15011
rect 21358 15008 21364 15020
rect 21319 14980 21364 15008
rect 21094 14971 21152 14977
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 17000 14776 19012 14804
rect 19337 14807 19395 14813
rect 17000 14764 17006 14776
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19886 14804 19892 14816
rect 19383 14776 19892 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20036 14776 20081 14804
rect 20036 14764 20042 14776
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 2501 14603 2559 14609
rect 2501 14600 2513 14603
rect 2280 14572 2513 14600
rect 2280 14560 2286 14572
rect 2501 14569 2513 14572
rect 2547 14569 2559 14603
rect 2501 14563 2559 14569
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 3510 14600 3516 14612
rect 3200 14572 3516 14600
rect 3200 14560 3206 14572
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 3970 14600 3976 14612
rect 3931 14572 3976 14600
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 5350 14600 5356 14612
rect 5311 14572 5356 14600
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14600 5871 14603
rect 5994 14600 6000 14612
rect 5859 14572 6000 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6638 14600 6644 14612
rect 6595 14572 6644 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 6822 14600 6828 14612
rect 6783 14572 6828 14600
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7466 14600 7472 14612
rect 7331 14572 7472 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7650 14600 7656 14612
rect 7611 14572 7656 14600
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14600 8355 14603
rect 8478 14600 8484 14612
rect 8343 14572 8484 14600
rect 8343 14569 8355 14572
rect 8297 14563 8355 14569
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9306 14600 9312 14612
rect 8987 14572 9312 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 16209 14603 16267 14609
rect 13648 14572 15884 14600
rect 2682 14492 2688 14544
rect 2740 14492 2746 14544
rect 3421 14535 3479 14541
rect 3421 14501 3433 14535
rect 3467 14532 3479 14535
rect 4338 14532 4344 14544
rect 3467 14504 4344 14532
rect 3467 14501 3479 14504
rect 3421 14495 3479 14501
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 5077 14535 5135 14541
rect 5077 14532 5089 14535
rect 4632 14504 5089 14532
rect 2700 14464 2728 14492
rect 4632 14476 4660 14504
rect 5077 14501 5089 14504
rect 5123 14532 5135 14535
rect 10870 14532 10876 14544
rect 5123 14504 10876 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 4430 14464 4436 14476
rect 2700 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4672 14436 4765 14464
rect 4672 14424 4678 14436
rect 5534 14424 5540 14476
rect 5592 14424 5598 14476
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6546 14464 6552 14476
rect 6227 14436 6552 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 6972 14436 8248 14464
rect 6972 14424 6978 14436
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14396 2743 14399
rect 3142 14396 3148 14408
rect 2731 14368 3148 14396
rect 2731 14365 2743 14368
rect 2685 14359 2743 14365
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 4338 14396 4344 14408
rect 4251 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14396 4402 14408
rect 4706 14396 4712 14408
rect 4396 14368 4712 14396
rect 4396 14356 4402 14368
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 5552 14328 5580 14424
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 7616 14368 8125 14396
rect 7616 14356 7622 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8220 14396 8248 14436
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 8444 14436 9413 14464
rect 8444 14424 8450 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10502 14464 10508 14476
rect 9631 14436 10508 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 12434 14464 12440 14476
rect 10735 14436 12440 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 13648 14396 13676 14572
rect 15856 14541 15884 14572
rect 16209 14569 16221 14603
rect 16255 14600 16267 14603
rect 16298 14600 16304 14612
rect 16255 14572 16304 14600
rect 16255 14569 16267 14572
rect 16209 14563 16267 14569
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 16577 14603 16635 14609
rect 16577 14569 16589 14603
rect 16623 14600 16635 14603
rect 17034 14600 17040 14612
rect 16623 14572 17040 14600
rect 16623 14569 16635 14572
rect 16577 14563 16635 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 18230 14600 18236 14612
rect 18191 14572 18236 14600
rect 18230 14560 18236 14572
rect 18288 14560 18294 14612
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19702 14600 19708 14612
rect 19383 14572 19708 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 15841 14535 15899 14541
rect 15841 14501 15853 14535
rect 15887 14532 15899 14535
rect 16942 14532 16948 14544
rect 15887 14504 16948 14532
rect 15887 14501 15899 14504
rect 15841 14495 15899 14501
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 17957 14467 18015 14473
rect 17957 14433 17969 14467
rect 18003 14464 18015 14467
rect 18248 14464 18276 14560
rect 19889 14535 19947 14541
rect 19889 14501 19901 14535
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 19904 14464 19932 14495
rect 18003 14436 18276 14464
rect 18340 14436 19932 14464
rect 21269 14467 21327 14473
rect 18003 14433 18015 14436
rect 17957 14427 18015 14433
rect 8220 14368 13676 14396
rect 13725 14399 13783 14405
rect 8113 14359 8171 14365
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 13814 14396 13820 14408
rect 13771 14368 13820 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 13814 14356 13820 14368
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14139 14368 14473 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 18340 14396 18368 14436
rect 21269 14433 21281 14467
rect 21315 14464 21327 14467
rect 21358 14464 21364 14476
rect 21315 14436 21364 14464
rect 21315 14433 21327 14436
rect 21269 14427 21327 14433
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 15160 14368 18368 14396
rect 15160 14356 15166 14368
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 21002 14399 21060 14405
rect 21002 14396 21014 14399
rect 19944 14368 21014 14396
rect 19944 14356 19950 14368
rect 21002 14365 21014 14368
rect 21048 14365 21060 14399
rect 21002 14359 21060 14365
rect 14274 14328 14280 14340
rect 2464 14300 5488 14328
rect 5552 14300 14280 14328
rect 2464 14288 2470 14300
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2038 14260 2044 14272
rect 1999 14232 2044 14260
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 2958 14260 2964 14272
rect 2919 14232 2964 14260
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 5460 14260 5488 14300
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 14706 14331 14764 14337
rect 14706 14328 14718 14331
rect 14424 14300 14718 14328
rect 14424 14288 14430 14300
rect 14706 14297 14718 14300
rect 14752 14297 14764 14331
rect 14706 14291 14764 14297
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 15344 14300 17632 14328
rect 15344 14288 15350 14300
rect 5626 14260 5632 14272
rect 5460 14232 5632 14260
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 6880 14232 9321 14260
rect 6880 14220 6886 14232
rect 9309 14229 9321 14232
rect 9355 14260 9367 14263
rect 9674 14260 9680 14272
rect 9355 14232 9680 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10778 14260 10784 14272
rect 10739 14232 10784 14260
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11517 14263 11575 14269
rect 11517 14260 11529 14263
rect 10919 14232 11529 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 11517 14229 11529 14232
rect 11563 14229 11575 14263
rect 11517 14223 11575 14229
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 14550 14260 14556 14272
rect 12032 14232 14556 14260
rect 12032 14220 12038 14232
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 17604 14260 17632 14300
rect 17678 14288 17684 14340
rect 17736 14337 17742 14340
rect 17736 14328 17748 14337
rect 19794 14328 19800 14340
rect 17736 14300 19800 14328
rect 17736 14291 17748 14300
rect 17736 14288 17742 14291
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 18506 14260 18512 14272
rect 17604 14232 18512 14260
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 18877 14263 18935 14269
rect 18877 14229 18889 14263
rect 18923 14260 18935 14263
rect 19058 14260 19064 14272
rect 18923 14232 19064 14260
rect 18923 14229 18935 14232
rect 18877 14223 18935 14229
rect 19058 14220 19064 14232
rect 19116 14220 19122 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 3053 14059 3111 14065
rect 3053 14056 3065 14059
rect 2455 14028 3065 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 3053 14025 3065 14028
rect 3099 14025 3111 14059
rect 3053 14019 3111 14025
rect 3326 14016 3332 14068
rect 3384 14056 3390 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 3384 14028 3525 14056
rect 3384 14016 3390 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 3513 14019 3571 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 5810 14056 5816 14068
rect 5675 14028 5816 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8110 14056 8116 14068
rect 8067 14028 8116 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8435 14028 9137 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 9125 14025 9137 14028
rect 9171 14056 9183 14059
rect 9214 14056 9220 14068
rect 9171 14028 9220 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9674 14056 9680 14068
rect 9539 14028 9680 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9824 14028 9873 14056
rect 9824 14016 9830 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 15010 14056 15016 14068
rect 9861 14019 9919 14025
rect 13924 14028 15016 14056
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 3344 13960 5181 13988
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1636 13892 1685 13920
rect 1636 13880 1642 13892
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13821 2191 13855
rect 2314 13852 2320 13864
rect 2275 13824 2320 13852
rect 2133 13815 2191 13821
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2148 13716 2176 13815
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 3344 13852 3372 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 10778 13988 10784 14000
rect 6052 13960 10784 13988
rect 6052 13948 6058 13960
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12802 13948 12808 14000
rect 12860 13988 12866 14000
rect 13924 13988 13952 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 16390 14056 16396 14068
rect 15243 14028 16396 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 12860 13960 13952 13988
rect 12860 13948 12866 13960
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3510 13920 3516 13932
rect 3467 13892 3516 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 4062 13920 4068 13932
rect 3568 13892 4068 13920
rect 3568 13880 3574 13892
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4212 13892 5273 13920
rect 4212 13880 4218 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 6871 13892 7481 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7469 13889 7481 13892
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8352 13892 8493 13920
rect 8352 13880 8358 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10275 13892 10885 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 13285 13923 13343 13929
rect 13285 13920 13297 13923
rect 12584 13892 13297 13920
rect 12584 13880 12590 13892
rect 13285 13889 13297 13892
rect 13331 13920 13343 13923
rect 13541 13923 13599 13929
rect 13331 13892 13501 13920
rect 13331 13889 13343 13892
rect 13285 13883 13343 13889
rect 2792 13824 3372 13852
rect 3697 13855 3755 13861
rect 2792 13793 2820 13824
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5997 13855 6055 13861
rect 5123 13824 5212 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 2777 13787 2835 13793
rect 2777 13753 2789 13787
rect 2823 13753 2835 13787
rect 3712 13784 3740 13815
rect 5184 13796 5212 13824
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6086 13852 6092 13864
rect 6043 13824 6092 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6086 13812 6092 13824
rect 6144 13852 6150 13864
rect 6546 13852 6552 13864
rect 6144 13824 6552 13852
rect 6144 13812 6150 13824
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 7834 13852 7840 13864
rect 6779 13824 7840 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 4065 13787 4123 13793
rect 4065 13784 4077 13787
rect 3712 13756 4077 13784
rect 2777 13747 2835 13753
rect 4065 13753 4077 13756
rect 4111 13784 4123 13787
rect 4614 13784 4620 13796
rect 4111 13756 4620 13784
rect 4111 13753 4123 13756
rect 4065 13747 4123 13753
rect 4614 13744 4620 13756
rect 4672 13744 4678 13796
rect 5166 13744 5172 13796
rect 5224 13744 5230 13796
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6656 13784 6684 13815
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 8665 13815 8723 13821
rect 6822 13784 6828 13796
rect 5592 13756 6828 13784
rect 5592 13744 5598 13756
rect 6822 13744 6828 13756
rect 6880 13744 6886 13796
rect 8680 13784 8708 13815
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13821 10563 13855
rect 13473 13852 13501 13892
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13814 13920 13820 13932
rect 13587 13892 13820 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 13924 13920 13952 13960
rect 14734 13948 14740 14000
rect 14792 13988 14798 14000
rect 15212 13988 15240 14019
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 16666 14056 16672 14068
rect 16627 14028 16672 14056
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17218 14056 17224 14068
rect 17083 14028 17224 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 18506 14016 18512 14068
rect 18564 14056 18570 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 18564 14028 20729 14056
rect 18564 14016 18570 14028
rect 20717 14025 20729 14028
rect 20763 14056 20775 14059
rect 20990 14056 20996 14068
rect 20763 14028 20996 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 21358 14056 21364 14068
rect 21223 14028 21364 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 21082 13988 21088 14000
rect 14792 13960 15240 13988
rect 18432 13960 21088 13988
rect 14792 13948 14798 13960
rect 14073 13923 14131 13929
rect 14073 13920 14085 13923
rect 13924 13892 14085 13920
rect 14073 13889 14085 13892
rect 14119 13889 14131 13923
rect 14073 13883 14131 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 15979 13892 16620 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 13473 13824 13584 13852
rect 10505 13815 10563 13821
rect 9214 13784 9220 13796
rect 8680 13756 9220 13784
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 10520 13784 10548 13815
rect 10520 13756 12434 13784
rect 2958 13716 2964 13728
rect 2148 13688 2964 13716
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 8478 13716 8484 13728
rect 5316 13688 8484 13716
rect 5316 13676 5322 13688
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 12158 13716 12164 13728
rect 12119 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12406 13716 12434 13756
rect 13354 13716 13360 13728
rect 12406 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13556 13716 13584 13824
rect 15286 13812 15292 13864
rect 15344 13852 15350 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 15344 13824 16313 13852
rect 15344 13812 15350 13824
rect 16301 13821 16313 13824
rect 16347 13852 16359 13855
rect 16482 13852 16488 13864
rect 16347 13824 16488 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16592 13852 16620 13892
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 18432 13920 18460 13960
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 16816 13892 18460 13920
rect 16816 13880 16822 13892
rect 18506 13880 18512 13932
rect 18564 13929 18570 13932
rect 18564 13920 18576 13929
rect 18785 13923 18843 13929
rect 18564 13892 18609 13920
rect 18564 13883 18576 13892
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 18874 13920 18880 13932
rect 18831 13892 18880 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 18564 13880 18570 13883
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 20185 13923 20243 13929
rect 20185 13889 20197 13923
rect 20231 13920 20243 13923
rect 20346 13920 20352 13932
rect 20231 13892 20352 13920
rect 20231 13889 20243 13892
rect 20185 13883 20243 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 20898 13920 20904 13932
rect 20487 13892 20904 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20898 13880 20904 13892
rect 20956 13920 20962 13932
rect 21192 13920 21220 14019
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 20956 13892 21220 13920
rect 20956 13880 20962 13892
rect 17586 13852 17592 13864
rect 16592 13824 17592 13852
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 15194 13744 15200 13796
rect 15252 13784 15258 13796
rect 15654 13784 15660 13796
rect 15252 13756 15660 13784
rect 15252 13744 15258 13756
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 18782 13744 18788 13796
rect 18840 13784 18846 13796
rect 18966 13784 18972 13796
rect 18840 13756 18972 13784
rect 18840 13744 18846 13756
rect 18966 13744 18972 13756
rect 19024 13784 19030 13796
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 19024 13756 19073 13784
rect 19024 13744 19030 13756
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 14918 13716 14924 13728
rect 13556 13688 14924 13716
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15565 13719 15623 13725
rect 15565 13685 15577 13719
rect 15611 13716 15623 13719
rect 16022 13716 16028 13728
rect 15611 13688 16028 13716
rect 15611 13685 15623 13688
rect 15565 13679 15623 13685
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2372 13484 2697 13512
rect 2372 13472 2378 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 3973 13515 4031 13521
rect 3973 13512 3985 13515
rect 3936 13484 3985 13512
rect 3936 13472 3942 13484
rect 3973 13481 3985 13484
rect 4019 13481 4031 13515
rect 3973 13475 4031 13481
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 4580 13484 6377 13512
rect 4580 13472 4586 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 6365 13475 6423 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9490 13512 9496 13524
rect 9272 13484 9496 13512
rect 9272 13472 9278 13484
rect 9490 13472 9496 13484
rect 9548 13512 9554 13524
rect 9548 13484 15056 13512
rect 9548 13472 9554 13484
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13444 2467 13447
rect 2498 13444 2504 13456
rect 2455 13416 2504 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 4614 13444 4620 13456
rect 3344 13416 4620 13444
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3344 13385 3372 13416
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 5810 13444 5816 13456
rect 5771 13416 5816 13444
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 9033 13447 9091 13453
rect 9033 13413 9045 13447
rect 9079 13444 9091 13447
rect 9306 13444 9312 13456
rect 9079 13416 9312 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 12158 13404 12164 13456
rect 12216 13404 12222 13456
rect 15028 13444 15056 13484
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 19576 13484 21189 13512
rect 19576 13472 19582 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21177 13475 21235 13481
rect 15194 13444 15200 13456
rect 15028 13416 15200 13444
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15436 13416 15485 13444
rect 15436 13404 15442 13416
rect 15473 13413 15485 13416
rect 15519 13444 15531 13447
rect 16942 13444 16948 13456
rect 15519 13416 16948 13444
rect 15519 13413 15531 13416
rect 15473 13407 15531 13413
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 18877 13447 18935 13453
rect 18877 13413 18889 13447
rect 18923 13444 18935 13447
rect 19610 13444 19616 13456
rect 18923 13416 19616 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2832 13348 3157 13376
rect 2832 13336 2838 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 4062 13376 4068 13388
rect 3936 13348 4068 13376
rect 3936 13336 3942 13348
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4430 13336 4436 13388
rect 4488 13336 4494 13388
rect 4525 13379 4583 13385
rect 4525 13345 4537 13379
rect 4571 13376 4583 13379
rect 4798 13376 4804 13388
rect 4571 13348 4804 13376
rect 4571 13345 4583 13348
rect 4525 13339 4583 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5261 13379 5319 13385
rect 5261 13345 5273 13379
rect 5307 13376 5319 13379
rect 6086 13376 6092 13388
rect 5307 13348 6092 13376
rect 5307 13345 5319 13348
rect 5261 13339 5319 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6788 13348 6929 13376
rect 6788 13336 6794 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 8202 13336 8208 13388
rect 8260 13376 8266 13388
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 8260 13348 8401 13376
rect 8260 13336 8266 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11204 13348 11345 13376
rect 11204 13336 11210 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13376 11575 13379
rect 11882 13376 11888 13388
rect 11563 13348 11888 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12176 13376 12204 13404
rect 12084 13348 12204 13376
rect 15841 13379 15899 13385
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13308 1458 13320
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1452 13280 1869 13308
rect 1452 13268 1458 13280
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 4338 13308 4344 13320
rect 3099 13280 4344 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4448 13308 4476 13336
rect 5350 13308 5356 13320
rect 4448 13280 5356 13308
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 6880 13280 11376 13308
rect 6880 13268 6886 13280
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 4433 13243 4491 13249
rect 4433 13240 4445 13243
rect 4120 13212 4445 13240
rect 4120 13200 4126 13212
rect 4433 13209 4445 13212
rect 4479 13209 4491 13243
rect 4433 13203 4491 13209
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 5445 13243 5503 13249
rect 5445 13240 5457 13243
rect 4580 13212 5457 13240
rect 4580 13200 4586 13212
rect 5445 13209 5457 13212
rect 5491 13209 5503 13243
rect 5445 13203 5503 13209
rect 6733 13243 6791 13249
rect 6733 13209 6745 13243
rect 6779 13240 6791 13243
rect 7377 13243 7435 13249
rect 7377 13240 7389 13243
rect 6779 13212 7389 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 7377 13209 7389 13212
rect 7423 13209 7435 13243
rect 7377 13203 7435 13209
rect 8297 13243 8355 13249
rect 8297 13209 8309 13243
rect 8343 13240 8355 13243
rect 9306 13240 9312 13252
rect 8343 13212 9312 13240
rect 8343 13209 8355 13212
rect 8297 13203 8355 13209
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10505 13243 10563 13249
rect 10505 13240 10517 13243
rect 10468 13212 10517 13240
rect 10468 13200 10474 13212
rect 10505 13209 10517 13212
rect 10551 13240 10563 13243
rect 10962 13240 10968 13252
rect 10551 13212 10968 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11241 13243 11299 13249
rect 11241 13240 11253 13243
rect 11020 13212 11253 13240
rect 11020 13200 11026 13212
rect 11241 13209 11253 13212
rect 11287 13209 11299 13243
rect 11241 13203 11299 13209
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2958 13172 2964 13184
rect 1627 13144 2964 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 3936 13144 4353 13172
rect 3936 13132 3942 13144
rect 4341 13141 4353 13144
rect 4387 13172 4399 13175
rect 5534 13172 5540 13184
rect 4387 13144 5540 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 6880 13144 6925 13172
rect 6880 13132 6886 13144
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7524 13144 8217 13172
rect 7524 13132 7530 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 8205 13135 8263 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11348 13172 11376 13280
rect 12084 13240 12112 13348
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16022 13376 16028 13388
rect 15887 13348 16028 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16022 13336 16028 13348
rect 16080 13376 16086 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 16080 13348 16405 13376
rect 16080 13336 16086 13348
rect 16393 13345 16405 13348
rect 16439 13376 16451 13379
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16439 13348 16865 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 16853 13345 16865 13348
rect 16899 13376 16911 13379
rect 17221 13379 17279 13385
rect 17221 13376 17233 13379
rect 16899 13348 17233 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17221 13345 17233 13348
rect 17267 13376 17279 13379
rect 17402 13376 17408 13388
rect 17267 13348 17408 13376
rect 17267 13345 17279 13348
rect 17221 13339 17279 13345
rect 17402 13336 17408 13348
rect 17460 13376 17466 13388
rect 17497 13379 17555 13385
rect 17497 13376 17509 13379
rect 17460 13348 17509 13376
rect 17460 13336 17466 13348
rect 17497 13345 17509 13348
rect 17543 13345 17555 13379
rect 20898 13376 20904 13388
rect 20859 13348 20904 13376
rect 17497 13339 17555 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 13814 13308 13820 13320
rect 12207 13280 13820 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 13814 13268 13820 13280
rect 13872 13308 13878 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13872 13280 14105 13308
rect 13872 13268 13878 13280
rect 14093 13277 14105 13280
rect 14139 13308 14151 13311
rect 14826 13308 14832 13320
rect 14139 13280 14832 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 17753 13311 17811 13317
rect 17753 13308 17765 13311
rect 16540 13280 17765 13308
rect 16540 13268 16546 13280
rect 17753 13277 17765 13280
rect 17799 13308 17811 13311
rect 17799 13280 19012 13308
rect 17799 13277 17811 13280
rect 17753 13271 17811 13277
rect 12406 13243 12464 13249
rect 12406 13240 12418 13243
rect 12084 13212 12418 13240
rect 12406 13209 12418 13212
rect 12452 13209 12464 13243
rect 13998 13240 14004 13252
rect 12406 13203 12464 13209
rect 13280 13212 14004 13240
rect 13280 13172 13308 13212
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14360 13243 14418 13249
rect 14360 13209 14372 13243
rect 14406 13209 14418 13243
rect 18984 13240 19012 13280
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 19116 13280 21373 13308
rect 19116 13268 19122 13280
rect 21361 13277 21373 13280
rect 21407 13308 21419 13311
rect 21450 13308 21456 13320
rect 21407 13280 21456 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 19334 13240 19340 13252
rect 18984 13212 19340 13240
rect 14360 13203 14418 13209
rect 11348 13144 13308 13172
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13412 13144 13553 13172
rect 13412 13132 13418 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 14384 13172 14412 13203
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 19978 13240 19984 13252
rect 19392 13212 19984 13240
rect 19392 13200 19398 13212
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20070 13200 20076 13252
rect 20128 13240 20134 13252
rect 20656 13243 20714 13249
rect 20656 13240 20668 13243
rect 20128 13212 20668 13240
rect 20128 13200 20134 13212
rect 20656 13209 20668 13212
rect 20702 13240 20714 13243
rect 20806 13240 20812 13252
rect 20702 13212 20812 13240
rect 20702 13209 20714 13212
rect 20656 13203 20714 13209
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 14550 13172 14556 13184
rect 14384 13144 14556 13172
rect 13541 13135 13599 13141
rect 14550 13132 14556 13144
rect 14608 13172 14614 13184
rect 15010 13172 15016 13184
rect 14608 13144 15016 13172
rect 14608 13132 14614 13144
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 19521 13175 19579 13181
rect 19521 13141 19533 13175
rect 19567 13172 19579 13175
rect 20346 13172 20352 13184
rect 19567 13144 20352 13172
rect 19567 13141 19579 13144
rect 19521 13135 19579 13141
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 4062 12968 4068 12980
rect 3384 12940 4068 12968
rect 3384 12928 3390 12940
rect 4062 12928 4068 12940
rect 4120 12968 4126 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4120 12940 5273 12968
rect 4120 12928 4126 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5261 12931 5319 12937
rect 5721 12971 5779 12977
rect 5721 12937 5733 12971
rect 5767 12968 5779 12971
rect 5994 12968 6000 12980
rect 5767 12940 6000 12968
rect 5767 12937 5779 12940
rect 5721 12931 5779 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 7101 12971 7159 12977
rect 7101 12937 7113 12971
rect 7147 12968 7159 12971
rect 7282 12968 7288 12980
rect 7147 12940 7288 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8159 12940 8677 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 8665 12931 8723 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 12805 12971 12863 12977
rect 12805 12937 12817 12971
rect 12851 12968 12863 12971
rect 13814 12968 13820 12980
rect 12851 12940 13820 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 14976 12940 16681 12968
rect 14976 12928 14982 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 18417 12971 18475 12977
rect 18417 12937 18429 12971
rect 18463 12968 18475 12971
rect 18874 12968 18880 12980
rect 18463 12940 18880 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 1780 12872 4200 12900
rect 1780 12841 1808 12872
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 2096 12804 2237 12832
rect 2096 12792 2102 12804
rect 2225 12801 2237 12804
rect 2271 12832 2283 12835
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 2271 12804 2697 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3108 12736 3525 12764
rect 3108 12724 3114 12736
rect 3513 12733 3525 12736
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 1394 12696 1400 12708
rect 1355 12668 1400 12696
rect 1394 12656 1400 12668
rect 1452 12656 1458 12708
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 4062 12696 4068 12708
rect 2455 12668 4068 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 4172 12696 4200 12872
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 6641 12903 6699 12909
rect 6641 12900 6653 12903
rect 4488 12872 6653 12900
rect 4488 12860 4494 12872
rect 6641 12869 6653 12872
rect 6687 12869 6699 12903
rect 8570 12900 8576 12912
rect 6641 12863 6699 12869
rect 7944 12872 8576 12900
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 4672 12804 5365 12832
rect 4672 12792 4678 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6328 12804 6745 12832
rect 6328 12792 6334 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 4338 12764 4344 12776
rect 4299 12736 4344 12764
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5258 12764 5264 12776
rect 5215 12736 5264 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 6549 12767 6607 12773
rect 6549 12733 6561 12767
rect 6595 12764 6607 12767
rect 7944 12764 7972 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9677 12903 9735 12909
rect 9677 12900 9689 12903
rect 9048 12872 9689 12900
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 8386 12832 8392 12844
rect 8067 12804 8392 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 9048 12841 9076 12872
rect 9677 12869 9689 12872
rect 9723 12869 9735 12903
rect 13538 12900 13544 12912
rect 9677 12863 9735 12869
rect 11072 12872 13544 12900
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8536 12804 9045 12832
rect 8536 12792 8542 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 11072 12832 11100 12872
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 14216 12903 14274 12909
rect 14216 12869 14228 12903
rect 14262 12900 14274 12903
rect 15930 12900 15936 12912
rect 14262 12872 14412 12900
rect 14262 12869 14274 12872
rect 14216 12863 14274 12869
rect 14384 12844 14412 12872
rect 15120 12872 15936 12900
rect 9033 12795 9091 12801
rect 9232 12804 11100 12832
rect 11149 12835 11207 12841
rect 6595 12736 7972 12764
rect 8205 12767 8263 12773
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 8205 12733 8217 12767
rect 8251 12764 8263 12767
rect 9232 12764 9260 12804
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11195 12804 11897 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 14366 12832 14372 12844
rect 14279 12804 14372 12832
rect 11885 12795 11943 12801
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14826 12832 14832 12844
rect 14507 12804 14832 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 8251 12736 9260 12764
rect 9309 12767 9367 12773
rect 8251 12733 8263 12736
rect 8205 12727 8263 12733
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9582 12764 9588 12776
rect 9355 12736 9588 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 11974 12764 11980 12776
rect 11935 12736 11980 12764
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12158 12764 12164 12776
rect 12119 12736 12164 12764
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 14384 12764 14412 12792
rect 15120 12764 15148 12872
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 17402 12900 17408 12912
rect 16816 12872 17408 12900
rect 16816 12860 16822 12872
rect 17402 12860 17408 12872
rect 17460 12900 17466 12912
rect 17460 12872 18092 12900
rect 17460 12860 17466 12872
rect 18064 12841 18092 12872
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 14384 12736 15148 12764
rect 15580 12804 17794 12832
rect 15580 12696 15608 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 17782 12795 17840 12801
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18432 12832 18460 12931
rect 18874 12928 18880 12940
rect 18932 12968 18938 12980
rect 18969 12971 19027 12977
rect 18969 12968 18981 12971
rect 18932 12940 18981 12968
rect 18932 12928 18938 12940
rect 18969 12937 18981 12940
rect 19015 12937 19027 12971
rect 19334 12968 19340 12980
rect 19295 12940 19340 12968
rect 18969 12931 19027 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 19794 12968 19800 12980
rect 19755 12940 19800 12968
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 20898 12928 20904 12980
rect 20956 12928 20962 12980
rect 20916 12900 20944 12928
rect 20916 12872 21220 12900
rect 18095 12804 18460 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 19610 12792 19616 12844
rect 19668 12832 19674 12844
rect 21192 12841 21220 12872
rect 20910 12835 20968 12841
rect 20910 12832 20922 12835
rect 19668 12804 20922 12832
rect 19668 12792 19674 12804
rect 20910 12801 20922 12804
rect 20956 12801 20968 12835
rect 20910 12795 20968 12801
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12832 21235 12835
rect 21358 12832 21364 12844
rect 21223 12804 21364 12832
rect 21223 12801 21235 12804
rect 21177 12795 21235 12801
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 4172 12668 7788 12696
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4706 12628 4712 12640
rect 4019 12600 4712 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 5684 12600 7665 12628
rect 5684 12588 5690 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 7760 12628 7788 12668
rect 14476 12668 15608 12696
rect 8202 12628 8208 12640
rect 7760 12600 8208 12628
rect 7653 12591 7711 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 9180 12600 13093 12628
rect 9180 12588 9186 12600
rect 13081 12597 13093 12600
rect 13127 12628 13139 12631
rect 14476 12628 14504 12668
rect 14826 12628 14832 12640
rect 13127 12600 14504 12628
rect 14787 12600 14832 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 19518 12628 19524 12640
rect 15068 12600 19524 12628
rect 15068 12588 15074 12600
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 4154 12424 4160 12436
rect 3467 12396 4160 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 5902 12424 5908 12436
rect 4571 12396 5908 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 8294 12424 8300 12436
rect 7208 12396 8300 12424
rect 2866 12356 2872 12368
rect 2779 12328 2872 12356
rect 2792 12297 2820 12328
rect 2866 12316 2872 12328
rect 2924 12356 2930 12368
rect 3602 12356 3608 12368
rect 2924 12328 3608 12356
rect 2924 12316 2930 12328
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 4798 12356 4804 12368
rect 3896 12328 4804 12356
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2958 12288 2964 12300
rect 2919 12260 2964 12288
rect 2777 12251 2835 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 3896 12297 3924 12328
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 5537 12359 5595 12365
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 7208 12356 7236 12396
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9950 12424 9956 12436
rect 9723 12396 9956 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 12032 12396 12081 12424
rect 12032 12384 12038 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 17310 12424 17316 12436
rect 12069 12387 12127 12393
rect 14752 12396 17316 12424
rect 5583 12328 7236 12356
rect 7285 12359 7343 12365
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 7285 12325 7297 12359
rect 7331 12325 7343 12359
rect 14553 12359 14611 12365
rect 7285 12319 7343 12325
rect 9140 12328 9352 12356
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12257 3939 12291
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 3881 12251 3939 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5350 12288 5356 12300
rect 5123 12260 5356 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4338 12220 4344 12232
rect 4203 12192 4344 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5000 12220 5028 12251
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 6914 12288 6920 12300
rect 6779 12260 6920 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7098 12220 7104 12232
rect 5000 12192 7104 12220
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7300 12220 7328 12319
rect 8386 12288 8392 12300
rect 8347 12260 8392 12288
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 9140 12297 9168 12328
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9324 12288 9352 12328
rect 14553 12325 14565 12359
rect 14599 12356 14611 12359
rect 14752 12356 14780 12396
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18874 12424 18880 12436
rect 18835 12396 18880 12424
rect 18874 12384 18880 12396
rect 18932 12424 18938 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18932 12396 19257 12424
rect 18932 12384 18938 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 14599 12328 14780 12356
rect 14599 12325 14611 12328
rect 14553 12319 14611 12325
rect 10778 12288 10784 12300
rect 9324 12260 10784 12288
rect 9125 12251 9183 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 12526 12288 12532 12300
rect 11563 12260 12532 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 14568 12288 14596 12319
rect 16298 12316 16304 12368
rect 16356 12356 16362 12368
rect 16758 12356 16764 12368
rect 16356 12328 16764 12356
rect 16356 12316 16362 12328
rect 16758 12316 16764 12328
rect 16816 12356 16822 12368
rect 16816 12328 17172 12356
rect 16816 12316 16822 12328
rect 17144 12297 17172 12328
rect 13648 12260 14596 12288
rect 17129 12291 17187 12297
rect 10318 12220 10324 12232
rect 7300 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11112 12192 11621 12220
rect 11112 12180 11118 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 13469 12223 13527 12229
rect 13469 12220 13481 12223
rect 12032 12192 13481 12220
rect 12032 12180 12038 12192
rect 13469 12189 13481 12192
rect 13515 12220 13527 12223
rect 13648 12220 13676 12260
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 21358 12288 21364 12300
rect 21319 12260 21364 12288
rect 17129 12251 17187 12257
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 13515 12192 13676 12220
rect 13725 12223 13783 12229
rect 13515 12189 13527 12192
rect 13469 12183 13527 12189
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14182 12220 14188 12232
rect 13771 12192 14188 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14182 12180 14188 12192
rect 14240 12220 14246 12232
rect 14826 12220 14832 12232
rect 14240 12192 14832 12220
rect 14240 12180 14246 12192
rect 14826 12180 14832 12192
rect 14884 12220 14890 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14884 12192 15025 12220
rect 14884 12180 14890 12192
rect 15013 12189 15025 12192
rect 15059 12220 15071 12223
rect 16298 12220 16304 12232
rect 15059 12192 16304 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 6825 12155 6883 12161
rect 6825 12152 6837 12155
rect 5132 12124 6837 12152
rect 5132 12112 5138 12124
rect 6825 12121 6837 12124
rect 6871 12121 6883 12155
rect 6825 12115 6883 12121
rect 9309 12155 9367 12161
rect 9309 12121 9321 12155
rect 9355 12152 9367 12155
rect 9953 12155 10011 12161
rect 9953 12152 9965 12155
rect 9355 12124 9965 12152
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 9953 12121 9965 12124
rect 9999 12121 10011 12155
rect 11790 12152 11796 12164
rect 9953 12115 10011 12121
rect 10060 12124 11796 12152
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 1946 12084 1952 12096
rect 1627 12056 1952 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 5166 12084 5172 12096
rect 5127 12056 5172 12084
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 5776 12056 6929 12084
rect 5776 12044 5782 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 7340 12056 9229 12084
rect 7340 12044 7346 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10060 12084 10088 12124
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 15286 12161 15292 12164
rect 15280 12152 15292 12161
rect 15247 12124 15292 12152
rect 15280 12115 15292 12124
rect 15286 12112 15292 12115
rect 15344 12112 15350 12164
rect 17374 12155 17432 12161
rect 17374 12152 17386 12155
rect 17236 12124 17386 12152
rect 9456 12056 10088 12084
rect 11057 12087 11115 12093
rect 9456 12044 9462 12056
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11146 12084 11152 12096
rect 11103 12056 11152 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11146 12044 11152 12056
rect 11204 12084 11210 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11204 12056 11713 12084
rect 11204 12044 11210 12056
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 11701 12047 11759 12053
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 12124 12056 12357 12084
rect 12124 12044 12130 12056
rect 12345 12053 12357 12056
rect 12391 12053 12403 12087
rect 12345 12047 12403 12053
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 15470 12084 15476 12096
rect 13596 12056 15476 12084
rect 13596 12044 13602 12056
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 16390 12044 16396 12056
rect 16448 12084 16454 12096
rect 17236 12084 17264 12124
rect 17374 12121 17386 12124
rect 17420 12121 17432 12155
rect 21094 12155 21152 12161
rect 21094 12152 21106 12155
rect 17374 12115 17432 12121
rect 18524 12124 21106 12152
rect 16448 12056 17264 12084
rect 16448 12044 16454 12056
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18524 12093 18552 12124
rect 21094 12121 21106 12124
rect 21140 12152 21152 12155
rect 21266 12152 21272 12164
rect 21140 12124 21272 12152
rect 21140 12121 21152 12124
rect 21094 12115 21152 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 17920 12056 18521 12084
rect 17920 12044 17926 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 18966 12084 18972 12096
rect 18840 12056 18972 12084
rect 18840 12044 18846 12056
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19610 12084 19616 12096
rect 19571 12056 19616 12084
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20530 12084 20536 12096
rect 20027 12056 20536 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 1949 11883 2007 11889
rect 1949 11880 1961 11883
rect 1912 11852 1961 11880
rect 1912 11840 1918 11852
rect 1949 11849 1961 11852
rect 1995 11849 2007 11883
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 1949 11843 2007 11849
rect 2056 11852 2789 11880
rect 1210 11772 1216 11824
rect 1268 11812 1274 11824
rect 2056 11812 2084 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4890 11880 4896 11892
rect 4295 11852 4896 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6380 11812 6408 11843
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7834 11880 7840 11892
rect 7432 11852 7840 11880
rect 7432 11840 7438 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 8260 11852 10425 11880
rect 8260 11840 8266 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10413 11843 10471 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 11020 11852 12434 11880
rect 11020 11840 11026 11852
rect 1268 11784 2084 11812
rect 2148 11784 6408 11812
rect 12406 11812 12434 11852
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13504 11852 13829 11880
rect 13504 11840 13510 11852
rect 13817 11849 13829 11852
rect 13863 11880 13875 11883
rect 14182 11880 14188 11892
rect 13863 11852 14188 11880
rect 13863 11849 13875 11852
rect 13817 11843 13875 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15930 11880 15936 11892
rect 15891 11852 15936 11880
rect 15930 11840 15936 11852
rect 15988 11880 15994 11892
rect 17034 11880 17040 11892
rect 15988 11852 17040 11880
rect 15988 11840 15994 11852
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 17678 11880 17684 11892
rect 17639 11852 17684 11880
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19576 11852 19625 11880
rect 19576 11840 19582 11852
rect 19613 11849 19625 11852
rect 19659 11849 19671 11883
rect 21266 11880 21272 11892
rect 21227 11852 21272 11880
rect 19613 11843 19671 11849
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 16390 11812 16396 11824
rect 12406 11784 16396 11812
rect 1268 11772 1274 11784
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 2148 11753 2176 11784
rect 16390 11772 16396 11784
rect 16448 11772 16454 11824
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 18932 11784 19104 11812
rect 18932 11772 18938 11784
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 4755 11716 5365 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 7374 11744 7380 11756
rect 6595 11716 7380 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 10042 11744 10048 11756
rect 10003 11716 10048 11744
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10827 11716 11529 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 12066 11744 12072 11756
rect 11848 11716 12072 11744
rect 11848 11704 11854 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 13193 11747 13251 11753
rect 13193 11744 13205 11747
rect 12676 11716 13205 11744
rect 12676 11704 12682 11716
rect 13193 11713 13205 11716
rect 13239 11744 13251 11747
rect 13354 11744 13360 11756
rect 13239 11716 13360 11744
rect 13239 11713 13251 11716
rect 13193 11707 13251 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 13504 11716 13549 11744
rect 13504 11704 13510 11716
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 14809 11747 14867 11753
rect 14809 11744 14821 11747
rect 14516 11716 14821 11744
rect 14516 11704 14522 11716
rect 14809 11713 14821 11716
rect 14855 11713 14867 11747
rect 16298 11744 16304 11756
rect 16259 11716 16304 11744
rect 14809 11707 14867 11713
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16356 11716 16681 11744
rect 16356 11704 16362 11716
rect 16669 11713 16681 11716
rect 16715 11744 16727 11747
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16715 11716 17233 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 17221 11713 17233 11716
rect 17267 11744 17279 11747
rect 17402 11744 17408 11756
rect 17267 11716 17408 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 18782 11744 18788 11756
rect 18840 11753 18846 11756
rect 19076 11753 19104 11784
rect 20530 11772 20536 11824
rect 20588 11812 20594 11824
rect 20726 11815 20784 11821
rect 20726 11812 20738 11815
rect 20588 11784 20738 11812
rect 20588 11772 20594 11784
rect 20726 11781 20738 11784
rect 20772 11781 20784 11815
rect 20726 11775 20784 11781
rect 18752 11716 18788 11744
rect 18782 11704 18788 11716
rect 18840 11707 18852 11753
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11744 21051 11747
rect 21358 11744 21364 11756
rect 21039 11716 21364 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 18840 11704 18846 11707
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 1412 11676 1440 11704
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 1412 11648 2421 11676
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 3602 11676 3608 11688
rect 3563 11648 3608 11676
rect 2409 11639 2467 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 5442 11676 5448 11688
rect 5403 11648 5448 11676
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 4430 11608 4436 11620
rect 1627 11580 4436 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 4430 11568 4436 11580
rect 4488 11568 4494 11620
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 5552 11608 5580 11639
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 10962 11676 10968 11688
rect 6788 11648 10968 11676
rect 6788 11636 6794 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 12434 11676 12440 11688
rect 11103 11648 12440 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14240 11648 14565 11676
rect 14240 11636 14246 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 5408 11580 5580 11608
rect 5408 11568 5414 11580
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 6972 11580 12434 11608
rect 6972 11568 6978 11580
rect 1302 11500 1308 11552
rect 1360 11540 1366 11552
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 1360 11512 3157 11540
rect 1360 11500 1366 11512
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 4982 11540 4988 11552
rect 4943 11512 4988 11540
rect 3145 11503 3203 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 12066 11540 12072 11552
rect 12027 11512 12072 11540
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12406 11540 12434 11580
rect 13078 11540 13084 11552
rect 12406 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 14734 11540 14740 11552
rect 13780 11512 14740 11540
rect 13780 11500 13786 11512
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 19702 11540 19708 11552
rect 17552 11512 19708 11540
rect 17552 11500 17558 11512
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 1949 11339 2007 11345
rect 1949 11336 1961 11339
rect 1728 11308 1961 11336
rect 1728 11296 1734 11308
rect 1949 11305 1961 11308
rect 1995 11305 2007 11339
rect 2590 11336 2596 11348
rect 2551 11308 2596 11336
rect 1949 11299 2007 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3292 11308 3801 11336
rect 3292 11296 3298 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5500 11308 5549 11336
rect 5500 11296 5506 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 7282 11336 7288 11348
rect 6779 11308 7288 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8720 11308 8953 11336
rect 8720 11296 8726 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 14458 11336 14464 11348
rect 11756 11308 14464 11336
rect 11756 11296 11762 11308
rect 14458 11296 14464 11308
rect 14516 11336 14522 11348
rect 15470 11336 15476 11348
rect 14516 11308 15056 11336
rect 15431 11308 15476 11336
rect 14516 11296 14522 11308
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 4522 11268 4528 11280
rect 1627 11240 4528 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 4522 11228 4528 11240
rect 4580 11228 4586 11280
rect 5994 11268 6000 11280
rect 4908 11240 6000 11268
rect 4908 11209 4936 11240
rect 5994 11228 6000 11240
rect 6052 11268 6058 11280
rect 11974 11268 11980 11280
rect 6052 11240 11980 11268
rect 6052 11228 6058 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12526 11268 12532 11280
rect 12391 11240 12532 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 15028 11268 15056 11308
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 16132 11308 17417 11336
rect 15749 11271 15807 11277
rect 15749 11268 15761 11271
rect 15028 11240 15761 11268
rect 15749 11237 15761 11240
rect 15795 11237 15807 11271
rect 15749 11231 15807 11237
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 5534 11160 5540 11212
rect 5592 11160 5598 11212
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 9490 11200 9496 11212
rect 9451 11172 9496 11200
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 10686 11200 10692 11212
rect 10647 11172 10692 11200
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 12618 11200 12624 11212
rect 10919 11172 12624 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13814 11200 13820 11212
rect 13648 11172 13820 11200
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2774 11132 2780 11144
rect 2455 11104 2780 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2148 11064 2176 11095
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2832 11104 2881 11132
rect 2832 11092 2838 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4982 11132 4988 11144
rect 4019 11104 4988 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5552 11132 5580 11160
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 5552 11104 6285 11132
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6788 11104 7021 11132
rect 6788 11092 6794 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 7156 11104 9413 11132
rect 7156 11092 7162 11104
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10100 11104 10609 11132
rect 10100 11092 10106 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 13469 11135 13527 11141
rect 13469 11132 13481 11135
rect 11940 11104 13481 11132
rect 11940 11092 11946 11104
rect 13469 11101 13481 11104
rect 13515 11132 13527 11135
rect 13648 11132 13676 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 16132 11200 16160 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 19426 11336 19432 11348
rect 17736 11308 19432 11336
rect 17736 11296 17742 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21358 11336 21364 11348
rect 21319 11308 21364 11336
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 15160 11172 16160 11200
rect 17129 11203 17187 11209
rect 15160 11160 15166 11172
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17402 11200 17408 11212
rect 17175 11172 17408 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 18874 11200 18880 11212
rect 18831 11172 18880 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 18874 11160 18880 11172
rect 18932 11200 18938 11212
rect 18932 11172 19334 11200
rect 18932 11160 18938 11172
rect 13515 11104 13676 11132
rect 13725 11135 13783 11141
rect 13515 11101 13527 11104
rect 13469 11095 13527 11101
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13771 11104 14105 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14093 11101 14105 11104
rect 14139 11132 14151 11135
rect 14182 11132 14188 11144
rect 14139 11104 14188 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 19306 11132 19334 11172
rect 19610 11132 19616 11144
rect 19306 11104 19616 11132
rect 19610 11092 19616 11104
rect 19668 11092 19674 11144
rect 19702 11092 19708 11144
rect 19760 11132 19766 11144
rect 19869 11135 19927 11141
rect 19869 11132 19881 11135
rect 19760 11104 19881 11132
rect 19760 11092 19766 11104
rect 19869 11101 19881 11104
rect 19915 11101 19927 11135
rect 19869 11095 19927 11101
rect 4062 11064 4068 11076
rect 2148 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 5077 11067 5135 11073
rect 5077 11064 5089 11067
rect 4304 11036 5089 11064
rect 4304 11024 4310 11036
rect 5077 11033 5089 11036
rect 5123 11033 5135 11067
rect 5077 11027 5135 11033
rect 5169 11067 5227 11073
rect 5169 11033 5181 11067
rect 5215 11033 5227 11067
rect 6365 11067 6423 11073
rect 6365 11064 6377 11067
rect 5169 11027 5227 11033
rect 5644 11036 6377 11064
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 5184 10996 5212 11027
rect 5644 11008 5672 11036
rect 6365 11033 6377 11036
rect 6411 11033 6423 11067
rect 6365 11027 6423 11033
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8619 11036 9321 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 13078 11064 13084 11076
rect 10560 11036 13084 11064
rect 10560 11024 10566 11036
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 14338 11067 14396 11073
rect 14338 11064 14350 11067
rect 13556 11036 14350 11064
rect 5040 10968 5212 10996
rect 5040 10956 5046 10968
rect 5626 10956 5632 11008
rect 5684 10956 5690 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8110 10996 8116 11008
rect 7708 10968 8116 10996
rect 7708 10956 7714 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 10226 10996 10232 11008
rect 10187 10968 10232 10996
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 12434 10996 12440 11008
rect 10744 10968 12440 10996
rect 10744 10956 10750 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 13556 10996 13584 11036
rect 14338 11033 14350 11036
rect 14384 11033 14396 11067
rect 16850 11064 16856 11076
rect 16908 11073 16914 11076
rect 16820 11036 16856 11064
rect 14338 11027 14396 11033
rect 16850 11024 16856 11036
rect 16908 11027 16920 11073
rect 16908 11024 16914 11027
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 18518 11067 18576 11073
rect 18518 11064 18530 11067
rect 17276 11036 18530 11064
rect 17276 11024 17282 11036
rect 18518 11033 18530 11036
rect 18564 11064 18576 11067
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18564 11036 19257 11064
rect 18564 11033 18576 11036
rect 18518 11027 18576 11033
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 12676 10968 13584 10996
rect 12676 10956 12682 10968
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 1452 10764 2513 10792
rect 1452 10752 1458 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 3142 10792 3148 10804
rect 3103 10764 3148 10792
rect 2501 10755 2559 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3476 10764 3617 10792
rect 3476 10752 3482 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 4120 10764 5365 10792
rect 4120 10752 4126 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 6730 10792 6736 10804
rect 6691 10764 6736 10792
rect 5353 10755 5411 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7147 10764 7757 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 7745 10755 7803 10761
rect 7852 10764 9873 10792
rect 7852 10724 7880 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10284 10764 10333 10792
rect 10284 10752 10290 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 12986 10792 12992 10804
rect 12947 10764 12992 10792
rect 10321 10755 10379 10761
rect 12986 10752 12992 10764
rect 13044 10792 13050 10804
rect 13262 10792 13268 10804
rect 13044 10764 13268 10792
rect 13044 10752 13050 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14645 10795 14703 10801
rect 14645 10792 14657 10795
rect 13872 10764 14657 10792
rect 13872 10752 13878 10764
rect 14645 10761 14657 10764
rect 14691 10761 14703 10795
rect 14645 10755 14703 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18414 10792 18420 10804
rect 18371 10764 18420 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 19981 10795 20039 10801
rect 19981 10761 19993 10795
rect 20027 10792 20039 10795
rect 20070 10792 20076 10804
rect 20027 10764 20076 10792
rect 20027 10761 20039 10764
rect 19981 10755 20039 10761
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 3344 10696 7880 10724
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1486 10656 1492 10668
rect 1443 10628 1492 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 3344 10665 3372 10696
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 8536 10696 8769 10724
rect 8536 10684 8542 10696
rect 8757 10693 8769 10696
rect 8803 10724 8815 10727
rect 10134 10724 10140 10736
rect 8803 10696 10140 10724
rect 8803 10693 8815 10696
rect 8757 10687 8815 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 12713 10727 12771 10733
rect 12713 10693 12725 10727
rect 12759 10724 12771 10727
rect 13446 10724 13452 10736
rect 12759 10696 13452 10724
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 16936 10727 16994 10733
rect 16936 10693 16948 10727
rect 16982 10724 16994 10727
rect 17034 10724 17040 10736
rect 16982 10696 17040 10724
rect 16982 10693 16994 10696
rect 16936 10687 16994 10693
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 19426 10684 19432 10736
rect 19484 10733 19490 10736
rect 19484 10724 19496 10733
rect 19484 10696 19529 10724
rect 19484 10687 19496 10696
rect 19484 10684 19490 10687
rect 19610 10684 19616 10736
rect 19668 10724 19674 10736
rect 19668 10696 21404 10724
rect 19668 10684 19674 10696
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 4154 10656 4160 10668
rect 3835 10628 4160 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 5902 10656 5908 10668
rect 5583 10628 5908 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 7742 10656 7748 10668
rect 6043 10628 7748 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 9490 10656 9496 10668
rect 7883 10628 9496 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10275 10628 10885 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13814 10656 13820 10668
rect 13136 10628 13820 10656
rect 13136 10616 13142 10628
rect 13814 10616 13820 10628
rect 13872 10656 13878 10668
rect 14102 10659 14160 10665
rect 14102 10656 14114 10659
rect 13872 10628 14114 10656
rect 13872 10616 13878 10628
rect 14102 10625 14114 10628
rect 14148 10625 14160 10659
rect 14102 10619 14160 10625
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 14332 10628 14381 10656
rect 14332 10616 14338 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 15758 10659 15816 10665
rect 15758 10656 15770 10659
rect 14369 10619 14427 10625
rect 14476 10628 15770 10656
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2682 10588 2688 10600
rect 2271 10560 2688 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 6546 10588 6552 10600
rect 6507 10560 6552 10588
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7466 10588 7472 10600
rect 6687 10560 7472 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 9122 10588 9128 10600
rect 8067 10560 9128 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9306 10588 9312 10600
rect 9267 10560 9312 10588
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 12066 10588 12072 10600
rect 10551 10560 12072 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 12066 10548 12072 10560
rect 12124 10588 12130 10600
rect 12124 10560 12434 10588
rect 12124 10548 12130 10560
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 1670 10520 1676 10532
rect 1627 10492 1676 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 1854 10480 1860 10532
rect 1912 10520 1918 10532
rect 7006 10520 7012 10532
rect 1912 10492 7012 10520
rect 1912 10480 1918 10492
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7374 10520 7380 10532
rect 7335 10492 7380 10520
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 12406 10520 12434 10560
rect 12406 10492 13492 10520
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9122 10452 9128 10464
rect 8352 10424 9128 10452
rect 8352 10412 8358 10424
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 12342 10452 12348 10464
rect 11112 10424 12348 10452
rect 11112 10412 11118 10424
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 13464 10452 13492 10492
rect 14476 10452 14504 10628
rect 15758 10625 15770 10628
rect 15804 10625 15816 10659
rect 15758 10619 15816 10625
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16298 10656 16304 10668
rect 16071 10628 16304 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16298 10616 16304 10628
rect 16356 10656 16362 10668
rect 19720 10665 19748 10696
rect 21376 10668 21404 10696
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16356 10628 16681 10656
rect 16356 10616 16362 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 21082 10616 21088 10668
rect 21140 10665 21146 10668
rect 21140 10656 21152 10665
rect 21358 10656 21364 10668
rect 21140 10628 21185 10656
rect 21319 10628 21364 10656
rect 21140 10619 21152 10628
rect 21140 10616 21146 10619
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 13464 10424 14504 10452
rect 14826 10412 14832 10464
rect 14884 10452 14890 10464
rect 17310 10452 17316 10464
rect 14884 10424 17316 10452
rect 14884 10412 14890 10424
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1820 10220 1961 10248
rect 1820 10208 1826 10220
rect 1949 10217 1961 10220
rect 1995 10217 2007 10251
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 1949 10211 2007 10217
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 5442 10248 5448 10260
rect 5040 10220 5448 10248
rect 5040 10208 5046 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 5994 10248 6000 10260
rect 5767 10220 6000 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10594 10248 10600 10260
rect 9723 10220 10600 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 10744 10220 10789 10248
rect 10744 10208 10750 10220
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11296 10220 13768 10248
rect 11296 10208 11302 10220
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 2409 10183 2467 10189
rect 2409 10180 2421 10183
rect 1544 10152 2421 10180
rect 1544 10140 1550 10152
rect 2409 10149 2421 10152
rect 2455 10149 2467 10183
rect 7190 10180 7196 10192
rect 2409 10143 2467 10149
rect 4632 10152 7196 10180
rect 4632 10121 4660 10152
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 7484 10152 9076 10180
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 1412 10084 2789 10112
rect 1412 10056 1440 10084
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 5258 10112 5264 10124
rect 4847 10084 5264 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 7282 10112 7288 10124
rect 5500 10084 6960 10112
rect 7243 10084 7288 10112
rect 5500 10072 5506 10084
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 5810 10044 5816 10056
rect 2179 10016 5816 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6932 10044 6960 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7484 10121 7512 10152
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10081 7527 10115
rect 8478 10112 8484 10124
rect 8439 10084 8484 10112
rect 7469 10075 7527 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 6932 10016 7205 10044
rect 7193 10013 7205 10016
rect 7239 10044 7251 10047
rect 8570 10044 8576 10056
rect 7239 10016 8576 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 4525 9979 4583 9985
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 6730 9976 6736 9988
rect 4571 9948 6736 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 9048 9976 9076 10152
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 12345 10183 12403 10189
rect 12345 10180 12357 10183
rect 9640 10152 12357 10180
rect 9640 10140 9646 10152
rect 12345 10149 12357 10152
rect 12391 10180 12403 10183
rect 12618 10180 12624 10192
rect 12391 10152 12624 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13740 10180 13768 10220
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13872 10220 14105 10248
rect 13872 10208 13878 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14568 10220 17448 10248
rect 14568 10180 14596 10220
rect 13740 10152 14596 10180
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 11054 10112 11060 10124
rect 9171 10084 11060 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14274 10112 14280 10124
rect 13771 10084 14280 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 17420 10112 17448 10220
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 18840 10220 19349 10248
rect 18840 10208 18846 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 21082 10208 21088 10260
rect 21140 10248 21146 10260
rect 21361 10251 21419 10257
rect 21361 10248 21373 10251
rect 21140 10220 21373 10248
rect 21140 10208 21146 10220
rect 21361 10217 21373 10220
rect 21407 10217 21419 10251
rect 21361 10211 21419 10217
rect 17420 10084 17540 10112
rect 9306 10044 9312 10056
rect 9267 10016 9312 10044
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 13458 10047 13516 10053
rect 13458 10044 13470 10047
rect 12584 10016 13470 10044
rect 12584 10004 12590 10016
rect 13458 10013 13470 10016
rect 13504 10013 13516 10047
rect 13458 10007 13516 10013
rect 15217 10047 15275 10053
rect 15217 10013 15229 10047
rect 15263 10044 15275 10047
rect 15378 10044 15384 10056
rect 15263 10016 15384 10044
rect 15263 10013 15275 10016
rect 15217 10007 15275 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 16022 10044 16028 10056
rect 15519 10016 16028 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16862 10047 16920 10053
rect 16862 10013 16874 10047
rect 16908 10013 16920 10047
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 16862 10007 16920 10013
rect 16868 9976 16896 10007
rect 17126 10004 17132 10016
rect 17184 10044 17190 10056
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 17184 10016 17417 10044
rect 17184 10004 17190 10016
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17512 10044 17540 10084
rect 17661 10047 17719 10053
rect 17661 10044 17673 10047
rect 17512 10016 17673 10044
rect 17405 10007 17463 10013
rect 17661 10013 17673 10016
rect 17707 10044 17719 10047
rect 18046 10044 18052 10056
rect 17707 10016 18052 10044
rect 17707 10013 17719 10016
rect 17661 10007 17719 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 21358 10044 21364 10056
rect 20027 10016 21364 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 16942 9976 16948 9988
rect 9048 9948 15792 9976
rect 16868 9948 16948 9976
rect 15304 9920 15332 9948
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1854 9908 1860 9920
rect 1627 9880 1860 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7098 9908 7104 9920
rect 6595 9880 7104 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 8202 9908 8208 9920
rect 8163 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8352 9880 8397 9908
rect 8352 9868 8358 9880
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 9180 9880 9229 9908
rect 9180 9868 9186 9880
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 9732 9880 10333 9908
rect 9732 9868 9738 9880
rect 10321 9877 10333 9880
rect 10367 9908 10379 9911
rect 10778 9908 10784 9920
rect 10367 9880 10784 9908
rect 10367 9877 10379 9880
rect 10321 9871 10379 9877
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 14826 9908 14832 9920
rect 12492 9880 14832 9908
rect 12492 9868 12498 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15286 9868 15292 9920
rect 15344 9868 15350 9920
rect 15764 9917 15792 9948
rect 16942 9936 16948 9948
rect 17000 9936 17006 9988
rect 20226 9979 20284 9985
rect 20226 9976 20238 9979
rect 18800 9948 20238 9976
rect 15749 9911 15807 9917
rect 15749 9877 15761 9911
rect 15795 9877 15807 9911
rect 15749 9871 15807 9877
rect 18690 9868 18696 9920
rect 18748 9908 18754 9920
rect 18800 9917 18828 9948
rect 20226 9945 20238 9948
rect 20272 9945 20284 9979
rect 20226 9939 20284 9945
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18748 9880 18797 9908
rect 18748 9868 18754 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9673 1639 9707
rect 6730 9704 6736 9716
rect 6691 9676 6736 9704
rect 1581 9667 1639 9673
rect 1596 9636 1624 9667
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 9401 9707 9459 9713
rect 9401 9704 9413 9707
rect 8352 9676 9413 9704
rect 8352 9664 8358 9676
rect 9401 9673 9413 9676
rect 9447 9673 9459 9707
rect 9401 9667 9459 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 9815 9676 10425 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10778 9704 10784 9716
rect 10739 9676 10784 9704
rect 10413 9667 10471 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10873 9707 10931 9713
rect 10873 9673 10885 9707
rect 10919 9704 10931 9707
rect 10962 9704 10968 9716
rect 10919 9676 10968 9704
rect 10919 9673 10931 9676
rect 10873 9667 10931 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 17034 9704 17040 9716
rect 16995 9676 17040 9704
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 20257 9707 20315 9713
rect 20257 9673 20269 9707
rect 20303 9704 20315 9707
rect 20993 9707 21051 9713
rect 20993 9704 21005 9707
rect 20303 9676 21005 9704
rect 20303 9673 20315 9676
rect 20257 9667 20315 9673
rect 20993 9673 21005 9676
rect 21039 9704 21051 9707
rect 21358 9704 21364 9716
rect 21039 9676 21364 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 4614 9636 4620 9648
rect 1596 9608 4620 9636
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 7098 9636 7104 9648
rect 7059 9608 7104 9636
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7193 9639 7251 9645
rect 7193 9605 7205 9639
rect 7239 9636 7251 9639
rect 7466 9636 7472 9648
rect 7239 9608 7472 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 9861 9639 9919 9645
rect 7984 9608 9812 9636
rect 7984 9596 7990 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2087 9540 2544 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2222 9432 2228 9444
rect 2183 9404 2228 9432
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 2516 9432 2544 9540
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2648 9540 2693 9568
rect 2648 9528 2654 9540
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2832 9540 2877 9568
rect 2832 9528 2838 9540
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4580 9540 4721 9568
rect 4580 9528 4586 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 7374 9568 7380 9580
rect 5951 9540 7380 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9582 9568 9588 9580
rect 8803 9540 9588 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9784 9568 9812 9608
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 12434 9636 12440 9648
rect 9907 9608 12440 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 14706 9639 14764 9645
rect 14706 9636 14718 9639
rect 13188 9608 14718 9636
rect 13188 9568 13216 9608
rect 14706 9605 14718 9608
rect 14752 9605 14764 9639
rect 14706 9599 14764 9605
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 16080 9608 16221 9636
rect 16080 9596 16086 9608
rect 16209 9605 16221 9608
rect 16255 9636 16267 9639
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16255 9608 16773 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 16761 9605 16773 9608
rect 16807 9636 16819 9639
rect 17126 9636 17132 9648
rect 16807 9608 17132 9636
rect 16807 9605 16819 9608
rect 16761 9599 16819 9605
rect 17126 9596 17132 9608
rect 17184 9636 17190 9648
rect 17497 9639 17555 9645
rect 17497 9636 17509 9639
rect 17184 9608 17509 9636
rect 17184 9596 17190 9608
rect 17497 9605 17509 9608
rect 17543 9636 17555 9639
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17543 9608 18245 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 18233 9605 18245 9608
rect 18279 9636 18291 9639
rect 18969 9639 19027 9645
rect 18969 9636 18981 9639
rect 18279 9608 18981 9636
rect 18279 9605 18291 9608
rect 18233 9599 18291 9605
rect 18969 9605 18981 9608
rect 19015 9636 19027 9639
rect 20272 9636 20300 9667
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 19015 9608 20300 9636
rect 19015 9605 19027 9608
rect 18969 9599 19027 9605
rect 9784 9540 13216 9568
rect 2746 9472 5764 9500
rect 2746 9432 2774 9472
rect 5736 9441 5764 9472
rect 7282 9460 7288 9512
rect 7340 9500 7346 9512
rect 8849 9503 8907 9509
rect 7340 9472 7385 9500
rect 7340 9460 7346 9472
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 9030 9500 9036 9512
rect 8991 9472 9036 9500
rect 8849 9463 8907 9469
rect 2516 9404 2774 9432
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9401 5779 9435
rect 5721 9395 5779 9401
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 8389 9435 8447 9441
rect 8389 9432 8401 9435
rect 5960 9404 8401 9432
rect 5960 9392 5966 9404
rect 8389 9401 8401 9404
rect 8435 9401 8447 9435
rect 8864 9432 8892 9463
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 10042 9500 10048 9512
rect 9955 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9500 10106 9512
rect 10100 9472 10640 9500
rect 10100 9460 10106 9472
rect 10612 9444 10640 9472
rect 9674 9432 9680 9444
rect 8864 9404 9680 9432
rect 8389 9395 8447 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10594 9392 10600 9444
rect 10652 9392 10658 9444
rect 10888 9432 10916 9540
rect 13262 9528 13268 9580
rect 13320 9577 13326 9580
rect 13320 9568 13332 9577
rect 13541 9571 13599 9577
rect 13320 9540 13365 9568
rect 13320 9531 13332 9540
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13814 9568 13820 9580
rect 13587 9540 13820 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13320 9528 13326 9531
rect 13814 9528 13820 9540
rect 13872 9568 13878 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13872 9540 13921 9568
rect 13872 9528 13878 9540
rect 13909 9537 13921 9540
rect 13955 9568 13967 9571
rect 14274 9568 14280 9580
rect 13955 9540 14280 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14274 9528 14280 9540
rect 14332 9568 14338 9580
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 14332 9540 14473 9568
rect 14332 9528 14338 9540
rect 14461 9537 14473 9540
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 18104 9540 19809 9568
rect 18104 9528 18110 9540
rect 19797 9537 19809 9540
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 19521 9503 19579 9509
rect 11011 9472 12434 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 10888 9404 12173 9432
rect 12161 9401 12173 9404
rect 12207 9401 12219 9435
rect 12161 9395 12219 9401
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 3476 9336 4537 9364
rect 3476 9324 3482 9336
rect 4525 9333 4537 9336
rect 4571 9333 4583 9367
rect 6454 9364 6460 9376
rect 6415 9336 6460 9364
rect 4525 9327 4583 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7340 9336 7849 9364
rect 7340 9324 7346 9336
rect 7837 9333 7849 9336
rect 7883 9364 7895 9367
rect 7926 9364 7932 9376
rect 7883 9336 7932 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 7926 9324 7932 9336
rect 7984 9364 7990 9376
rect 10686 9364 10692 9376
rect 7984 9336 10692 9364
rect 7984 9324 7990 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11020 9336 11529 9364
rect 11020 9324 11026 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 12406 9364 12434 9472
rect 19521 9469 19533 9503
rect 19567 9500 19579 9503
rect 19702 9500 19708 9512
rect 19567 9472 19708 9500
rect 19567 9469 19579 9472
rect 19521 9463 19579 9469
rect 19702 9460 19708 9472
rect 19760 9460 19766 9512
rect 15838 9432 15844 9444
rect 15799 9404 15844 9432
rect 15838 9392 15844 9404
rect 15896 9432 15902 9444
rect 16942 9432 16948 9444
rect 15896 9404 16948 9432
rect 15896 9392 15902 9404
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 20530 9432 20536 9444
rect 19392 9404 20536 9432
rect 19392 9392 19398 9404
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 13170 9364 13176 9376
rect 12406 9336 13176 9364
rect 11517 9327 11575 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 18601 9367 18659 9373
rect 18601 9333 18613 9367
rect 18647 9364 18659 9367
rect 19518 9364 19524 9376
rect 18647 9336 19524 9364
rect 18647 9333 18659 9336
rect 18601 9327 18659 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1578 9120 1584 9172
rect 1636 9160 1642 9172
rect 2041 9163 2099 9169
rect 2041 9160 2053 9163
rect 1636 9132 2053 9160
rect 1636 9120 1642 9132
rect 2041 9129 2053 9132
rect 2087 9129 2099 9163
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 2041 9123 2099 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 5718 9160 5724 9172
rect 4816 9132 5724 9160
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 2501 9095 2559 9101
rect 2501 9092 2513 9095
rect 1544 9064 2513 9092
rect 1544 9052 1550 9064
rect 2501 9061 2513 9064
rect 2547 9061 2559 9095
rect 2501 9055 2559 9061
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 1412 8996 2881 9024
rect 1412 8968 1440 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 3418 8956 3424 8968
rect 2271 8928 3424 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 4816 8820 4844 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7064 9132 7297 9160
rect 7064 9120 7070 9132
rect 7285 9129 7297 9132
rect 7331 9160 7343 9163
rect 8018 9160 8024 9172
rect 7331 9132 8024 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9582 9160 9588 9172
rect 9543 9132 9588 9160
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9732 9132 10609 9160
rect 9732 9120 9738 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 13725 9163 13783 9169
rect 10744 9132 12434 9160
rect 10744 9120 10750 9132
rect 5442 9092 5448 9104
rect 5184 9064 5448 9092
rect 5184 9033 5212 9064
rect 5442 9052 5448 9064
rect 5500 9092 5506 9104
rect 7650 9092 7656 9104
rect 5500 9064 7656 9092
rect 5500 9052 5506 9064
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 12406 9092 12434 9132
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 13814 9160 13820 9172
rect 13771 9132 13820 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 16022 9160 16028 9172
rect 15983 9132 16028 9160
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 19337 9163 19395 9169
rect 19337 9129 19349 9163
rect 19383 9160 19395 9163
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 19383 9132 20453 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 20441 9129 20453 9132
rect 20487 9160 20499 9163
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 20487 9132 20821 9160
rect 20487 9129 20499 9132
rect 20441 9123 20499 9129
rect 20809 9129 20821 9132
rect 20855 9160 20867 9163
rect 21177 9163 21235 9169
rect 21177 9160 21189 9163
rect 20855 9132 21189 9160
rect 20855 9129 20867 9132
rect 20809 9123 20867 9129
rect 21177 9129 21189 9132
rect 21223 9160 21235 9163
rect 21358 9160 21364 9172
rect 21223 9132 21364 9160
rect 21223 9129 21235 9132
rect 21177 9123 21235 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 17862 9092 17868 9104
rect 11020 9064 12112 9092
rect 12406 9064 17868 9092
rect 11020 9052 11026 9064
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6454 9024 6460 9036
rect 6227 8996 6460 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6454 8984 6460 8996
rect 6512 9024 6518 9036
rect 6638 9024 6644 9036
rect 6512 8996 6644 9024
rect 6512 8984 6518 8996
rect 6638 8984 6644 8996
rect 6696 9024 6702 9036
rect 9858 9024 9864 9036
rect 6696 8996 9864 9024
rect 6696 8984 6702 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 12084 9033 12112 9064
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 19797 9095 19855 9101
rect 19797 9092 19809 9095
rect 18748 9064 19809 9092
rect 18748 9052 18754 9064
rect 19797 9061 19809 9064
rect 19843 9061 19855 9095
rect 19797 9055 19855 9061
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 10275 8996 11253 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 11241 8993 11253 8996
rect 11287 8993 11299 9027
rect 11241 8987 11299 8993
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12802 9024 12808 9036
rect 12299 8996 12808 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5994 8956 6000 8968
rect 5031 8928 6000 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 11256 8956 11284 8987
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 13722 8956 13728 8968
rect 11256 8928 13728 8956
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 5905 8891 5963 8897
rect 4939 8860 5580 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 5552 8829 5580 8860
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 5951 8860 6561 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 9309 8891 9367 8897
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 9953 8891 10011 8897
rect 9953 8888 9965 8891
rect 9355 8860 9965 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9953 8857 9965 8860
rect 9999 8857 10011 8891
rect 9953 8851 10011 8857
rect 10965 8891 11023 8897
rect 10965 8857 10977 8891
rect 11011 8888 11023 8891
rect 11011 8860 11652 8888
rect 11011 8857 11023 8860
rect 10965 8851 11023 8857
rect 1627 8792 4844 8820
rect 5537 8823 5595 8829
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 5537 8789 5549 8823
rect 5583 8789 5595 8823
rect 5537 8783 5595 8789
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8820 6055 8823
rect 6914 8820 6920 8832
rect 6043 8792 6920 8820
rect 6043 8789 6055 8792
rect 5997 8783 6055 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9398 8820 9404 8832
rect 8619 8792 9404 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 9640 8792 10057 8820
rect 9640 8780 9646 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 10045 8783 10103 8789
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11624 8829 11652 8860
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8789 11667 8823
rect 11974 8820 11980 8832
rect 11935 8792 11980 8820
rect 11609 8783 11667 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 2041 8619 2099 8625
rect 2041 8585 2053 8619
rect 2087 8616 2099 8619
rect 2130 8616 2136 8628
rect 2087 8588 2136 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 5442 8616 5448 8628
rect 5403 8588 5448 8616
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8260 8588 9045 8616
rect 8260 8576 8266 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9398 8616 9404 8628
rect 9359 8588 9404 8616
rect 9033 8579 9091 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 9548 8588 10425 8616
rect 9548 8576 9554 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10413 8579 10471 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 10962 8576 10968 8628
rect 11020 8576 11026 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 20993 8619 21051 8625
rect 12492 8588 12537 8616
rect 12492 8576 12498 8588
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21082 8616 21088 8628
rect 21039 8588 21088 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21358 8616 21364 8628
rect 21319 8588 21364 8616
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 2685 8551 2743 8557
rect 2685 8548 2697 8551
rect 1412 8520 2697 8548
rect 1412 8492 1440 8520
rect 2685 8517 2697 8520
rect 2731 8517 2743 8551
rect 2685 8511 2743 8517
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 8662 8548 8668 8560
rect 7791 8520 8668 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 10980 8548 11008 8576
rect 10183 8520 11008 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12897 8551 12955 8557
rect 12897 8548 12909 8551
rect 12216 8520 12909 8548
rect 12216 8508 12222 8520
rect 12897 8517 12909 8520
rect 12943 8517 12955 8551
rect 12897 8511 12955 8517
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8480 1918 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1912 8452 2329 8480
rect 1912 8440 1918 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7098 8480 7104 8492
rect 6779 8452 7104 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 8386 8480 8392 8492
rect 7883 8452 8392 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 8628 8452 9505 8480
rect 8628 8440 8634 8452
rect 9493 8449 9505 8452
rect 9539 8480 9551 8483
rect 9582 8480 9588 8492
rect 9539 8452 9588 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10744 8452 10793 8480
rect 10744 8440 10750 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 10781 8443 10839 8449
rect 12084 8452 12817 8480
rect 7006 8412 7012 8424
rect 6967 8384 7012 8412
rect 7006 8372 7012 8384
rect 7064 8412 7070 8424
rect 7558 8412 7564 8424
rect 7064 8384 7564 8412
rect 7064 8372 7070 8384
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8294 8412 8300 8424
rect 8067 8384 8300 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 9306 8412 9312 8424
rect 8803 8384 9312 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10042 8412 10048 8424
rect 9723 8384 10048 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10962 8412 10968 8424
rect 10923 8384 10968 8412
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 5626 8344 5632 8356
rect 1627 8316 5632 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 10928 8316 11529 8344
rect 10928 8304 10934 8316
rect 11517 8313 11529 8316
rect 11563 8344 11575 8347
rect 11974 8344 11980 8356
rect 11563 8316 11980 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 6362 8276 6368 8288
rect 6323 8248 6368 8276
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12084 8285 12112 8452
rect 12805 8449 12817 8452
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 13170 8412 13176 8424
rect 13127 8384 13176 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11940 8248 12081 8276
rect 11940 8236 11946 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 5994 8072 6000 8084
rect 5955 8044 6000 8072
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7248 8044 7297 8072
rect 7248 8032 7254 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8720 8044 8953 8072
rect 8720 8032 8726 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 8941 8035 8999 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11112 8044 12265 8072
rect 11112 8032 11118 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 5166 8004 5172 8016
rect 1627 7976 5172 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8389 8007 8447 8013
rect 8389 8004 8401 8007
rect 8352 7976 8401 8004
rect 8352 7964 8358 7976
rect 8389 7973 8401 7976
rect 8435 8004 8447 8007
rect 9214 8004 9220 8016
rect 8435 7976 9220 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 2685 7939 2743 7945
rect 2685 7936 2697 7939
rect 1412 7908 2697 7936
rect 1412 7880 1440 7908
rect 2685 7905 2697 7908
rect 2731 7905 2743 7939
rect 2685 7899 2743 7905
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6457 7939 6515 7945
rect 6457 7936 6469 7939
rect 6420 7908 6469 7936
rect 6420 7896 6426 7908
rect 6457 7905 6469 7908
rect 6503 7905 6515 7939
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 6457 7899 6515 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7926 7936 7932 7948
rect 7887 7908 7932 7936
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9548 7908 9597 7936
rect 9548 7896 9554 7908
rect 9585 7905 9597 7908
rect 9631 7936 9643 7939
rect 12710 7936 12716 7948
rect 9631 7908 10456 7936
rect 12671 7908 12716 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7868 1918 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1912 7840 2329 7868
rect 1912 7828 1918 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 2317 7831 2375 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 7834 7760 7840 7812
rect 7892 7800 7898 7812
rect 8018 7800 8024 7812
rect 7892 7772 8024 7800
rect 7892 7760 7898 7772
rect 8018 7760 8024 7772
rect 8076 7800 8082 7812
rect 10428 7809 10456 7908
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 12860 7908 12905 7936
rect 12860 7896 12866 7908
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 11940 7840 12633 7868
rect 11940 7828 11946 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 10413 7803 10471 7809
rect 8076 7772 10364 7800
rect 8076 7760 8082 7772
rect 6365 7735 6423 7741
rect 6365 7701 6377 7735
rect 6411 7732 6423 7735
rect 7006 7732 7012 7744
rect 6411 7704 7012 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7653 7735 7711 7741
rect 7653 7732 7665 7735
rect 7248 7704 7665 7732
rect 7248 7692 7254 7704
rect 7653 7701 7665 7704
rect 7699 7701 7711 7735
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 7653 7695 7711 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 10336 7732 10364 7772
rect 10413 7769 10425 7803
rect 10459 7800 10471 7803
rect 19886 7800 19892 7812
rect 10459 7772 19892 7800
rect 10459 7769 10471 7772
rect 10413 7763 10471 7769
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 11146 7732 11152 7744
rect 10336 7704 11152 7732
rect 11146 7692 11152 7704
rect 11204 7732 11210 7744
rect 11882 7732 11888 7744
rect 11204 7704 11888 7732
rect 11204 7692 11210 7704
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 2590 7528 2596 7540
rect 1627 7500 2596 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7984 7500 8033 7528
rect 7984 7488 7990 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8386 7528 8392 7540
rect 8347 7500 8392 7528
rect 8021 7491 8079 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9490 7528 9496 7540
rect 9451 7500 9496 7528
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 8849 7463 8907 7469
rect 8849 7429 8861 7463
rect 8895 7460 8907 7463
rect 10318 7460 10324 7472
rect 8895 7432 10324 7460
rect 8895 7429 8907 7432
rect 8849 7423 8907 7429
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7392 1918 7404
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 1912 7364 2329 7392
rect 1912 7352 1918 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8294 7392 8300 7404
rect 7423 7364 8300 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8294 7352 8300 7364
rect 8352 7392 8358 7404
rect 8478 7392 8484 7404
rect 8352 7364 8484 7392
rect 8352 7352 8358 7364
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 9122 7392 9128 7404
rect 8803 7364 9128 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 5166 7256 5172 7268
rect 2087 7228 5172 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5868 7160 5917 7188
rect 5868 7148 5874 7160
rect 5905 7157 5917 7160
rect 5951 7188 5963 7191
rect 6730 7188 6736 7200
rect 5951 7160 6736 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6730 7148 6736 7160
rect 6788 7188 6794 7200
rect 7484 7188 7512 7287
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 9033 7327 9091 7333
rect 7616 7296 7661 7324
rect 7616 7284 7622 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9490 7324 9496 7336
rect 9079 7296 9496 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 6788 7160 7512 7188
rect 9953 7191 10011 7197
rect 6788 7148 6794 7160
rect 9953 7157 9965 7191
rect 9999 7188 10011 7191
rect 10226 7188 10232 7200
rect 9999 7160 10232 7188
rect 9999 7157 10011 7160
rect 9953 7151 10011 7157
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1857 6987 1915 6993
rect 1857 6984 1869 6987
rect 1452 6956 1869 6984
rect 1452 6944 1458 6956
rect 1857 6953 1869 6956
rect 1903 6953 1915 6987
rect 1857 6947 1915 6953
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 8021 6987 8079 6993
rect 8021 6984 8033 6987
rect 7616 6956 8033 6984
rect 7616 6944 7622 6956
rect 7300 6888 7604 6916
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 7300 6848 7328 6888
rect 5399 6820 7328 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6780 1458 6792
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1452 6752 2237 6780
rect 1452 6740 1458 6752
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 2225 6743 2283 6749
rect 2746 6752 5733 6780
rect 2746 6712 2774 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5902 6780 5908 6792
rect 5863 6752 5908 6780
rect 5721 6743 5779 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 7064 6752 7481 6780
rect 7064 6740 7070 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7576 6780 7604 6888
rect 7668 6857 7696 6956
rect 8021 6953 8033 6956
rect 8067 6953 8079 6987
rect 8021 6947 8079 6953
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9398 6984 9404 6996
rect 9079 6956 9404 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10318 6984 10324 6996
rect 10279 6956 10324 6984
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8260 6820 8493 6848
rect 8260 6808 8266 6820
rect 8481 6817 8493 6820
rect 8527 6848 8539 6851
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 8527 6820 9505 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10226 6848 10232 6860
rect 9723 6820 10232 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10226 6808 10232 6820
rect 10284 6848 10290 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10284 6820 10977 6848
rect 10284 6808 10290 6820
rect 10965 6817 10977 6820
rect 11011 6848 11023 6851
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 11011 6820 11437 6848
rect 11011 6817 11023 6820
rect 10965 6811 11023 6817
rect 11425 6817 11437 6820
rect 11471 6848 11483 6851
rect 18598 6848 18604 6860
rect 11471 6820 18604 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 7576 6752 12434 6780
rect 7469 6743 7527 6749
rect 5166 6712 5172 6724
rect 1596 6684 2774 6712
rect 5127 6684 5172 6712
rect 1596 6653 1624 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5350 6672 5356 6724
rect 5408 6712 5414 6724
rect 6273 6715 6331 6721
rect 6273 6712 6285 6715
rect 5408 6684 6285 6712
rect 5408 6672 5414 6684
rect 6273 6681 6285 6684
rect 6319 6681 6331 6715
rect 6273 6675 6331 6681
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6712 6515 6715
rect 12406 6712 12434 6752
rect 15562 6712 15568 6724
rect 6503 6684 11468 6712
rect 12406 6684 15568 6712
rect 6503 6681 6515 6684
rect 6457 6675 6515 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7009 6647 7067 6653
rect 7009 6644 7021 6647
rect 6972 6616 7021 6644
rect 6972 6604 6978 6616
rect 7009 6613 7021 6616
rect 7055 6613 7067 6647
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7009 6607 7067 6613
rect 7374 6604 7380 6616
rect 7432 6644 7438 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 7432 6616 9413 6644
rect 7432 6604 7438 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 10686 6644 10692 6656
rect 10647 6616 10692 6644
rect 9401 6607 9459 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6644 10839 6647
rect 11054 6644 11060 6656
rect 10827 6616 11060 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11440 6644 11468 6684
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 15930 6644 15936 6656
rect 11440 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 5350 6440 5356 6452
rect 1627 6412 5356 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7616 6412 7849 6440
rect 7616 6400 7622 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 7837 6403 7895 6409
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9232 6412 9597 6440
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 1854 6304 1860 6316
rect 1815 6276 1860 6304
rect 1854 6264 1860 6276
rect 1912 6304 1918 6316
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1912 6276 2329 6304
rect 1912 6264 1918 6276
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 5868 6276 8769 6304
rect 5868 6264 5874 6276
rect 8757 6273 8769 6276
rect 8803 6304 8815 6307
rect 9232 6304 9260 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 10226 6440 10232 6452
rect 10187 6412 10232 6440
rect 9585 6403 9643 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 12250 6440 12256 6452
rect 11112 6412 12256 6440
rect 11112 6400 11118 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 10686 6372 10692 6384
rect 8803 6276 9260 6304
rect 9416 6344 10692 6372
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 9416 6236 9444 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 7248 6208 9444 6236
rect 7248 6196 7254 6208
rect 8294 6168 8300 6180
rect 6656 6140 8300 6168
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 6656 6109 6684 6140
rect 8294 6128 8300 6140
rect 8352 6168 8358 6180
rect 8389 6171 8447 6177
rect 8389 6168 8401 6171
rect 8352 6140 8401 6168
rect 8352 6128 8358 6140
rect 8389 6137 8401 6140
rect 8435 6168 8447 6171
rect 9508 6168 9536 6267
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 10226 6236 10232 6248
rect 9815 6208 10232 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 8435 6140 9536 6168
rect 8435 6137 8447 6140
rect 8389 6131 8447 6137
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 4120 6072 6653 6100
rect 4120 6060 4126 6072
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 7006 6100 7012 6112
rect 6967 6072 7012 6100
rect 6641 6063 6699 6069
rect 7006 6060 7012 6072
rect 7064 6100 7070 6112
rect 8202 6100 8208 6112
rect 7064 6072 8208 6100
rect 7064 6060 7070 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1857 5899 1915 5905
rect 1857 5896 1869 5899
rect 1452 5868 1869 5896
rect 1452 5856 1458 5868
rect 1857 5865 1869 5868
rect 1903 5865 1915 5899
rect 1857 5859 1915 5865
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 10962 5896 10968 5908
rect 2096 5868 10968 5896
rect 2096 5856 2102 5868
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 7650 5828 7656 5840
rect 1627 5800 7656 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 7650 5788 7656 5800
rect 7708 5788 7714 5840
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5692 1458 5704
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 1452 5664 2237 5692
rect 1452 5652 1458 5664
rect 2225 5661 2237 5664
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 10962 5284 10968 5296
rect 10923 5256 10968 5284
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11149 5287 11207 5293
rect 11149 5253 11161 5287
rect 11195 5284 11207 5287
rect 16206 5284 16212 5296
rect 11195 5256 16212 5284
rect 11195 5253 11207 5256
rect 11149 5247 11207 5253
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 7374 5216 7380 5228
rect 1995 5188 7380 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 2222 5148 2228 5160
rect 2183 5120 2228 5148
rect 2222 5108 2228 5120
rect 2280 5148 2286 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2280 5120 2513 5148
rect 2280 5108 2286 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 4982 4672 4988 4684
rect 1995 4644 4988 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4604 2286 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2280 4576 2513 4604
rect 2280 4564 2286 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 1486 4128 1492 4140
rect 1447 4100 1492 4128
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4128 2102 4140
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 2096 4100 2513 4128
rect 2096 4088 2102 4100
rect 2501 4097 2513 4100
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 7006 4060 7012 4072
rect 1719 4032 7012 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 10870 3992 10876 4004
rect 2271 3964 10876 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1544 3692 1961 3720
rect 1544 3680 1550 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 1673 3655 1731 3661
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 4062 3652 4068 3664
rect 1719 3624 4068 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 1486 3448 1492 3460
rect 1447 3420 1492 3448
rect 1486 3408 1492 3420
rect 1544 3448 1550 3460
rect 2317 3451 2375 3457
rect 2317 3448 2329 3451
rect 1544 3420 2329 3448
rect 1544 3408 1550 3420
rect 2317 3417 2329 3420
rect 2363 3417 2375 3451
rect 2317 3411 2375 3417
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 5810 3176 5816 3188
rect 2179 3148 5816 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 5534 3108 5540 3120
rect 1719 3080 5540 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 1486 3040 1492 3052
rect 1447 3012 1492 3040
rect 1486 3000 1492 3012
rect 1544 3000 1550 3052
rect 2038 3040 2044 3052
rect 1999 3012 2044 3040
rect 2038 3000 2044 3012
rect 2096 3040 2102 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2096 3012 2513 3040
rect 2096 3000 2102 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 1504 2972 1532 3000
rect 2869 2975 2927 2981
rect 2869 2972 2881 2975
rect 1504 2944 2881 2972
rect 2869 2941 2881 2944
rect 2915 2941 2927 2975
rect 2869 2935 2927 2941
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 7926 2564 7932 2576
rect 2823 2536 7932 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 7190 2496 7196 2508
rect 1995 2468 7196 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2428 2286 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2280 2400 3801 2428
rect 2280 2388 2286 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 11790 2428 11796 2440
rect 11751 2400 11796 2428
rect 3789 2391 3847 2397
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 2774 2360 2780 2372
rect 2639 2332 2780 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 2774 2320 2780 2332
rect 2832 2360 2838 2372
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 2832 2332 3065 2360
rect 2832 2320 2838 2332
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 11609 2295 11667 2301
rect 11609 2261 11621 2295
rect 11655 2292 11667 2295
rect 11698 2292 11704 2304
rect 11655 2264 11704 2292
rect 11655 2261 11667 2264
rect 11609 2255 11667 2261
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
<< via1 >>
rect 8484 20748 8536 20800
rect 8668 20748 8720 20800
rect 9680 20748 9732 20800
rect 18972 20748 19024 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 3148 20587 3200 20596
rect 3148 20553 3157 20587
rect 3157 20553 3191 20587
rect 3191 20553 3200 20587
rect 3148 20544 3200 20553
rect 3976 20587 4028 20596
rect 3976 20553 3985 20587
rect 3985 20553 4019 20587
rect 4019 20553 4028 20587
rect 3976 20544 4028 20553
rect 5632 20544 5684 20596
rect 7104 20544 7156 20596
rect 7380 20544 7432 20596
rect 204 20408 256 20460
rect 1308 20408 1360 20460
rect 3332 20451 3384 20460
rect 2688 20340 2740 20392
rect 3332 20417 3341 20451
rect 3341 20417 3375 20451
rect 3375 20417 3384 20451
rect 3332 20408 3384 20417
rect 3884 20408 3936 20460
rect 4528 20408 4580 20460
rect 4712 20340 4764 20392
rect 5448 20408 5500 20460
rect 7288 20476 7340 20528
rect 8024 20476 8076 20528
rect 9404 20544 9456 20596
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 11060 20544 11112 20596
rect 13084 20544 13136 20596
rect 13820 20544 13872 20596
rect 14464 20544 14516 20596
rect 15844 20544 15896 20596
rect 17040 20544 17092 20596
rect 6552 20408 6604 20460
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 6092 20340 6144 20392
rect 7748 20340 7800 20392
rect 4804 20272 4856 20324
rect 8208 20408 8260 20460
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 8576 20408 8628 20460
rect 9864 20476 9916 20528
rect 9956 20476 10008 20528
rect 9588 20408 9640 20460
rect 10324 20408 10376 20460
rect 10784 20408 10836 20460
rect 11244 20408 11296 20460
rect 11704 20408 11756 20460
rect 12164 20408 12216 20460
rect 12624 20408 12676 20460
rect 14372 20476 14424 20528
rect 13268 20408 13320 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 8024 20340 8076 20392
rect 16764 20408 16816 20460
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 17868 20408 17920 20460
rect 20720 20408 20772 20460
rect 22284 20408 22336 20460
rect 8668 20272 8720 20324
rect 2780 20204 2832 20256
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 5540 20247 5592 20256
rect 5540 20213 5549 20247
rect 5549 20213 5583 20247
rect 5583 20213 5592 20247
rect 5540 20204 5592 20213
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 6184 20204 6236 20256
rect 6828 20204 6880 20256
rect 7748 20204 7800 20256
rect 8300 20204 8352 20256
rect 8484 20204 8536 20256
rect 9128 20204 9180 20256
rect 9312 20204 9364 20256
rect 10600 20272 10652 20324
rect 17592 20340 17644 20392
rect 19800 20340 19852 20392
rect 21364 20340 21416 20392
rect 14004 20272 14056 20324
rect 14924 20272 14976 20324
rect 16304 20272 16356 20324
rect 17500 20272 17552 20324
rect 21272 20272 21324 20324
rect 9772 20204 9824 20256
rect 10692 20204 10744 20256
rect 10968 20247 11020 20256
rect 10968 20213 10977 20247
rect 10977 20213 11011 20247
rect 11011 20213 11020 20247
rect 10968 20204 11020 20213
rect 12072 20204 12124 20256
rect 12256 20247 12308 20256
rect 12256 20213 12265 20247
rect 12265 20213 12299 20247
rect 12299 20213 12308 20247
rect 12256 20204 12308 20213
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 17224 20204 17276 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 8024 20000 8076 20052
rect 8668 20000 8720 20052
rect 9956 20000 10008 20052
rect 10600 20043 10652 20052
rect 10600 20009 10609 20043
rect 10609 20009 10643 20043
rect 10643 20009 10652 20043
rect 10600 20000 10652 20009
rect 11244 20000 11296 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 12624 20043 12676 20052
rect 12624 20009 12633 20043
rect 12633 20009 12667 20043
rect 12667 20009 12676 20043
rect 12624 20000 12676 20009
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 15384 20000 15436 20052
rect 17500 20000 17552 20052
rect 18236 20000 18288 20052
rect 6092 19975 6144 19984
rect 6092 19941 6101 19975
rect 6101 19941 6135 19975
rect 6135 19941 6144 19975
rect 6092 19932 6144 19941
rect 6368 19932 6420 19984
rect 6920 19932 6972 19984
rect 9404 19932 9456 19984
rect 9680 19975 9732 19984
rect 9680 19941 9689 19975
rect 9689 19941 9723 19975
rect 9723 19941 9732 19975
rect 9680 19932 9732 19941
rect 664 19864 716 19916
rect 1216 19864 1268 19916
rect 2688 19864 2740 19916
rect 5264 19864 5316 19916
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 3516 19796 3568 19848
rect 4436 19839 4488 19848
rect 2412 19728 2464 19780
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 4620 19796 4672 19848
rect 6184 19796 6236 19848
rect 10048 19864 10100 19916
rect 10416 19932 10468 19984
rect 16764 19932 16816 19984
rect 8024 19839 8076 19848
rect 2780 19660 2832 19712
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 3976 19703 4028 19712
rect 3976 19669 3985 19703
rect 3985 19669 4019 19703
rect 4019 19669 4028 19703
rect 3976 19660 4028 19669
rect 6368 19728 6420 19780
rect 6552 19728 6604 19780
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 9128 19796 9180 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 10140 19796 10192 19848
rect 10232 19796 10284 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 19984 19864 20036 19916
rect 21364 19907 21416 19916
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 15844 19796 15896 19848
rect 5356 19660 5408 19712
rect 5816 19660 5868 19712
rect 7472 19660 7524 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7932 19703 7984 19712
rect 7564 19660 7616 19669
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 9404 19728 9456 19780
rect 10508 19660 10560 19712
rect 11888 19660 11940 19712
rect 13728 19771 13780 19780
rect 13728 19737 13737 19771
rect 13737 19737 13771 19771
rect 13771 19737 13780 19771
rect 13728 19728 13780 19737
rect 15752 19728 15804 19780
rect 18972 19796 19024 19848
rect 14372 19660 14424 19712
rect 15200 19703 15252 19712
rect 15200 19669 15209 19703
rect 15209 19669 15243 19703
rect 15243 19669 15252 19703
rect 15200 19660 15252 19669
rect 15476 19660 15528 19712
rect 17316 19660 17368 19712
rect 18328 19771 18380 19780
rect 18328 19737 18346 19771
rect 18346 19737 18380 19771
rect 18328 19728 18380 19737
rect 21272 19728 21324 19780
rect 19892 19660 19944 19712
rect 20076 19660 20128 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 4988 19456 5040 19508
rect 5356 19456 5408 19508
rect 4528 19388 4580 19440
rect 5908 19388 5960 19440
rect 6092 19456 6144 19508
rect 6644 19456 6696 19508
rect 7472 19499 7524 19508
rect 6368 19388 6420 19440
rect 6460 19388 6512 19440
rect 6920 19388 6972 19440
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 2872 19320 2924 19372
rect 3240 19320 3292 19372
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 4344 19320 4396 19372
rect 4804 19363 4856 19372
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 5724 19320 5776 19372
rect 6644 19363 6696 19372
rect 1124 19252 1176 19304
rect 4528 19252 4580 19304
rect 2136 19227 2188 19236
rect 2136 19193 2145 19227
rect 2145 19193 2179 19227
rect 2179 19193 2188 19227
rect 2136 19184 2188 19193
rect 4160 19184 4212 19236
rect 6092 19252 6144 19304
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 7472 19465 7481 19499
rect 7481 19465 7515 19499
rect 7515 19465 7524 19499
rect 7472 19456 7524 19465
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 9404 19456 9456 19508
rect 9864 19456 9916 19508
rect 10416 19456 10468 19508
rect 10784 19499 10836 19508
rect 7564 19388 7616 19440
rect 9680 19388 9732 19440
rect 10784 19465 10793 19499
rect 10793 19465 10827 19499
rect 10827 19465 10836 19499
rect 10784 19456 10836 19465
rect 13820 19456 13872 19508
rect 15200 19456 15252 19508
rect 15752 19456 15804 19508
rect 17408 19456 17460 19508
rect 18604 19456 18656 19508
rect 14648 19388 14700 19440
rect 19984 19388 20036 19440
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 9864 19363 9916 19372
rect 7104 19252 7156 19304
rect 7564 19252 7616 19304
rect 8116 19252 8168 19304
rect 8576 19252 8628 19304
rect 9312 19252 9364 19304
rect 7380 19184 7432 19236
rect 8668 19184 8720 19236
rect 9864 19329 9873 19363
rect 9873 19329 9907 19363
rect 9907 19329 9916 19363
rect 9864 19320 9916 19329
rect 9680 19252 9732 19304
rect 13544 19363 13596 19372
rect 13544 19329 13562 19363
rect 13562 19329 13596 19363
rect 13544 19320 13596 19329
rect 13728 19320 13780 19372
rect 14464 19320 14516 19372
rect 10784 19252 10836 19304
rect 12808 19252 12860 19304
rect 9772 19184 9824 19236
rect 16120 19252 16172 19304
rect 17960 19320 18012 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 20812 19363 20864 19372
rect 20812 19329 20830 19363
rect 20830 19329 20864 19363
rect 20812 19320 20864 19329
rect 21364 19320 21416 19372
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 3148 19159 3200 19168
rect 3148 19125 3157 19159
rect 3157 19125 3191 19159
rect 3191 19125 3200 19159
rect 3148 19116 3200 19125
rect 4252 19116 4304 19168
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 5448 19116 5500 19168
rect 7656 19116 7708 19168
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 9220 19116 9272 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 13636 19116 13688 19168
rect 15476 19116 15528 19168
rect 17684 19184 17736 19236
rect 15844 19116 15896 19168
rect 17592 19116 17644 19168
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 22744 19116 22796 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1676 18912 1728 18964
rect 3332 18912 3384 18964
rect 2044 18844 2096 18896
rect 2228 18844 2280 18896
rect 5172 18912 5224 18964
rect 5540 18912 5592 18964
rect 5816 18912 5868 18964
rect 1584 18776 1636 18828
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1860 18708 1912 18760
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 4160 18708 4212 18760
rect 6736 18776 6788 18828
rect 6920 18776 6972 18828
rect 8392 18912 8444 18964
rect 8116 18844 8168 18896
rect 9588 18912 9640 18964
rect 10324 18955 10376 18964
rect 10324 18921 10333 18955
rect 10333 18921 10367 18955
rect 10367 18921 10376 18955
rect 10324 18912 10376 18921
rect 11888 18912 11940 18964
rect 4988 18708 5040 18760
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 2688 18572 2740 18624
rect 3792 18572 3844 18624
rect 4068 18572 4120 18624
rect 5264 18640 5316 18692
rect 4712 18615 4764 18624
rect 4712 18581 4721 18615
rect 4721 18581 4755 18615
rect 4755 18581 4764 18615
rect 4712 18572 4764 18581
rect 8208 18708 8260 18760
rect 8576 18776 8628 18828
rect 10784 18776 10836 18828
rect 6920 18683 6972 18692
rect 6920 18649 6929 18683
rect 6929 18649 6963 18683
rect 6963 18649 6972 18683
rect 6920 18640 6972 18649
rect 7932 18640 7984 18692
rect 8116 18640 8168 18692
rect 5724 18572 5776 18624
rect 5816 18572 5868 18624
rect 6828 18572 6880 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 8208 18615 8260 18624
rect 7012 18572 7064 18581
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 9588 18708 9640 18760
rect 9956 18751 10008 18760
rect 9956 18717 9965 18751
rect 9965 18717 9999 18751
rect 9999 18717 10008 18751
rect 9956 18708 10008 18717
rect 10048 18708 10100 18760
rect 10324 18708 10376 18760
rect 12624 18844 12676 18896
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 13728 18776 13780 18785
rect 18144 18776 18196 18828
rect 15476 18751 15528 18760
rect 9036 18572 9088 18624
rect 13452 18683 13504 18692
rect 13452 18649 13470 18683
rect 13470 18649 13504 18683
rect 13452 18640 13504 18649
rect 13636 18640 13688 18692
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 19064 18912 19116 18964
rect 19524 18912 19576 18964
rect 19984 18708 20036 18760
rect 21180 18708 21232 18760
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 12164 18572 12216 18624
rect 13084 18572 13136 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 17132 18640 17184 18692
rect 19708 18640 19760 18692
rect 17960 18572 18012 18624
rect 20444 18572 20496 18624
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 3240 18368 3292 18420
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 2320 18232 2372 18284
rect 2596 18232 2648 18284
rect 3240 18164 3292 18216
rect 3884 18368 3936 18420
rect 4528 18368 4580 18420
rect 4068 18275 4120 18284
rect 4068 18241 4077 18275
rect 4077 18241 4111 18275
rect 4111 18241 4120 18275
rect 4068 18232 4120 18241
rect 5264 18232 5316 18284
rect 6920 18368 6972 18420
rect 7840 18368 7892 18420
rect 5908 18300 5960 18352
rect 6184 18300 6236 18352
rect 6828 18300 6880 18352
rect 7196 18300 7248 18352
rect 7656 18343 7708 18352
rect 7656 18309 7665 18343
rect 7665 18309 7699 18343
rect 7699 18309 7708 18343
rect 7656 18300 7708 18309
rect 6000 18232 6052 18284
rect 8208 18368 8260 18420
rect 9496 18368 9548 18420
rect 12808 18368 12860 18420
rect 9036 18300 9088 18352
rect 13084 18300 13136 18352
rect 13544 18368 13596 18420
rect 14832 18300 14884 18352
rect 15660 18300 15712 18352
rect 4528 18207 4580 18216
rect 2872 18096 2924 18148
rect 4528 18173 4537 18207
rect 4537 18173 4571 18207
rect 4571 18173 4580 18207
rect 4528 18164 4580 18173
rect 6184 18164 6236 18216
rect 7472 18207 7524 18216
rect 5172 18096 5224 18148
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9496 18164 9548 18216
rect 10048 18164 10100 18216
rect 16212 18232 16264 18284
rect 20076 18368 20128 18420
rect 20996 18368 21048 18420
rect 21364 18411 21416 18420
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 19616 18300 19668 18352
rect 21640 18300 21692 18352
rect 17408 18232 17460 18284
rect 19432 18275 19484 18284
rect 19432 18241 19450 18275
rect 19450 18241 19484 18275
rect 19432 18232 19484 18241
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 20076 18232 20128 18284
rect 20628 18232 20680 18284
rect 18052 18207 18104 18216
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 3332 18028 3384 18080
rect 4712 18028 4764 18080
rect 5448 18028 5500 18080
rect 6368 18071 6420 18080
rect 6368 18037 6377 18071
rect 6377 18037 6411 18071
rect 6411 18037 6420 18071
rect 6368 18028 6420 18037
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 6828 18028 6880 18037
rect 7840 18096 7892 18148
rect 9680 18096 9732 18148
rect 11336 18096 11388 18148
rect 10048 18028 10100 18080
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 12900 18028 12952 18080
rect 13452 18028 13504 18080
rect 16212 18096 16264 18148
rect 14188 18028 14240 18080
rect 14280 18028 14332 18080
rect 17132 18028 17184 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1676 17824 1728 17876
rect 3424 17824 3476 17876
rect 4160 17824 4212 17876
rect 9680 17824 9732 17876
rect 10324 17824 10376 17876
rect 11244 17824 11296 17876
rect 3884 17756 3936 17808
rect 7196 17756 7248 17808
rect 11428 17756 11480 17808
rect 18052 17824 18104 17876
rect 19984 17824 20036 17876
rect 19432 17756 19484 17808
rect 19616 17799 19668 17808
rect 19616 17765 19625 17799
rect 19625 17765 19659 17799
rect 19659 17765 19668 17799
rect 19616 17756 19668 17765
rect 4068 17688 4120 17740
rect 4896 17688 4948 17740
rect 6828 17688 6880 17740
rect 8208 17688 8260 17740
rect 9680 17688 9732 17740
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 1952 17663 2004 17672
rect 1952 17629 1961 17663
rect 1961 17629 1995 17663
rect 1995 17629 2004 17663
rect 1952 17620 2004 17629
rect 3884 17620 3936 17672
rect 4528 17620 4580 17672
rect 7472 17620 7524 17672
rect 7288 17552 7340 17604
rect 9220 17620 9272 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 14188 17688 14240 17740
rect 17132 17688 17184 17740
rect 19708 17688 19760 17740
rect 11428 17552 11480 17604
rect 11796 17552 11848 17604
rect 12164 17552 12216 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2136 17527 2188 17536
rect 2136 17493 2145 17527
rect 2145 17493 2179 17527
rect 2179 17493 2188 17527
rect 2136 17484 2188 17493
rect 2412 17484 2464 17536
rect 2688 17484 2740 17536
rect 3608 17484 3660 17536
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 4528 17484 4580 17493
rect 4804 17484 4856 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6368 17484 6420 17536
rect 6828 17484 6880 17536
rect 7012 17484 7064 17536
rect 7932 17484 7984 17536
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 9036 17484 9088 17536
rect 11704 17527 11756 17536
rect 11704 17493 11713 17527
rect 11713 17493 11747 17527
rect 11747 17493 11756 17527
rect 11704 17484 11756 17493
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 12900 17484 12952 17536
rect 14004 17620 14056 17672
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 16212 17620 16264 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 14924 17552 14976 17604
rect 15568 17552 15620 17604
rect 20812 17552 20864 17604
rect 20996 17552 21048 17604
rect 14372 17484 14424 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 17684 17484 17736 17536
rect 19340 17484 19392 17536
rect 19524 17484 19576 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2320 17280 2372 17332
rect 3240 17323 3292 17332
rect 3240 17289 3249 17323
rect 3249 17289 3283 17323
rect 3283 17289 3292 17323
rect 3240 17280 3292 17289
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 4896 17280 4948 17332
rect 5356 17280 5408 17332
rect 5908 17280 5960 17332
rect 6552 17280 6604 17332
rect 7656 17280 7708 17332
rect 8944 17280 8996 17332
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 9680 17280 9732 17332
rect 11244 17280 11296 17332
rect 11704 17280 11756 17332
rect 12900 17280 12952 17332
rect 13268 17280 13320 17332
rect 13820 17280 13872 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 15476 17280 15528 17332
rect 13912 17212 13964 17264
rect 1768 17144 1820 17196
rect 2872 17144 2924 17196
rect 4160 17144 4212 17196
rect 4528 17144 4580 17196
rect 5816 17187 5868 17196
rect 3332 17076 3384 17128
rect 3792 17119 3844 17128
rect 3792 17085 3801 17119
rect 3801 17085 3835 17119
rect 3835 17085 3844 17119
rect 3792 17076 3844 17085
rect 2964 17008 3016 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6828 17144 6880 17196
rect 8576 17144 8628 17196
rect 10508 17144 10560 17196
rect 5172 17119 5224 17128
rect 5172 17085 5181 17119
rect 5181 17085 5215 17119
rect 5215 17085 5224 17119
rect 5172 17076 5224 17085
rect 5724 17076 5776 17128
rect 6552 17076 6604 17128
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 6644 17008 6696 17060
rect 5172 16940 5224 16992
rect 7564 17076 7616 17128
rect 14004 17144 14056 17196
rect 14188 17212 14240 17264
rect 16396 17212 16448 17264
rect 17040 17144 17092 17196
rect 18052 17212 18104 17264
rect 17684 17144 17736 17196
rect 18144 17144 18196 17196
rect 19064 17280 19116 17332
rect 19984 17280 20036 17332
rect 20996 17212 21048 17264
rect 19800 17144 19852 17196
rect 21364 17187 21416 17196
rect 21364 17153 21373 17187
rect 21373 17153 21407 17187
rect 21407 17153 21416 17187
rect 21364 17144 21416 17153
rect 7380 17008 7432 17060
rect 10784 17008 10836 17060
rect 11244 16940 11296 16992
rect 13728 17008 13780 17060
rect 15200 17008 15252 17060
rect 13820 16940 13872 16992
rect 15384 16940 15436 16992
rect 15476 16940 15528 16992
rect 16396 16940 16448 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 19340 17008 19392 17060
rect 20352 17008 20404 17060
rect 17960 16940 18012 16992
rect 18972 16983 19024 16992
rect 18972 16949 18981 16983
rect 18981 16949 19015 16983
rect 19015 16949 19024 16983
rect 18972 16940 19024 16949
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 19892 16940 19944 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1676 16736 1728 16788
rect 2872 16736 2924 16788
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 5080 16736 5132 16788
rect 4528 16668 4580 16720
rect 6000 16668 6052 16720
rect 7840 16736 7892 16788
rect 8760 16736 8812 16788
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 1952 16532 2004 16584
rect 2780 16532 2832 16584
rect 3240 16464 3292 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 1860 16396 1912 16448
rect 4068 16396 4120 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 7104 16396 7156 16448
rect 7840 16600 7892 16652
rect 7380 16532 7432 16584
rect 8116 16532 8168 16584
rect 9128 16600 9180 16652
rect 20076 16736 20128 16788
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 10968 16464 11020 16516
rect 12164 16668 12216 16720
rect 15476 16600 15528 16652
rect 19064 16600 19116 16652
rect 19708 16575 19760 16584
rect 13820 16464 13872 16516
rect 19708 16541 19731 16575
rect 19731 16541 19760 16575
rect 21088 16575 21140 16584
rect 19708 16532 19760 16541
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 9588 16439 9640 16448
rect 9588 16405 9597 16439
rect 9597 16405 9631 16439
rect 9631 16405 9640 16439
rect 9588 16396 9640 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 10324 16396 10376 16448
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 11888 16396 11940 16448
rect 12348 16396 12400 16448
rect 13544 16396 13596 16448
rect 16028 16507 16080 16516
rect 16028 16473 16062 16507
rect 16062 16473 16080 16507
rect 16028 16464 16080 16473
rect 15660 16396 15712 16448
rect 17224 16464 17276 16516
rect 17500 16439 17552 16448
rect 17500 16405 17509 16439
rect 17509 16405 17543 16439
rect 17543 16405 17552 16439
rect 17500 16396 17552 16405
rect 18236 16464 18288 16516
rect 20996 16464 21048 16516
rect 20812 16439 20864 16448
rect 20812 16405 20821 16439
rect 20821 16405 20855 16439
rect 20855 16405 20864 16439
rect 20812 16396 20864 16405
rect 20904 16396 20956 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 3332 16235 3384 16244
rect 2780 16192 2832 16201
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 3976 16192 4028 16244
rect 5540 16235 5592 16244
rect 5540 16201 5549 16235
rect 5549 16201 5583 16235
rect 5583 16201 5592 16235
rect 5540 16192 5592 16201
rect 6000 16192 6052 16244
rect 6736 16192 6788 16244
rect 7012 16192 7064 16244
rect 7196 16192 7248 16244
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 9220 16192 9272 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 6828 16124 6880 16176
rect 8024 16124 8076 16176
rect 3332 16056 3384 16108
rect 4528 16099 4580 16108
rect 4528 16065 4537 16099
rect 4537 16065 4571 16099
rect 4571 16065 4580 16099
rect 4528 16056 4580 16065
rect 4068 15988 4120 16040
rect 4160 15988 4212 16040
rect 5080 15988 5132 16040
rect 5724 16056 5776 16108
rect 2044 15963 2096 15972
rect 2044 15929 2053 15963
rect 2053 15929 2087 15963
rect 2087 15929 2096 15963
rect 2044 15920 2096 15929
rect 3884 15920 3936 15972
rect 5448 15920 5500 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4988 15852 5040 15904
rect 5632 15852 5684 15904
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 6000 15920 6052 15972
rect 8116 16056 8168 16108
rect 8668 16056 8720 16108
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 7656 15920 7708 15972
rect 15108 16124 15160 16176
rect 15476 16192 15528 16244
rect 16304 16235 16356 16244
rect 16304 16201 16313 16235
rect 16313 16201 16347 16235
rect 16347 16201 16356 16235
rect 16304 16192 16356 16201
rect 20352 16192 20404 16244
rect 17408 16124 17460 16176
rect 18972 16124 19024 16176
rect 12992 16056 13044 16108
rect 15476 16056 15528 16108
rect 15016 15988 15068 16040
rect 17500 16056 17552 16108
rect 17776 16099 17828 16108
rect 17776 16065 17794 16099
rect 17794 16065 17828 16099
rect 17776 16056 17828 16065
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 19892 16056 19944 16108
rect 13544 15920 13596 15972
rect 6092 15852 6144 15904
rect 10416 15852 10468 15904
rect 13176 15895 13228 15904
rect 13176 15861 13185 15895
rect 13185 15861 13219 15895
rect 13219 15861 13228 15895
rect 16028 15920 16080 15972
rect 21088 15920 21140 15972
rect 13176 15852 13228 15861
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 15108 15852 15160 15904
rect 15936 15852 15988 15904
rect 19984 15852 20036 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2596 15648 2648 15700
rect 3332 15648 3384 15700
rect 3516 15648 3568 15700
rect 4620 15648 4672 15700
rect 6092 15648 6144 15700
rect 7656 15648 7708 15700
rect 1768 15580 1820 15632
rect 5448 15580 5500 15632
rect 8208 15648 8260 15700
rect 9404 15648 9456 15700
rect 9680 15648 9732 15700
rect 20720 15648 20772 15700
rect 5632 15512 5684 15564
rect 7196 15512 7248 15564
rect 13452 15580 13504 15632
rect 15568 15580 15620 15632
rect 18880 15623 18932 15632
rect 8300 15512 8352 15564
rect 1860 15444 1912 15496
rect 1952 15444 2004 15496
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3424 15444 3476 15496
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5540 15444 5592 15496
rect 8116 15444 8168 15496
rect 8576 15444 8628 15496
rect 10416 15487 10468 15496
rect 4160 15419 4212 15428
rect 4160 15385 4169 15419
rect 4169 15385 4203 15419
rect 4203 15385 4212 15419
rect 4160 15376 4212 15385
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 3516 15308 3568 15360
rect 5448 15308 5500 15360
rect 6736 15376 6788 15428
rect 7840 15376 7892 15428
rect 8668 15376 8720 15428
rect 8760 15376 8812 15428
rect 9496 15376 9548 15428
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 8116 15351 8168 15360
rect 7012 15308 7064 15317
rect 8116 15317 8125 15351
rect 8125 15317 8159 15351
rect 8159 15317 8168 15351
rect 8116 15308 8168 15317
rect 10324 15308 10376 15360
rect 10508 15308 10560 15360
rect 16304 15444 16356 15496
rect 18880 15589 18889 15623
rect 18889 15589 18923 15623
rect 18923 15589 18932 15623
rect 18880 15580 18932 15589
rect 19064 15580 19116 15632
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 14188 15376 14240 15428
rect 15016 15376 15068 15428
rect 16396 15376 16448 15428
rect 20812 15376 20864 15428
rect 21088 15419 21140 15428
rect 21088 15385 21106 15419
rect 21106 15385 21140 15419
rect 21088 15376 21140 15385
rect 15568 15308 15620 15360
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 18604 15308 18656 15360
rect 18972 15308 19024 15360
rect 19708 15351 19760 15360
rect 19708 15317 19717 15351
rect 19717 15317 19751 15351
rect 19751 15317 19760 15351
rect 19708 15308 19760 15317
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1676 15104 1728 15156
rect 2596 15147 2648 15156
rect 2596 15113 2605 15147
rect 2605 15113 2639 15147
rect 2639 15113 2648 15147
rect 2596 15104 2648 15113
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 6000 15147 6052 15156
rect 6000 15113 6009 15147
rect 6009 15113 6043 15147
rect 6043 15113 6052 15147
rect 6000 15104 6052 15113
rect 6736 15104 6788 15156
rect 6920 15104 6972 15156
rect 7104 15104 7156 15156
rect 9864 15104 9916 15156
rect 1768 14968 1820 15020
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 4160 15036 4212 15088
rect 4712 15036 4764 15088
rect 3884 14968 3936 15020
rect 3976 14900 4028 14952
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 2596 14832 2648 14884
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 5540 14900 5592 14952
rect 5908 14900 5960 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 7748 15036 7800 15088
rect 9680 15036 9732 15088
rect 10876 15104 10928 15156
rect 14188 15104 14240 15156
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 17500 15104 17552 15156
rect 7656 14968 7708 15020
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11244 14968 11296 15020
rect 5448 14832 5500 14884
rect 8300 14900 8352 14952
rect 9312 14943 9364 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 5264 14764 5316 14816
rect 6828 14764 6880 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 7932 14832 7984 14884
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 12992 14900 13044 14952
rect 9404 14764 9456 14816
rect 15108 15036 15160 15088
rect 19432 15104 19484 15156
rect 14832 14968 14884 15020
rect 15200 14968 15252 15020
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 17960 15011 18012 15020
rect 17960 14977 17978 15011
rect 17978 14977 18012 15011
rect 19984 15104 20036 15156
rect 19708 15079 19760 15088
rect 19708 15045 19717 15079
rect 19717 15045 19751 15079
rect 19751 15045 19760 15079
rect 19708 15036 19760 15045
rect 17960 14968 18012 14977
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18880 15011 18932 15020
rect 18236 14968 18288 14977
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 14280 14900 14332 14952
rect 15016 14900 15068 14952
rect 14188 14832 14240 14884
rect 15292 14832 15344 14884
rect 13820 14764 13872 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15016 14764 15068 14816
rect 16948 14764 17000 14816
rect 21364 15011 21416 15020
rect 21364 14977 21373 15011
rect 21373 14977 21407 15011
rect 21407 14977 21416 15011
rect 21364 14968 21416 14977
rect 19892 14764 19944 14816
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 2228 14560 2280 14612
rect 3148 14560 3200 14612
rect 3516 14560 3568 14612
rect 3976 14603 4028 14612
rect 3976 14569 3985 14603
rect 3985 14569 4019 14603
rect 4019 14569 4028 14603
rect 3976 14560 4028 14569
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 6000 14560 6052 14612
rect 6644 14560 6696 14612
rect 6828 14603 6880 14612
rect 6828 14569 6837 14603
rect 6837 14569 6871 14603
rect 6871 14569 6880 14603
rect 6828 14560 6880 14569
rect 7472 14560 7524 14612
rect 7656 14603 7708 14612
rect 7656 14569 7665 14603
rect 7665 14569 7699 14603
rect 7699 14569 7708 14603
rect 7656 14560 7708 14569
rect 8484 14560 8536 14612
rect 9312 14560 9364 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 2688 14492 2740 14544
rect 4344 14492 4396 14544
rect 10876 14492 10928 14544
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 5540 14424 5592 14476
rect 6552 14424 6604 14476
rect 6920 14424 6972 14476
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 3148 14356 3200 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4712 14356 4764 14408
rect 2412 14288 2464 14340
rect 7564 14356 7616 14408
rect 8392 14424 8444 14476
rect 10508 14424 10560 14476
rect 12440 14424 12492 14476
rect 16304 14560 16356 14612
rect 17040 14560 17092 14612
rect 18236 14603 18288 14612
rect 18236 14569 18245 14603
rect 18245 14569 18279 14603
rect 18279 14569 18288 14603
rect 18236 14560 18288 14569
rect 19708 14560 19760 14612
rect 16948 14492 17000 14544
rect 13820 14356 13872 14408
rect 15108 14356 15160 14408
rect 21364 14424 21416 14476
rect 19892 14356 19944 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 2964 14263 3016 14272
rect 2964 14229 2973 14263
rect 2973 14229 3007 14263
rect 3007 14229 3016 14263
rect 2964 14220 3016 14229
rect 14280 14288 14332 14340
rect 14372 14288 14424 14340
rect 15292 14288 15344 14340
rect 5632 14220 5684 14272
rect 6828 14220 6880 14272
rect 9680 14220 9732 14272
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 11980 14220 12032 14272
rect 14556 14220 14608 14272
rect 17684 14331 17736 14340
rect 17684 14297 17702 14331
rect 17702 14297 17736 14331
rect 17684 14288 17736 14297
rect 19800 14288 19852 14340
rect 18512 14220 18564 14272
rect 19064 14220 19116 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 3332 14016 3384 14068
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 5816 14016 5868 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 8116 14016 8168 14068
rect 9220 14016 9272 14068
rect 9680 14016 9732 14068
rect 9772 14016 9824 14068
rect 1584 13880 1636 13932
rect 2320 13855 2372 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 6000 13948 6052 14000
rect 10784 13948 10836 14000
rect 12808 13948 12860 14000
rect 15016 14016 15068 14068
rect 3516 13880 3568 13932
rect 4068 13880 4120 13932
rect 4160 13880 4212 13932
rect 8300 13880 8352 13932
rect 12532 13880 12584 13932
rect 6092 13812 6144 13864
rect 6552 13812 6604 13864
rect 4620 13744 4672 13796
rect 5172 13744 5224 13796
rect 5540 13744 5592 13796
rect 7840 13812 7892 13864
rect 10324 13855 10376 13864
rect 6828 13744 6880 13796
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 14740 13948 14792 14000
rect 16396 14016 16448 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 17224 14016 17276 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 18512 14016 18564 14068
rect 20996 14016 21048 14068
rect 9220 13744 9272 13796
rect 2964 13676 3016 13728
rect 5264 13676 5316 13728
rect 8484 13676 8536 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 13360 13676 13412 13728
rect 15292 13812 15344 13864
rect 16488 13812 16540 13864
rect 16764 13880 16816 13932
rect 21088 13948 21140 14000
rect 18512 13923 18564 13932
rect 18512 13889 18530 13923
rect 18530 13889 18564 13923
rect 18512 13880 18564 13889
rect 18880 13880 18932 13932
rect 20352 13880 20404 13932
rect 20904 13880 20956 13932
rect 21364 14016 21416 14068
rect 17592 13812 17644 13864
rect 15200 13744 15252 13796
rect 15660 13744 15712 13796
rect 18788 13744 18840 13796
rect 18972 13744 19024 13796
rect 14924 13676 14976 13728
rect 16028 13676 16080 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2320 13472 2372 13524
rect 3884 13472 3936 13524
rect 4528 13472 4580 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 9220 13472 9272 13524
rect 9496 13472 9548 13524
rect 2504 13404 2556 13456
rect 2780 13336 2832 13388
rect 4620 13404 4672 13456
rect 5816 13447 5868 13456
rect 5816 13413 5825 13447
rect 5825 13413 5859 13447
rect 5859 13413 5868 13447
rect 5816 13404 5868 13413
rect 9312 13404 9364 13456
rect 12164 13404 12216 13456
rect 19524 13472 19576 13524
rect 15200 13404 15252 13456
rect 15384 13404 15436 13456
rect 16948 13404 17000 13456
rect 19616 13404 19668 13456
rect 3884 13336 3936 13388
rect 4068 13336 4120 13388
rect 4436 13336 4488 13388
rect 4804 13336 4856 13388
rect 6092 13336 6144 13388
rect 6736 13336 6788 13388
rect 8208 13336 8260 13388
rect 11152 13336 11204 13388
rect 11888 13336 11940 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 4344 13268 4396 13320
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 6828 13268 6880 13320
rect 4068 13200 4120 13252
rect 4528 13200 4580 13252
rect 9312 13200 9364 13252
rect 10416 13200 10468 13252
rect 10968 13200 11020 13252
rect 2964 13132 3016 13184
rect 3884 13132 3936 13184
rect 5540 13132 5592 13184
rect 6828 13175 6880 13184
rect 6828 13141 6837 13175
rect 6837 13141 6871 13175
rect 6871 13141 6880 13175
rect 6828 13132 6880 13141
rect 7472 13132 7524 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 16028 13336 16080 13388
rect 17408 13336 17460 13388
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 13820 13268 13872 13320
rect 14832 13268 14884 13320
rect 16488 13268 16540 13320
rect 14004 13200 14056 13252
rect 19064 13268 19116 13320
rect 21456 13268 21508 13320
rect 13360 13132 13412 13184
rect 19340 13200 19392 13252
rect 19984 13200 20036 13252
rect 20076 13200 20128 13252
rect 20812 13200 20864 13252
rect 14556 13132 14608 13184
rect 15016 13132 15068 13184
rect 20352 13132 20404 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3332 12928 3384 12980
rect 4068 12928 4120 12980
rect 6000 12928 6052 12980
rect 7288 12928 7340 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 13820 12928 13872 12980
rect 14924 12928 14976 12980
rect 2044 12792 2096 12844
rect 3056 12724 3108 12776
rect 1400 12699 1452 12708
rect 1400 12665 1409 12699
rect 1409 12665 1443 12699
rect 1443 12665 1452 12699
rect 1400 12656 1452 12665
rect 4068 12656 4120 12708
rect 4436 12860 4488 12912
rect 4620 12792 4672 12844
rect 6276 12792 6328 12844
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 5264 12724 5316 12776
rect 8576 12860 8628 12912
rect 8392 12792 8444 12844
rect 8484 12792 8536 12844
rect 13544 12860 13596 12912
rect 14372 12792 14424 12844
rect 14832 12792 14884 12844
rect 9588 12724 9640 12776
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 15936 12860 15988 12912
rect 16764 12860 16816 12912
rect 17408 12860 17460 12912
rect 18880 12928 18932 12980
rect 19340 12971 19392 12980
rect 19340 12937 19349 12971
rect 19349 12937 19383 12971
rect 19383 12937 19392 12971
rect 19340 12928 19392 12937
rect 19800 12971 19852 12980
rect 19800 12937 19809 12971
rect 19809 12937 19843 12971
rect 19843 12937 19852 12971
rect 19800 12928 19852 12937
rect 20904 12928 20956 12980
rect 19616 12792 19668 12844
rect 21364 12792 21416 12844
rect 4712 12588 4764 12640
rect 5632 12588 5684 12640
rect 8208 12588 8260 12640
rect 9128 12588 9180 12640
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 15016 12588 15068 12640
rect 19524 12588 19576 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 4160 12384 4212 12436
rect 5908 12384 5960 12436
rect 2872 12316 2924 12368
rect 3608 12316 3660 12368
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 4804 12316 4856 12368
rect 8300 12384 8352 12436
rect 9956 12384 10008 12436
rect 11980 12384 12032 12436
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 4344 12180 4396 12232
rect 5356 12248 5408 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 6920 12248 6972 12300
rect 7104 12180 7156 12232
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 17316 12384 17368 12436
rect 18880 12427 18932 12436
rect 18880 12393 18889 12427
rect 18889 12393 18923 12427
rect 18923 12393 18932 12427
rect 18880 12384 18932 12393
rect 10784 12248 10836 12300
rect 12532 12248 12584 12300
rect 16304 12316 16356 12368
rect 16764 12359 16816 12368
rect 16764 12325 16773 12359
rect 16773 12325 16807 12359
rect 16807 12325 16816 12359
rect 16764 12316 16816 12325
rect 10324 12180 10376 12232
rect 11060 12180 11112 12232
rect 11980 12180 12032 12232
rect 21364 12291 21416 12300
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 14832 12180 14884 12232
rect 16304 12180 16356 12232
rect 5080 12112 5132 12164
rect 1952 12044 2004 12096
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 5724 12044 5776 12096
rect 7288 12044 7340 12096
rect 9404 12044 9456 12096
rect 11796 12112 11848 12164
rect 15292 12155 15344 12164
rect 15292 12121 15326 12155
rect 15326 12121 15344 12155
rect 15292 12112 15344 12121
rect 11152 12044 11204 12096
rect 12072 12044 12124 12096
rect 13544 12044 13596 12096
rect 15476 12044 15528 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 17868 12044 17920 12096
rect 21272 12112 21324 12164
rect 18788 12044 18840 12096
rect 18972 12044 19024 12096
rect 19616 12087 19668 12096
rect 19616 12053 19625 12087
rect 19625 12053 19659 12087
rect 19659 12053 19668 12087
rect 19616 12044 19668 12053
rect 20536 12044 20588 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1860 11840 1912 11892
rect 1216 11772 1268 11824
rect 4896 11840 4948 11892
rect 7380 11840 7432 11892
rect 7840 11840 7892 11892
rect 8208 11840 8260 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 10968 11840 11020 11892
rect 13452 11840 13504 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 15936 11883 15988 11892
rect 15936 11849 15945 11883
rect 15945 11849 15979 11883
rect 15979 11849 15988 11883
rect 15936 11840 15988 11849
rect 17040 11840 17092 11892
rect 17684 11883 17736 11892
rect 17684 11849 17693 11883
rect 17693 11849 17727 11883
rect 17727 11849 17736 11883
rect 17684 11840 17736 11849
rect 19524 11840 19576 11892
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 16396 11772 16448 11824
rect 18880 11772 18932 11824
rect 7380 11704 7432 11756
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 11796 11704 11848 11756
rect 12072 11704 12124 11756
rect 12624 11704 12676 11756
rect 13360 11704 13412 11756
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 14464 11704 14516 11756
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 17408 11704 17460 11756
rect 18788 11747 18840 11756
rect 20536 11772 20588 11824
rect 18788 11713 18806 11747
rect 18806 11713 18840 11747
rect 18788 11704 18840 11713
rect 21364 11704 21416 11756
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 4436 11568 4488 11620
rect 5356 11568 5408 11620
rect 6736 11636 6788 11688
rect 10968 11636 11020 11688
rect 12440 11636 12492 11688
rect 14188 11636 14240 11688
rect 6920 11568 6972 11620
rect 1308 11500 1360 11552
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 4988 11500 5040 11509
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 13084 11500 13136 11552
rect 13728 11500 13780 11552
rect 14740 11500 14792 11552
rect 17500 11500 17552 11552
rect 19708 11500 19760 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1676 11296 1728 11348
rect 2596 11339 2648 11348
rect 2596 11305 2605 11339
rect 2605 11305 2639 11339
rect 2639 11305 2648 11339
rect 2596 11296 2648 11305
rect 3240 11296 3292 11348
rect 5448 11296 5500 11348
rect 7288 11296 7340 11348
rect 8668 11296 8720 11348
rect 11704 11296 11756 11348
rect 14464 11296 14516 11348
rect 15476 11339 15528 11348
rect 4528 11228 4580 11280
rect 6000 11228 6052 11280
rect 11980 11228 12032 11280
rect 12532 11228 12584 11280
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 5540 11160 5592 11212
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 12624 11160 12676 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2780 11092 2832 11144
rect 4988 11092 5040 11144
rect 6736 11092 6788 11144
rect 7104 11092 7156 11144
rect 10048 11092 10100 11144
rect 11888 11092 11940 11144
rect 13820 11160 13872 11212
rect 15108 11160 15160 11212
rect 17684 11296 17736 11348
rect 19432 11296 19484 11348
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 17408 11160 17460 11212
rect 18880 11160 18932 11212
rect 14188 11092 14240 11144
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 19708 11092 19760 11144
rect 4068 11024 4120 11076
rect 4252 11024 4304 11076
rect 4988 10956 5040 11008
rect 10508 11024 10560 11076
rect 13084 11024 13136 11076
rect 5632 10956 5684 11008
rect 7656 10956 7708 11008
rect 8116 10956 8168 11008
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 10692 10956 10744 11008
rect 12440 10956 12492 11008
rect 12624 10956 12676 11008
rect 16856 11067 16908 11076
rect 16856 11033 16874 11067
rect 16874 11033 16908 11067
rect 16856 11024 16908 11033
rect 17224 11024 17276 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1400 10752 1452 10804
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 3424 10752 3476 10804
rect 4068 10752 4120 10804
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 10232 10752 10284 10804
rect 12992 10795 13044 10804
rect 12992 10761 13001 10795
rect 13001 10761 13035 10795
rect 13035 10761 13044 10795
rect 12992 10752 13044 10761
rect 13268 10752 13320 10804
rect 13820 10752 13872 10804
rect 18420 10752 18472 10804
rect 20076 10752 20128 10804
rect 1492 10616 1544 10668
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 8484 10684 8536 10736
rect 10140 10684 10192 10736
rect 13452 10684 13504 10736
rect 17040 10684 17092 10736
rect 19432 10727 19484 10736
rect 19432 10693 19450 10727
rect 19450 10693 19484 10727
rect 19432 10684 19484 10693
rect 19616 10684 19668 10736
rect 4160 10616 4212 10668
rect 5908 10616 5960 10668
rect 7748 10616 7800 10668
rect 9496 10616 9548 10668
rect 13084 10616 13136 10668
rect 13820 10616 13872 10668
rect 14280 10616 14332 10668
rect 2688 10548 2740 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 7472 10548 7524 10600
rect 9128 10548 9180 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 12072 10548 12124 10600
rect 1676 10480 1728 10532
rect 1860 10480 1912 10532
rect 7012 10480 7064 10532
rect 7380 10523 7432 10532
rect 7380 10489 7389 10523
rect 7389 10489 7423 10523
rect 7423 10489 7432 10523
rect 7380 10480 7432 10489
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 8300 10412 8352 10464
rect 9128 10412 9180 10464
rect 11060 10412 11112 10464
rect 12348 10412 12400 10464
rect 16304 10616 16356 10668
rect 21088 10659 21140 10668
rect 21088 10625 21106 10659
rect 21106 10625 21140 10659
rect 21364 10659 21416 10668
rect 21088 10616 21140 10625
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 14832 10412 14884 10464
rect 17316 10412 17368 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1768 10208 1820 10260
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 4988 10208 5040 10260
rect 5448 10208 5500 10260
rect 6000 10208 6052 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 7748 10208 7800 10260
rect 10600 10208 10652 10260
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 11244 10208 11296 10260
rect 1492 10140 1544 10192
rect 7196 10140 7248 10192
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5448 10072 5500 10124
rect 7288 10115 7340 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 5816 10004 5868 10056
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 8576 10004 8628 10056
rect 6736 9936 6788 9988
rect 9588 10140 9640 10192
rect 12624 10140 12676 10192
rect 13820 10208 13872 10260
rect 11060 10072 11112 10124
rect 14280 10072 14332 10124
rect 18788 10208 18840 10260
rect 21088 10208 21140 10260
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 12532 10004 12584 10056
rect 15384 10004 15436 10056
rect 16028 10004 16080 10056
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 18052 10004 18104 10056
rect 21364 10004 21416 10056
rect 1860 9868 1912 9920
rect 7104 9868 7156 9920
rect 8208 9911 8260 9920
rect 8208 9877 8217 9911
rect 8217 9877 8251 9911
rect 8251 9877 8260 9911
rect 8208 9868 8260 9877
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 9128 9868 9180 9920
rect 9680 9868 9732 9920
rect 10784 9868 10836 9920
rect 12440 9868 12492 9920
rect 14832 9868 14884 9920
rect 15292 9868 15344 9920
rect 16948 9936 17000 9988
rect 18696 9868 18748 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 8300 9664 8352 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 10968 9664 11020 9716
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 21364 9707 21416 9716
rect 4620 9596 4672 9648
rect 7104 9639 7156 9648
rect 7104 9605 7113 9639
rect 7113 9605 7147 9639
rect 7147 9605 7156 9639
rect 7104 9596 7156 9605
rect 7472 9596 7524 9648
rect 7932 9596 7984 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2228 9435 2280 9444
rect 2228 9401 2237 9435
rect 2237 9401 2271 9435
rect 2271 9401 2280 9435
rect 2228 9392 2280 9401
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 4528 9528 4580 9580
rect 7380 9528 7432 9580
rect 9588 9528 9640 9580
rect 12440 9596 12492 9648
rect 16028 9596 16080 9648
rect 17132 9596 17184 9648
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 9036 9503 9088 9512
rect 5908 9392 5960 9444
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 9680 9392 9732 9444
rect 10600 9392 10652 9444
rect 13268 9571 13320 9580
rect 13268 9537 13286 9571
rect 13286 9537 13320 9571
rect 13268 9528 13320 9537
rect 13820 9528 13872 9580
rect 14280 9528 14332 9580
rect 18052 9528 18104 9580
rect 3424 9324 3476 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 7288 9324 7340 9376
rect 7932 9324 7984 9376
rect 10692 9324 10744 9376
rect 10968 9324 11020 9376
rect 19708 9460 19760 9512
rect 15844 9435 15896 9444
rect 15844 9401 15853 9435
rect 15853 9401 15887 9435
rect 15887 9401 15896 9435
rect 15844 9392 15896 9401
rect 16948 9392 17000 9444
rect 19340 9392 19392 9444
rect 20536 9435 20588 9444
rect 20536 9401 20545 9435
rect 20545 9401 20579 9435
rect 20579 9401 20588 9435
rect 20536 9392 20588 9401
rect 13176 9324 13228 9376
rect 19524 9324 19576 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1584 9120 1636 9172
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 1492 9052 1544 9104
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3424 8916 3476 8968
rect 5724 9120 5776 9172
rect 7012 9120 7064 9172
rect 8024 9120 8076 9172
rect 9588 9163 9640 9172
rect 9588 9129 9597 9163
rect 9597 9129 9631 9163
rect 9631 9129 9640 9163
rect 9588 9120 9640 9129
rect 9680 9120 9732 9172
rect 10692 9120 10744 9172
rect 5448 9052 5500 9104
rect 7656 9052 7708 9104
rect 10968 9052 11020 9104
rect 13820 9120 13872 9172
rect 16028 9163 16080 9172
rect 16028 9129 16037 9163
rect 16037 9129 16071 9163
rect 16071 9129 16080 9163
rect 16028 9120 16080 9129
rect 21364 9120 21416 9172
rect 6460 8984 6512 9036
rect 6644 8984 6696 9036
rect 9864 8984 9916 9036
rect 17868 9052 17920 9104
rect 18696 9052 18748 9104
rect 6000 8916 6052 8968
rect 12808 8984 12860 9036
rect 13728 8916 13780 8968
rect 6920 8780 6972 8832
rect 9404 8780 9456 8832
rect 9588 8780 9640 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2136 8576 2188 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 8208 8576 8260 8628
rect 9404 8619 9456 8628
rect 9404 8585 9413 8619
rect 9413 8585 9447 8619
rect 9447 8585 9456 8619
rect 9404 8576 9456 8585
rect 9496 8576 9548 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 10968 8576 11020 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 21088 8576 21140 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 8668 8508 8720 8560
rect 12164 8508 12216 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 7104 8440 7156 8492
rect 8392 8440 8444 8492
rect 8576 8440 8628 8492
rect 9588 8440 9640 8492
rect 10692 8440 10744 8492
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7564 8372 7616 8424
rect 8300 8372 8352 8424
rect 9312 8372 9364 8424
rect 10048 8372 10100 8424
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 5632 8304 5684 8356
rect 10876 8304 10928 8356
rect 11980 8304 12032 8356
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 11888 8236 11940 8288
rect 13176 8372 13228 8424
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 6000 8075 6052 8084
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 7196 8032 7248 8084
rect 8668 8032 8720 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 11060 8032 11112 8084
rect 5172 7964 5224 8016
rect 8300 7964 8352 8016
rect 9220 7964 9272 8016
rect 6368 7896 6420 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 7932 7939 7984 7948
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 9496 7896 9548 7948
rect 12716 7939 12768 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 7840 7760 7892 7812
rect 8024 7760 8076 7812
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 11888 7828 11940 7880
rect 7012 7692 7064 7744
rect 7196 7692 7248 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 19892 7760 19944 7812
rect 11152 7692 11204 7744
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2596 7488 2648 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7932 7488 7984 7540
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 9496 7531 9548 7540
rect 9496 7497 9505 7531
rect 9505 7497 9539 7531
rect 9539 7497 9548 7531
rect 9496 7488 9548 7497
rect 10324 7420 10376 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 8300 7352 8352 7404
rect 8484 7352 8536 7404
rect 9128 7352 9180 7404
rect 5172 7216 5224 7268
rect 5816 7148 5868 7200
rect 6736 7148 6788 7200
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 9496 7284 9548 7336
rect 10232 7148 10284 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 1400 6944 1452 6996
rect 7564 6944 7616 6996
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 7012 6740 7064 6792
rect 9404 6944 9456 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 8208 6808 8260 6860
rect 10232 6808 10284 6860
rect 18604 6808 18656 6860
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 5356 6672 5408 6724
rect 6920 6604 6972 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 11060 6604 11112 6656
rect 15568 6672 15620 6724
rect 15936 6604 15988 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 5356 6400 5408 6452
rect 7564 6400 7616 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 5816 6264 5868 6316
rect 10232 6443 10284 6452
rect 10232 6409 10241 6443
rect 10241 6409 10275 6443
rect 10275 6409 10284 6443
rect 10232 6400 10284 6409
rect 11060 6400 11112 6452
rect 12256 6400 12308 6452
rect 7196 6196 7248 6248
rect 10692 6332 10744 6384
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 4068 6060 4120 6112
rect 8300 6128 8352 6180
rect 10232 6196 10284 6248
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 8208 6060 8260 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1400 5856 1452 5908
rect 2044 5856 2096 5908
rect 10968 5856 11020 5908
rect 7656 5788 7708 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 10968 5287 11020 5296
rect 10968 5253 10977 5287
rect 10977 5253 11011 5287
rect 11011 5253 11020 5287
rect 10968 5244 11020 5253
rect 16212 5244 16264 5296
rect 7380 5176 7432 5228
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 4988 4632 5040 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 7012 4020 7064 4072
rect 10876 3952 10928 4004
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1492 3680 1544 3732
rect 4068 3612 4120 3664
rect 1492 3451 1544 3460
rect 1492 3417 1501 3451
rect 1501 3417 1535 3451
rect 1535 3417 1544 3451
rect 1492 3408 1544 3417
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 5816 3136 5868 3188
rect 5540 3068 5592 3120
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 7932 2524 7984 2576
rect 7196 2456 7248 2508
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 2780 2320 2832 2372
rect 11704 2252 11756 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3528 22222 3832 22250
rect 216 20466 244 22200
rect 204 20460 256 20466
rect 204 20402 256 20408
rect 676 19922 704 22200
rect 664 19916 716 19922
rect 664 19858 716 19864
rect 1136 19310 1164 22200
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 1228 11830 1256 19858
rect 1216 11824 1268 11830
rect 1216 11766 1268 11772
rect 1320 11558 1348 20402
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1490 18864 1546 18873
rect 1596 18834 1624 22200
rect 2056 21434 2084 22200
rect 2056 21406 2268 21434
rect 2042 21312 2098 21321
rect 2042 21247 2098 21256
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1688 18970 1716 19314
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1490 18799 1546 18808
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1688 17882 1716 18226
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1688 16794 1716 17614
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1490 16759 1546 16768
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1688 15162 1716 16050
rect 1780 15638 1808 17138
rect 1872 16454 1900 18702
rect 1964 18426 1992 19314
rect 2056 18902 2084 21247
rect 2134 19272 2190 19281
rect 2134 19207 2136 19216
rect 2188 19207 2190 19216
rect 2136 19178 2188 19184
rect 2240 18902 2268 21406
rect 2516 19938 2544 22200
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2516 19910 2636 19938
rect 2700 19922 2728 20334
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2792 20097 2820 20198
rect 2778 20088 2834 20097
rect 2778 20023 2834 20032
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2044 18896 2096 18902
rect 2044 18838 2096 18844
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2134 17640 2190 17649
rect 1964 17338 1992 17614
rect 2134 17575 2190 17584
rect 2148 17542 2176 17575
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2332 17338 2360 18226
rect 2424 17542 2452 19722
rect 2516 19514 2544 19790
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2608 18306 2636 19910
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2780 19712 2832 19718
rect 2778 19680 2780 19689
rect 2832 19680 2834 19689
rect 2778 19615 2834 19624
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2516 18290 2636 18306
rect 2516 18284 2648 18290
rect 2516 18278 2596 18284
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1964 15706 1992 16526
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2042 16008 2098 16017
rect 2042 15943 2044 15952
rect 2096 15943 2098 15952
rect 2044 15914 2096 15920
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1490 15127 1546 15136
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13569 1532 13670
rect 1490 13560 1546 13569
rect 1490 13495 1546 13504
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 13161 1440 13262
rect 1398 13152 1454 13161
rect 1398 13087 1454 13096
rect 1398 12744 1454 12753
rect 1398 12679 1400 12688
rect 1452 12679 1454 12688
rect 1400 12650 1452 12656
rect 1412 12238 1440 12650
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1398 11928 1454 11937
rect 1398 11863 1454 11872
rect 1412 11762 1440 11863
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1308 11552 1360 11558
rect 1308 11494 1360 11500
rect 1398 11520 1454 11529
rect 1398 11455 1454 11464
rect 1412 11150 1440 11455
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1490 11112 1546 11121
rect 1412 10810 1440 11086
rect 1490 11047 1546 11056
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1504 10674 1532 11047
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1412 10062 1440 10231
rect 1504 10198 1532 10610
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1412 9602 1440 9823
rect 1412 9586 1532 9602
rect 1400 9580 1532 9586
rect 1452 9574 1532 9580
rect 1400 9522 1452 9528
rect 1398 9480 1454 9489
rect 1398 9415 1454 9424
rect 1412 8974 1440 9415
rect 1504 9110 1532 9574
rect 1596 9178 1624 13874
rect 1688 11354 1716 14350
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1674 10840 1730 10849
rect 1674 10775 1730 10784
rect 1688 10538 1716 10775
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1780 10266 1808 14962
rect 1872 11898 1900 15438
rect 1964 12986 1992 15438
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2042 14376 2098 14385
rect 2042 14311 2098 14320
rect 2056 14278 2084 14311
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12345 2084 12786
rect 2148 12442 2176 14962
rect 2240 14618 2268 16050
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2042 12336 2098 12345
rect 2042 12271 2098 12280
rect 1950 12200 2006 12209
rect 1950 12135 2006 12144
rect 1964 12102 1992 12135
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1872 9926 1900 10474
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1412 8498 1440 8735
rect 1858 8664 1914 8673
rect 1858 8599 1914 8608
rect 1872 8498 1900 8599
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1412 7886 1440 8191
rect 2056 8090 2084 10610
rect 2134 10024 2190 10033
rect 2134 9959 2190 9968
rect 2148 8634 2176 9959
rect 2240 9450 2268 14350
rect 2424 14346 2452 14962
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2332 13530 2360 13806
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2516 13462 2544 18278
rect 2596 18226 2648 18232
rect 2700 17660 2728 18566
rect 2884 18154 2912 19314
rect 2976 18850 3004 22200
rect 3436 20618 3464 22200
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3252 20590 3464 20618
rect 3160 20505 3188 20538
rect 3146 20496 3202 20505
rect 3146 20431 3202 20440
rect 3252 19378 3280 20590
rect 3528 20482 3556 22222
rect 3804 22114 3832 22222
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8588 22222 8892 22250
rect 3896 22114 3924 22200
rect 3804 22086 3924 22114
rect 3974 20904 4030 20913
rect 3974 20839 4030 20848
rect 3988 20602 4016 20839
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3436 20454 3556 20482
rect 3884 20460 3936 20466
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 2976 18822 3096 18850
rect 3068 18766 3096 18822
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2608 17632 2728 17660
rect 2608 15706 2636 17632
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15162 2636 15438
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2318 12336 2374 12345
rect 2318 12271 2374 12280
rect 2332 12238 2360 12271
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2608 11354 2636 14826
rect 2700 14550 2728 17478
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16794 2912 17138
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2792 16250 2820 16526
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2976 15162 3004 17002
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2700 13818 2728 14486
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2700 13790 2820 13818
rect 2792 13394 2820 13790
rect 2976 13734 3004 14214
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2976 13444 3004 13670
rect 2884 13416 3004 13444
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2884 12374 2912 13416
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2976 12306 3004 13126
rect 3068 12986 3096 18702
rect 3160 14618 3188 19110
rect 3252 18426 3280 19314
rect 3344 18970 3372 20402
rect 3436 19836 3464 20454
rect 3884 20402 3936 20408
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3516 19848 3568 19854
rect 3436 19808 3516 19836
rect 3516 19790 3568 19796
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 19553 3464 19654
rect 3422 19544 3478 19553
rect 3422 19479 3478 19488
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3252 17338 3280 18158
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3344 17218 3372 18022
rect 3436 17882 3464 19314
rect 3528 19281 3556 19790
rect 3514 19272 3570 19281
rect 3514 19207 3570 19216
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3804 18170 3832 18566
rect 3896 18426 3924 20402
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3804 18142 3924 18170
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3896 17814 3924 18142
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17338 3648 17478
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3790 17232 3846 17241
rect 3344 17190 3464 17218
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3240 16516 3292 16522
rect 3240 16458 3292 16464
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3068 12238 3096 12718
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2792 10713 2820 11086
rect 3160 10810 3188 14350
rect 3252 11354 3280 16458
rect 3344 16250 3372 17070
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15706 3372 16050
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15586 3464 17190
rect 3790 17167 3846 17176
rect 3804 17134 3832 17167
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3896 15978 3924 17614
rect 3988 16250 4016 19654
rect 4080 18630 4108 19751
rect 4356 19378 4384 22200
rect 4816 20482 4844 22200
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4632 20454 4844 20482
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4172 18766 4200 19178
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4080 17898 4108 18226
rect 4080 17882 4200 17898
rect 4080 17876 4212 17882
rect 4080 17870 4160 17876
rect 4160 17818 4212 17824
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4080 16538 4108 17682
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4172 16794 4200 17138
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4080 16510 4200 16538
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4080 16046 4108 16390
rect 4172 16046 4200 16510
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3344 15558 3464 15586
rect 3344 14074 3372 15558
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3344 12986 3372 14010
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3436 10810 3464 15438
rect 3528 15366 3556 15642
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 15065 3556 15302
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3528 13938 3556 14554
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3896 13530 3924 14962
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14618 4016 14894
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4080 14498 4108 15982
rect 4158 15464 4214 15473
rect 4158 15399 4160 15408
rect 4212 15399 4214 15408
rect 4160 15370 4212 15376
rect 4172 15094 4200 15370
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3988 14470 4108 14498
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3896 13190 3924 13330
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3620 11694 3648 12310
rect 3988 11801 4016 14470
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4080 13394 4108 13874
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12986 4108 13194
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4080 12306 4108 12650
rect 4172 12442 4200 13874
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3608 11688 3660 11694
rect 3606 11656 3608 11665
rect 3660 11656 3662 11665
rect 3606 11591 3662 11600
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 4264 11082 4292 19110
rect 4356 14550 4384 19314
rect 4448 16153 4476 19790
rect 4540 19446 4568 20402
rect 4632 19854 4660 20454
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4540 18426 4568 19246
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4540 17678 4568 18158
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4540 17338 4568 17478
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4540 16726 4568 17138
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4434 16144 4490 16153
rect 4434 16079 4490 16088
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4436 14952 4488 14958
rect 4434 14920 4436 14929
rect 4488 14920 4490 14929
rect 4434 14855 4490 14864
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 13326 4384 14350
rect 4448 13394 4476 14418
rect 4540 13530 4568 16050
rect 4632 15706 4660 19790
rect 4724 18630 4752 20334
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4816 19378 4844 20266
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 5000 18766 5028 19450
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4724 15094 4752 18022
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4816 16658 4844 17478
rect 4908 17338 4936 17682
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 16561 4844 16594
rect 4802 16552 4858 16561
rect 4802 16487 4858 16496
rect 4908 15881 4936 17274
rect 5092 16794 5120 20198
rect 5276 19922 5304 22200
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 19514 5396 19654
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5460 19174 5488 20402
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 19417 5580 20198
rect 5538 19408 5594 19417
rect 5538 19343 5594 19352
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5184 18766 5212 18906
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 18290 5304 18634
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5184 17134 5212 18090
rect 5172 17128 5224 17134
rect 5170 17096 5172 17105
rect 5224 17096 5226 17105
rect 5170 17031 5226 17040
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4988 15904 5040 15910
rect 4894 15872 4950 15881
rect 4988 15846 5040 15852
rect 4894 15807 4950 15816
rect 5000 15502 5028 15846
rect 4988 15496 5040 15502
rect 4894 15464 4950 15473
rect 4988 15438 5040 15444
rect 4894 15399 4950 15408
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 14074 4660 14418
rect 4724 14414 4752 15030
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4620 14068 4672 14074
rect 4672 14028 4844 14056
rect 4620 14010 4672 14016
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4632 13462 4660 13738
rect 4620 13456 4672 13462
rect 4618 13424 4620 13433
rect 4672 13424 4674 13433
rect 4436 13388 4488 13394
rect 4674 13382 4752 13410
rect 4816 13394 4844 14028
rect 4618 13359 4674 13368
rect 4436 13330 4488 13336
rect 4632 13333 4660 13359
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4356 12238 4384 12718
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4448 11626 4476 12854
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4540 11286 4568 13194
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4080 10810 4108 11018
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 2688 10600 2740 10606
rect 2686 10568 2688 10577
rect 2740 10568 2742 10577
rect 2686 10503 2742 10512
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 4172 10266 4200 10610
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4632 9654 4660 12786
rect 4724 12646 4752 13382
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4804 12368 4856 12374
rect 4908 12322 4936 15399
rect 4856 12316 4936 12322
rect 4804 12310 4936 12316
rect 4816 12294 4936 12310
rect 4908 11898 4936 12294
rect 5092 12170 5120 15982
rect 5184 13920 5212 16934
rect 5276 14822 5304 18226
rect 5368 17338 5396 19110
rect 5460 18086 5488 19110
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5552 16250 5580 18906
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 15638 5488 15914
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5552 15502 5580 16186
rect 5644 15910 5672 20538
rect 5736 19378 5764 22200
rect 6196 20890 6224 22200
rect 6012 20862 6224 20890
rect 6012 20482 6040 20862
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6656 20618 6684 22200
rect 6564 20590 6684 20618
rect 7116 20602 7144 22200
rect 7104 20596 7156 20602
rect 6012 20454 6224 20482
rect 6564 20466 6592 20590
rect 7104 20538 7156 20544
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7288 20528 7340 20534
rect 6642 20496 6698 20505
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5736 18850 5764 19314
rect 5828 18970 5856 19654
rect 5908 19440 5960 19446
rect 6012 19417 6040 20198
rect 6104 19990 6132 20334
rect 6196 20262 6224 20454
rect 6552 20460 6604 20466
rect 7288 20470 7340 20476
rect 6642 20431 6698 20440
rect 6736 20460 6788 20466
rect 6552 20402 6604 20408
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6196 19854 6224 20198
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6380 19786 6408 19926
rect 6550 19816 6606 19825
rect 6368 19780 6420 19786
rect 6550 19751 6552 19760
rect 6368 19722 6420 19728
rect 6604 19751 6606 19760
rect 6552 19722 6604 19728
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6656 19514 6684 20431
rect 6736 20402 6788 20408
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 5908 19382 5960 19388
rect 5998 19408 6054 19417
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5736 18822 5856 18850
rect 5828 18630 5856 18822
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5736 17134 5764 18566
rect 5920 18358 5948 19382
rect 5998 19343 6054 19352
rect 6104 19310 6132 19450
rect 6368 19440 6420 19446
rect 6366 19408 6368 19417
rect 6460 19440 6512 19446
rect 6420 19408 6422 19417
rect 6460 19382 6512 19388
rect 6550 19408 6606 19417
rect 6366 19343 6422 19352
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6472 18873 6500 19382
rect 6550 19343 6606 19352
rect 6644 19372 6696 19378
rect 6458 18864 6514 18873
rect 6458 18799 6514 18808
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17338 5948 17478
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6012 17218 6040 18226
rect 6196 18222 6224 18294
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6380 17542 6408 18022
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6564 17338 6592 19343
rect 6644 19314 6696 19320
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5920 17190 6040 17218
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16114 5764 16390
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5354 14920 5410 14929
rect 5460 14890 5488 15302
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5354 14855 5410 14864
rect 5448 14884 5500 14890
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5368 14618 5396 14855
rect 5448 14826 5500 14832
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5552 14482 5580 14894
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5644 14362 5672 15506
rect 5552 14334 5672 14362
rect 5184 13892 5304 13920
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5184 12889 5212 13738
rect 5276 13734 5304 13892
rect 5552 13802 5580 14334
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5262 13016 5318 13025
rect 5262 12951 5318 12960
rect 5170 12880 5226 12889
rect 5170 12815 5226 12824
rect 5276 12782 5304 12951
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5368 12306 5396 13262
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 11150 5028 11494
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10266 5028 10950
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1400 7880 1452 7886
rect 1860 7880 1912 7886
rect 1400 7822 1452 7828
rect 1858 7848 1860 7857
rect 1912 7848 1914 7857
rect 1858 7783 1914 7792
rect 2608 7546 2636 9522
rect 2792 9081 2820 9522
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 3436 8974 3464 9318
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 4540 9178 4568 9522
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 1398 7440 1454 7449
rect 1398 7375 1400 7384
rect 1452 7375 1454 7384
rect 1860 7404 1912 7410
rect 1400 7346 1452 7352
rect 1860 7346 1912 7352
rect 1412 7002 1440 7346
rect 1872 7041 1900 7346
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 1858 7032 1914 7041
rect 3549 7035 3857 7044
rect 1400 6996 1452 7002
rect 1858 6967 1914 6976
rect 1400 6938 1452 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6633 1440 6734
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1412 6225 1440 6258
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 1412 5914 1440 6151
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1872 5817 1900 6258
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 2056 5914 2084 6054
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5409 1440 5646
rect 1398 5400 1454 5409
rect 1398 5335 1454 5344
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2240 5001 2268 5102
rect 2226 4992 2282 5001
rect 2226 4927 2282 4936
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 2228 4616 2280 4622
rect 2226 4584 2228 4593
rect 2280 4584 2282 4593
rect 2226 4519 2282 4528
rect 1490 4176 1546 4185
rect 1490 4111 1492 4120
rect 1544 4111 1546 4120
rect 2044 4140 2096 4146
rect 1492 4082 1544 4088
rect 2044 4082 2096 4088
rect 1504 3738 1532 4082
rect 2056 3777 2084 4082
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 2042 3768 2098 3777
rect 3549 3771 3857 3780
rect 1492 3732 1544 3738
rect 2042 3703 2098 3712
rect 1492 3674 1544 3680
rect 4080 3670 4108 6054
rect 5000 4690 5028 10202
rect 5184 8022 5212 12038
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 11121 5396 11562
rect 5460 11354 5488 11630
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11218 5580 13126
rect 5644 12646 5672 14214
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5630 12472 5686 12481
rect 5630 12407 5686 12416
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5354 11112 5410 11121
rect 5644 11098 5672 12407
rect 5736 12209 5764 16050
rect 5828 14074 5856 17138
rect 5920 15042 5948 17190
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 16250 6040 16662
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 15162 6040 15914
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 15706 6132 15846
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 5920 15014 6040 15042
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5814 13968 5870 13977
rect 5814 13903 5870 13912
rect 5828 13462 5856 13903
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5920 13002 5948 14894
rect 6012 14618 6040 15014
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6564 14482 6592 17070
rect 6656 17066 6684 19314
rect 6748 18834 6776 20402
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6840 18714 6868 20198
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 6932 19446 6960 19926
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6918 18864 6974 18873
rect 6918 18799 6920 18808
rect 6972 18799 6974 18808
rect 6920 18770 6972 18776
rect 6748 18686 6868 18714
rect 6920 18692 6972 18698
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6748 16946 6776 18686
rect 6920 18634 6972 18640
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18358 6868 18566
rect 6932 18426 6960 18634
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6840 17785 6868 18022
rect 6826 17776 6882 17785
rect 6826 17711 6828 17720
rect 6880 17711 6882 17720
rect 6828 17682 6880 17688
rect 6840 17651 6868 17682
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 17202 6868 17478
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6656 16918 6776 16946
rect 6656 14618 6684 16918
rect 6840 16266 6868 17138
rect 6932 16402 6960 18362
rect 7024 18057 7052 18566
rect 7010 18048 7066 18057
rect 7010 17983 7066 17992
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 17134 7052 17478
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7116 16538 7144 19246
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7208 17814 7236 18294
rect 7300 18170 7328 20470
rect 7392 19242 7420 20538
rect 7576 19904 7604 22200
rect 8036 20534 8064 22200
rect 8496 20806 8524 22200
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8588 20618 8616 22222
rect 8864 22114 8892 22222
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 16868 22222 17080 22250
rect 8956 22114 8984 22200
rect 8864 22086 8984 22114
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8220 20590 8616 20618
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8220 20466 8248 20590
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 7748 20392 7800 20398
rect 8024 20392 8076 20398
rect 7800 20352 8024 20380
rect 7748 20334 7800 20340
rect 8024 20334 8076 20340
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7576 19876 7696 19904
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7484 19514 7512 19654
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7576 19446 7604 19654
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7472 18216 7524 18222
rect 7470 18184 7472 18193
rect 7524 18184 7526 18193
rect 7300 18142 7420 18170
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7194 17232 7250 17241
rect 7194 17167 7250 17176
rect 7208 16658 7236 17167
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7116 16510 7236 16538
rect 7104 16448 7156 16454
rect 6932 16374 7052 16402
rect 7104 16390 7156 16396
rect 6736 16244 6788 16250
rect 6840 16238 6960 16266
rect 7024 16250 7052 16374
rect 6736 16186 6788 16192
rect 6748 15434 6776 16186
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6550 14240 6606 14249
rect 6148 14172 6456 14181
rect 6550 14175 6606 14184
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5828 12974 5948 13002
rect 6012 12986 6040 13942
rect 6564 13870 6592 14175
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6104 13394 6132 13806
rect 6748 13512 6776 15098
rect 6840 14822 6868 16118
rect 6932 15688 6960 16238
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7012 16040 7064 16046
rect 7010 16008 7012 16017
rect 7064 16008 7066 16017
rect 7010 15943 7066 15952
rect 6932 15660 7052 15688
rect 7024 15450 7052 15660
rect 6932 15422 7052 15450
rect 6932 15162 6960 15422
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6826 14648 6882 14657
rect 6826 14583 6828 14592
rect 6880 14583 6882 14592
rect 6828 14554 6880 14560
rect 6840 14278 6868 14554
rect 6932 14482 6960 14894
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6656 13484 6776 13512
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6656 13297 6684 13484
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6642 13288 6698 13297
rect 6642 13223 6698 13232
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6000 12980 6052 12986
rect 5828 12730 5856 12974
rect 6000 12922 6052 12928
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5828 12702 5948 12730
rect 5920 12442 5948 12702
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6288 12306 6316 12786
rect 6656 12481 6684 13223
rect 6642 12472 6698 12481
rect 6642 12407 6698 12416
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 5722 12200 5778 12209
rect 5722 12135 5778 12144
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5354 11047 5410 11056
rect 5552 11070 5672 11098
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5262 10160 5318 10169
rect 5460 10130 5488 10202
rect 5262 10095 5264 10104
rect 5316 10095 5318 10104
rect 5448 10124 5500 10130
rect 5264 10066 5316 10072
rect 5448 10066 5500 10072
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8634 5488 9046
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5184 6730 5212 7210
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 6458 5396 6666
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1504 3369 1532 3402
rect 1490 3360 1546 3369
rect 1490 3295 1546 3304
rect 5552 3126 5580 11070
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 8362 5672 10950
rect 5736 9178 5764 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6642 11928 6698 11937
rect 6642 11863 6698 11872
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 6182 11248 6238 11257
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10062 5856 10406
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5920 9450 5948 10610
rect 6012 10266 6040 11222
rect 6182 11183 6184 11192
rect 6236 11183 6238 11192
rect 6184 11154 6236 11160
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 6472 9042 6500 9318
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 6012 8090 6040 8910
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8537 6592 10542
rect 6656 9602 6684 11863
rect 6748 11694 6776 13330
rect 6840 13326 6868 13738
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10810 6776 11086
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6840 10266 6868 13126
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6932 11626 6960 12242
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 7024 10538 7052 15302
rect 7116 15162 7144 16390
rect 7208 16250 7236 16510
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7194 15600 7250 15609
rect 7194 15535 7196 15544
rect 7248 15535 7250 15544
rect 7196 15506 7248 15512
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14074 7236 14962
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7300 12986 7328 17546
rect 7392 17066 7420 18142
rect 7470 18119 7526 18128
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7104 12232 7156 12238
rect 7102 12200 7104 12209
rect 7156 12200 7158 12209
rect 7102 12135 7158 12144
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11354 7328 12038
rect 7392 11898 7420 16526
rect 7484 16266 7512 17614
rect 7576 17134 7604 19246
rect 7668 19174 7696 19876
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7668 17338 7696 18294
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7484 16238 7604 16266
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7484 14618 7512 16079
rect 7576 14929 7604 16238
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7668 15706 7696 15914
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7760 15094 7788 20198
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8036 19854 8064 19994
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7852 18426 7880 19110
rect 7944 18698 7972 19654
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7852 16794 7880 18090
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7838 16688 7894 16697
rect 7838 16623 7840 16632
rect 7892 16623 7894 16632
rect 7840 16594 7892 16600
rect 7944 16250 7972 17478
rect 8036 16266 8064 19790
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 8128 18902 8156 19246
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8220 18766 8248 20402
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8128 16590 8156 18634
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18426 8248 18566
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17649 8248 17682
rect 8206 17640 8262 17649
rect 8206 17575 8262 17584
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 16244 7984 16250
rect 8036 16238 8156 16266
rect 7932 16186 7984 16192
rect 8024 16176 8076 16182
rect 7838 16144 7894 16153
rect 8024 16118 8076 16124
rect 7838 16079 7894 16088
rect 7852 15881 7880 16079
rect 7838 15872 7894 15881
rect 7838 15807 7894 15816
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7748 15088 7800 15094
rect 7654 15056 7710 15065
rect 7748 15030 7800 15036
rect 7654 14991 7656 15000
rect 7708 14991 7710 15000
rect 7656 14962 7708 14968
rect 7562 14920 7618 14929
rect 7562 14855 7618 14864
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14414 7604 14758
rect 7668 14618 7696 14962
rect 7746 14920 7802 14929
rect 7746 14855 7802 14864
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12434 7512 13126
rect 7484 12406 7604 12434
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7116 10033 7144 11086
rect 7392 10538 7420 11698
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7286 10296 7342 10305
rect 7286 10231 7342 10240
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7102 10024 7158 10033
rect 6736 9988 6788 9994
rect 7102 9959 7158 9968
rect 6736 9930 6788 9936
rect 6748 9722 6776 9930
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 7116 9654 7144 9862
rect 7104 9648 7156 9654
rect 6656 9574 6776 9602
rect 7104 9590 7156 9596
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6550 8528 6606 8537
rect 6550 8463 6606 8472
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6380 7954 6408 8230
rect 6656 7954 6684 8978
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6656 7546 6684 7890
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6748 7206 6776 9574
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6826 8936 6882 8945
rect 6826 8871 6882 8880
rect 6840 8634 6868 8871
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 5828 6322 5856 7142
rect 5908 6792 5960 6798
rect 5906 6760 5908 6769
rect 5960 6760 5962 6769
rect 5906 6695 5962 6704
rect 6932 6662 6960 8774
rect 7024 8430 7052 9114
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7116 7970 7144 8434
rect 7208 8090 7236 10134
rect 7300 10130 7328 10231
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7484 9654 7512 10542
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 9382 7328 9454
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7392 8634 7420 9522
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7484 8514 7512 9590
rect 7392 8486 7512 8514
rect 7576 8514 7604 12406
rect 7668 11014 7696 14554
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7760 10826 7788 14855
rect 7852 14793 7880 15370
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7838 14784 7894 14793
rect 7838 14719 7894 14728
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13530 7880 13806
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7668 10798 7788 10826
rect 7668 9110 7696 10798
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 10266 7788 10610
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7576 8486 7696 8514
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7116 7942 7236 7970
rect 7208 7750 7236 7942
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7024 7546 7052 7686
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5828 3194 5856 6258
rect 7024 6118 7052 6734
rect 7208 6254 7236 7686
rect 7392 6662 7420 8486
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 7342 7604 8366
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 7002 7604 7278
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 7024 4078 7052 6054
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1504 2961 1532 2994
rect 1490 2952 1546 2961
rect 1490 2887 1546 2896
rect 2056 2553 2084 2994
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 2042 2544 2098 2553
rect 7208 2514 7236 6190
rect 7392 5234 7420 6598
rect 7576 6458 7604 6938
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7668 5846 7696 8486
rect 7746 7984 7802 7993
rect 7746 7919 7748 7928
rect 7800 7919 7802 7928
rect 7748 7890 7800 7896
rect 7852 7818 7880 11834
rect 7944 9654 7972 14826
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 7954 7972 9318
rect 8036 9178 8064 16118
rect 8128 16114 8156 16238
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8128 15502 8156 16050
rect 8208 15700 8260 15706
rect 8312 15688 8340 20198
rect 8404 18970 8432 20402
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19553 8524 20198
rect 8482 19544 8538 19553
rect 8482 19479 8538 19488
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8312 15660 8432 15688
rect 8208 15642 8260 15648
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 14074 8156 15302
rect 8220 14385 8248 15642
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 14958 8340 15506
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8298 14784 8354 14793
rect 8298 14719 8354 14728
rect 8206 14376 8262 14385
rect 8206 14311 8262 14320
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 13394 8248 14311
rect 8312 13938 8340 14719
rect 8404 14482 8432 15660
rect 8496 14618 8524 19314
rect 8588 19310 8616 20402
rect 8680 20330 8708 20742
rect 9416 20602 9444 22200
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20602 9720 20742
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9876 20534 9904 22200
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 9128 20256 9180 20262
rect 9312 20256 9364 20262
rect 9180 20216 9260 20244
rect 9128 20198 9180 20204
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8680 19514 8708 19994
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18329 8616 18770
rect 8574 18320 8630 18329
rect 8574 18255 8630 18264
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17202 8616 17478
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8680 16114 8708 19178
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18358 9076 18566
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8956 17338 8984 17478
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9048 17105 9076 17478
rect 9140 17338 9168 19790
rect 9232 19174 9260 20216
rect 9312 20198 9364 20204
rect 9324 19394 9352 20198
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9416 19786 9444 19926
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9402 19544 9458 19553
rect 9402 19479 9404 19488
rect 9456 19479 9458 19488
rect 9404 19450 9456 19456
rect 9324 19366 9444 19394
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9034 17096 9090 17105
rect 9034 17031 9090 17040
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8576 16040 8628 16046
rect 8772 15994 8800 16730
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8576 15982 8628 15988
rect 8588 15502 8616 15982
rect 8680 15966 8800 15994
rect 8680 15688 8708 15966
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8680 15660 8800 15688
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8496 12850 8524 13670
rect 8588 12918 8616 15438
rect 8772 15434 8800 15660
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 11898 8248 12582
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8128 8514 8156 10950
rect 8312 10470 8340 12378
rect 8404 12306 8432 12786
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8496 10826 8524 12786
rect 8680 11354 8708 15370
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9140 13977 9168 16594
rect 9232 16250 9260 17614
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9232 14074 9260 16186
rect 9324 15314 9352 19246
rect 9416 18465 9444 19366
rect 9402 18456 9458 18465
rect 9508 18426 9536 19790
rect 9600 18970 9628 20402
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 20097 9812 20198
rect 9770 20088 9826 20097
rect 9770 20023 9826 20032
rect 9680 19984 9732 19990
rect 9678 19952 9680 19961
rect 9732 19952 9734 19961
rect 9678 19887 9734 19896
rect 9678 19816 9734 19825
rect 9678 19751 9734 19760
rect 9692 19446 9720 19751
rect 9876 19514 9904 20295
rect 9968 20058 9996 20470
rect 10336 20466 10364 22200
rect 10796 20466 10824 22200
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9402 18391 9458 18400
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9416 15706 9444 18226
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9508 15434 9536 18158
rect 9600 16454 9628 18702
rect 9692 18154 9720 19246
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9692 17746 9720 17818
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17338 9720 17682
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9784 16674 9812 19178
rect 9692 16646 9812 16674
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9692 15706 9720 16646
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9324 15286 9720 15314
rect 9692 15094 9720 15286
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14618 9352 14894
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9220 14068 9272 14074
rect 9272 14028 9352 14056
rect 9220 14010 9272 14016
rect 9126 13968 9182 13977
rect 9126 13903 9182 13912
rect 9126 13832 9182 13841
rect 9126 13767 9182 13776
rect 9220 13796 9272 13802
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9140 12986 9168 13767
rect 9220 13738 9272 13744
rect 9232 13530 9260 13738
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9324 13462 9352 14028
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9324 13258 9352 13398
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8404 10798 8524 10826
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8404 10010 8432 10798
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10130 8524 10678
rect 9140 10606 9168 12582
rect 9416 12434 9444 14758
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 14074 9720 14214
rect 9784 14074 9812 16526
rect 9876 15162 9904 19314
rect 10060 18766 10088 19858
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9232 12406 9444 12434
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8576 10056 8628 10062
rect 8404 9982 8524 10010
rect 8576 9998 8628 10004
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8220 8634 8248 9862
rect 8312 9722 8340 9862
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8128 8486 8248 8514
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7944 7546 7972 7890
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 8036 2774 8064 7754
rect 8220 6866 8248 8486
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 8022 8340 8366
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8404 7546 8432 8434
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7410 8524 9982
rect 8588 8498 8616 9998
rect 9140 9926 9168 10406
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9512 9088 9518
rect 9034 9480 9036 9489
rect 9088 9480 9090 9489
rect 9034 9415 9090 9424
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8680 8090 8708 8502
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9232 8022 9260 12406
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9416 12102 9444 12135
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9508 11218 9536 13466
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10062 9352 10542
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8634 9444 8774
rect 9508 8634 9536 10610
rect 9600 10198 9628 12718
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9692 9926 9720 14010
rect 9862 13968 9918 13977
rect 9862 13903 9918 13912
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9178 9628 9522
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 9178 9720 9386
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9876 9042 9904 13903
rect 9968 12442 9996 18702
rect 10048 18216 10100 18222
rect 10046 18184 10048 18193
rect 10100 18184 10102 18193
rect 10046 18119 10102 18128
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 16590 10088 18022
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10152 16250 10180 19790
rect 10244 16454 10272 19790
rect 10336 18970 10364 20402
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 20058 10640 20266
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10428 19514 10456 19926
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 17882 10364 18702
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10336 16114 10364 16390
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10428 15994 10456 19207
rect 10520 17202 10548 19654
rect 10598 19136 10654 19145
rect 10598 19071 10654 19080
rect 10612 18737 10640 19071
rect 10598 18728 10654 18737
rect 10598 18663 10654 18672
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10336 15966 10456 15994
rect 10336 15366 10364 15966
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15502 10456 15846
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15026 10548 15302
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10138 14512 10194 14521
rect 10138 14447 10194 14456
rect 10508 14476 10560 14482
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 10046 11928 10102 11937
rect 10046 11863 10102 11872
rect 10060 11762 10088 11863
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11150 10088 11698
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10152 10742 10180 14447
rect 10508 14418 10560 14424
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10336 12238 10364 13806
rect 10414 13288 10470 13297
rect 10414 13223 10416 13232
rect 10468 13223 10470 13232
rect 10416 13194 10468 13200
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10520 11082 10548 14418
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10810 10272 10950
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10612 10266 10640 17614
rect 10704 11218 10732 20198
rect 10796 19514 10824 20402
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10980 19417 11008 20198
rect 10966 19408 11022 19417
rect 10966 19343 11022 19352
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10796 18834 10824 19246
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10966 17912 11022 17921
rect 10966 17847 11022 17856
rect 10980 17377 11008 17847
rect 10966 17368 11022 17377
rect 10966 17303 11022 17312
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10796 14396 10824 17002
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16250 10916 16390
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 14550 10916 15098
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10796 14368 10916 14396
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14006 10824 14214
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10888 13852 10916 14368
rect 10980 14249 11008 16458
rect 10966 14240 11022 14249
rect 10966 14175 11022 14184
rect 10796 13824 10916 13852
rect 10796 12306 10824 13824
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10888 11898 10916 13126
rect 10980 12050 11008 13194
rect 11072 12238 11100 20538
rect 11256 20466 11284 22200
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11716 20466 11744 22200
rect 12176 20466 12204 22200
rect 12636 20466 12664 22200
rect 13096 20602 13124 22200
rect 13556 20618 13584 22200
rect 13556 20602 13860 20618
rect 13084 20596 13136 20602
rect 13556 20596 13872 20602
rect 13556 20590 13820 20596
rect 13084 20538 13136 20544
rect 13820 20538 13872 20544
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 11256 20058 11284 20402
rect 11716 20058 11744 20402
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11150 18456 11206 18465
rect 11150 18391 11206 18400
rect 11164 13394 11192 18391
rect 11256 17882 11284 19790
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11900 18970 11928 19654
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11978 18728 12034 18737
rect 11978 18663 12034 18672
rect 11992 18630 12020 18663
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11348 17762 11376 18090
rect 11992 17921 12020 18566
rect 11978 17912 12034 17921
rect 11978 17847 12034 17856
rect 11256 17734 11376 17762
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11256 17338 11284 17734
rect 11440 17610 11468 17750
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17338 11744 17478
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 15144 11284 16934
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11702 16008 11758 16017
rect 11702 15943 11758 15952
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11256 15116 11376 15144
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14618 11284 14962
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11348 14498 11376 15116
rect 11256 14470 11376 14498
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11152 12096 11204 12102
rect 10980 12022 11100 12050
rect 11152 12038 11204 12044
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10980 11694 11008 11834
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 11072 11506 11100 12022
rect 10980 11478 11100 11506
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10266 10732 10950
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10048 9512 10100 9518
rect 10704 9466 10732 10202
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9722 10824 9862
rect 10980 9722 11008 11478
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10130 11100 10406
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10048 9454 10100 9460
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 8498 9628 8774
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 10060 8430 10088 9454
rect 10612 9450 10732 9466
rect 10600 9444 10732 9450
rect 10652 9438 10732 9444
rect 10600 9386 10652 9392
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9178 10732 9318
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10796 8514 10824 9658
rect 10980 9382 11008 9658
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9110 11008 9318
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10874 8664 10930 8673
rect 10980 8634 11008 9046
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10874 8599 10876 8608
rect 10928 8599 10930 8608
rect 10968 8628 11020 8634
rect 10876 8570 10928 8576
rect 10968 8570 11020 8576
rect 10966 8528 11022 8537
rect 10692 8492 10744 8498
rect 10796 8486 10916 8514
rect 10692 8434 10744 8440
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9324 7886 9352 8366
rect 10060 8090 10088 8366
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6118 8248 6802
rect 8312 6186 8340 7346
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9140 6458 9168 7346
rect 9416 7002 9444 7686
rect 9508 7546 9536 7890
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9508 7342 9536 7482
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 10244 6866 10272 7142
rect 10336 7002 10364 7414
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10244 6458 10272 6802
rect 10704 6662 10732 8434
rect 10888 8362 10916 8486
rect 10966 8463 11022 8472
rect 10980 8430 11008 8463
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10244 6254 10272 6394
rect 10704 6390 10732 6598
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 10888 4010 10916 8298
rect 11072 8090 11100 8774
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7750 11192 12038
rect 11256 10266 11284 14470
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 12345 11560 12922
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11716 11354 11744 15943
rect 11808 12170 11836 17546
rect 11978 16688 12034 16697
rect 11978 16623 12034 16632
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16250 11928 16390
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11992 14278 12020 16623
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11808 11121 11836 11698
rect 11900 11150 11928 13330
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12442 12020 12718
rect 11980 12436 12032 12442
rect 12084 12434 12112 20198
rect 12176 20058 12204 20402
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 17610 12204 18566
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12164 16720 12216 16726
rect 12162 16688 12164 16697
rect 12216 16688 12218 16697
rect 12162 16623 12218 16632
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13462 12204 13670
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 12782 12204 13398
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12084 12406 12204 12434
rect 11980 12378 12032 12384
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11286 12020 12174
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11762 12112 12038
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11888 11144 11940 11150
rect 11794 11112 11850 11121
rect 11888 11086 11940 11092
rect 11794 11047 11850 11056
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6458 11100 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10980 5302 11008 5850
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 7944 2746 8064 2774
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 7944 2582 7972 2746
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 2042 2479 2098 2488
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 11808 2446 11836 11047
rect 12084 10606 12112 11494
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8362 12020 8774
rect 12176 8566 12204 12406
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7886 11928 8230
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 7750 11928 7822
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 12268 6458 12296 20198
rect 12636 20058 12664 20402
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 16454 12388 17478
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 10470 12388 16390
rect 12452 14482 12480 19110
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12636 17377 12664 18838
rect 12622 17368 12678 17377
rect 12622 17303 12678 17312
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 12306 12572 13874
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12440 11688 12492 11694
rect 12492 11636 12572 11642
rect 12440 11630 12572 11636
rect 12452 11614 12572 11630
rect 12544 11286 12572 11614
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12452 9926 12480 10950
rect 12544 10062 12572 11222
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10198 12664 10950
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 8634 12480 9590
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12728 7954 12756 20198
rect 12898 20088 12954 20097
rect 12898 20023 12900 20032
rect 12952 20023 12954 20032
rect 12900 19994 12952 20000
rect 12912 19825 12940 19994
rect 12898 19816 12954 19825
rect 12898 19751 12954 19760
rect 13280 19689 13308 20402
rect 14016 20330 14044 22200
rect 14476 20602 14504 22200
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13266 19680 13322 19689
rect 13266 19615 13322 19624
rect 13740 19378 13768 19722
rect 14384 19718 14412 20470
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12820 18426 12848 19246
rect 13556 19145 13584 19314
rect 13636 19168 13688 19174
rect 13542 19136 13598 19145
rect 13636 19110 13688 19116
rect 13542 19071 13598 19080
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 13096 18358 13124 18566
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12912 17542 12940 18022
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17338 12940 17478
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12990 16144 13046 16153
rect 12990 16079 12992 16088
rect 13044 16079 13046 16088
rect 12992 16050 13044 16056
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12820 9042 12848 13942
rect 13004 10810 13032 14894
rect 13096 11558 13124 18294
rect 13464 18086 13492 18634
rect 13556 18426 13584 19071
rect 13648 18698 13676 19110
rect 13740 18834 13768 19314
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13726 18320 13782 18329
rect 13726 18255 13782 18264
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13096 10674 13124 11018
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13188 9382 13216 15846
rect 13280 11257 13308 17274
rect 13464 15638 13492 18022
rect 13740 17066 13768 18255
rect 13832 17338 13860 19450
rect 14660 19446 14688 20402
rect 14936 20330 14964 22200
rect 15198 20496 15254 20505
rect 15198 20431 15200 20440
rect 15252 20431 15254 20440
rect 15200 20402 15252 20408
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 15396 20058 15424 22200
rect 15856 20602 15884 22200
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16316 20330 16344 22200
rect 16776 22114 16804 22200
rect 16868 22114 16896 22222
rect 16776 22086 16896 22114
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 17052 20602 17080 22222
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 16776 19990 16804 20402
rect 17236 20262 17264 22200
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17512 20058 17540 20266
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15212 19514 15240 19654
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14476 18170 14504 19314
rect 15488 19174 15516 19654
rect 15764 19514 15792 19722
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18766 15516 19110
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 14832 18352 14884 18358
rect 14832 18294 14884 18300
rect 14200 18142 14504 18170
rect 14200 18086 14228 18142
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13910 17368 13966 17377
rect 13820 17332 13872 17338
rect 14016 17338 14044 17614
rect 13910 17303 13966 17312
rect 14004 17332 14056 17338
rect 13820 17274 13872 17280
rect 13924 17270 13952 17303
rect 14004 17274 14056 17280
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 14016 17202 14044 17274
rect 14200 17270 14228 17682
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13634 16552 13690 16561
rect 13832 16522 13860 16934
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13634 16487 13690 16496
rect 13820 16516 13872 16522
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 15978 13584 16390
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13358 13832 13414 13841
rect 13358 13767 13414 13776
rect 13372 13734 13400 13767
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 11762 13400 13126
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13556 12102 13584 12854
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13648 11937 13676 16487
rect 13820 16458 13872 16464
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14292 15586 14320 18022
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14200 15558 14320 15586
rect 14200 15434 14228 15558
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14200 14890 14228 15098
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14414 13860 14758
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 13938 13860 14350
rect 14292 14346 14320 14894
rect 14384 14346 14412 17478
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13326 13860 13874
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 14384 13410 14412 14282
rect 14476 13841 14504 18142
rect 14554 18184 14610 18193
rect 14554 18119 14610 18128
rect 14568 15162 14596 18119
rect 14844 15910 14872 18294
rect 15488 17678 15516 18702
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14844 15026 14872 15846
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14936 14822 14964 17546
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15434 15056 15982
rect 15120 15910 15148 16118
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 14958 15056 15370
rect 15120 15094 15148 15846
rect 15212 15178 15240 17002
rect 15488 16998 15516 17274
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15396 15178 15424 16934
rect 15488 16658 15516 16934
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16250 15516 16594
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 16114 15516 16186
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15580 15638 15608 17546
rect 15672 16454 15700 18294
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 15366 15608 15574
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15212 15150 15332 15178
rect 15396 15150 15608 15178
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15304 15042 15332 15150
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14936 14385 14964 14758
rect 14922 14376 14978 14385
rect 14922 14311 14978 14320
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14016 13382 14412 13410
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12986 13860 13262
rect 14016 13258 14044 13382
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14568 13190 14596 14214
rect 15028 14074 15056 14758
rect 15120 14414 15148 15030
rect 15200 15020 15252 15026
rect 15304 15014 15424 15042
rect 15200 14962 15252 14968
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15212 14226 15240 14962
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14346 15332 14826
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15120 14198 15240 14226
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 13634 11928 13690 11937
rect 13452 11892 13504 11898
rect 14200 11898 14228 12174
rect 13634 11863 13690 11872
rect 14188 11892 14240 11898
rect 13452 11834 13504 11840
rect 14188 11834 14240 11840
rect 13464 11762 13492 11834
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 9586 13308 10746
rect 13464 10742 13492 11698
rect 14200 11694 14228 11834
rect 14188 11688 14240 11694
rect 14240 11648 14320 11676
rect 14188 11630 14240 11636
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 7954 12848 8978
rect 13188 8430 13216 9318
rect 13740 8974 13768 11494
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 10810 13860 11154
rect 14188 11144 14240 11150
rect 14292 11132 14320 11648
rect 14240 11104 14320 11132
rect 14188 11086 14240 11092
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 14292 10674 14320 11104
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13832 10266 13860 10610
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14292 10130 14320 10610
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 9586 14320 10066
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 13832 9178 13860 9522
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 14384 8537 14412 12786
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 11354 14504 11698
rect 14752 11558 14780 13942
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12850 14872 13262
rect 14936 12986 14964 13670
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14844 12646 14872 12786
rect 15028 12646 15056 13126
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14844 12238 14872 12582
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 15120 11218 15148 14198
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15212 13462 15240 13738
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15304 12434 15332 13806
rect 15396 13462 15424 15014
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15212 12406 15332 12434
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15212 10577 15240 12406
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 9926 14872 10406
rect 15304 9926 15332 12106
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11354 15516 12038
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15384 10056 15436 10062
rect 15488 10044 15516 11290
rect 15436 10016 15516 10044
rect 15384 9998 15436 10004
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14370 8528 14426 8537
rect 14370 8463 14426 8472
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 15580 6730 15608 15150
rect 15672 13802 15700 16390
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15764 9081 15792 19450
rect 15856 19174 15884 19790
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 9738 15884 19110
rect 16132 18630 16160 19246
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16040 15978 16068 16458
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 12918 15976 15846
rect 16132 15609 16160 18566
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 18154 16252 18226
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16224 17678 16252 18090
rect 17144 18086 17172 18634
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16212 17672 16264 17678
rect 16264 17632 16436 17660
rect 16212 17614 16264 17620
rect 16408 17270 16436 17632
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16408 16998 16436 17206
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16316 16250 16344 16487
rect 16960 16425 16988 16934
rect 16946 16416 17002 16425
rect 16544 16348 16852 16357
rect 16946 16351 17002 16360
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16118 15600 16174 15609
rect 16316 15586 16344 16186
rect 16118 15535 16174 15544
rect 16224 15558 16344 15586
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13394 16068 13670
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15934 11928 15990 11937
rect 15934 11863 15936 11872
rect 15988 11863 15990 11872
rect 15936 11834 15988 11840
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15856 9710 15976 9738
rect 15842 9616 15898 9625
rect 15842 9551 15898 9560
rect 15856 9450 15884 9551
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15750 9072 15806 9081
rect 15750 9007 15806 9016
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15948 6662 15976 9710
rect 16040 9654 16068 9998
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16040 9178 16068 9590
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 16224 5302 16252 15558
rect 16304 15496 16356 15502
rect 16960 15473 16988 16351
rect 16304 15438 16356 15444
rect 16946 15464 17002 15473
rect 16316 15026 16344 15438
rect 16396 15428 16448 15434
rect 16946 15399 17002 15408
rect 16396 15370 16448 15376
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16316 14618 16344 14962
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16408 14074 16436 15370
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 14550 16988 14758
rect 17052 14618 17080 17138
rect 17144 16697 17172 17682
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 17052 14226 17080 14554
rect 16960 14198 17080 14226
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16684 13977 16712 14010
rect 16670 13968 16726 13977
rect 16726 13938 16804 13954
rect 16726 13932 16816 13938
rect 16726 13926 16764 13932
rect 16670 13903 16726 13912
rect 16764 13874 16816 13880
rect 16488 13864 16540 13870
rect 16486 13832 16488 13841
rect 16960 13852 16988 14198
rect 17236 14074 17264 16458
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 16540 13832 16542 13841
rect 16960 13824 17172 13852
rect 16486 13767 16542 13776
rect 16948 13456 17000 13462
rect 16486 13424 16542 13433
rect 16948 13398 17000 13404
rect 16486 13359 16542 13368
rect 16500 13326 16528 13359
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16776 12374 16804 12854
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16316 12238 16344 12310
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 11762 16344 12174
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11830 16436 12038
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16396 11824 16448 11830
rect 16960 11778 16988 13398
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16396 11766 16448 11772
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16868 11750 16988 11778
rect 16316 10674 16344 11698
rect 16868 11082 16896 11750
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 17052 10742 17080 11834
rect 17144 11098 17172 13824
rect 17236 11234 17264 14010
rect 17328 12442 17356 19654
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17420 18290 17448 19450
rect 17604 19174 17632 20334
rect 17696 19242 17724 22200
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17788 20369 17816 20402
rect 17774 20360 17830 20369
rect 17774 20295 17830 20304
rect 17880 19417 17908 20402
rect 18156 20040 18184 22200
rect 18236 20052 18288 20058
rect 18156 20012 18236 20040
rect 18236 19994 18288 20000
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17866 19408 17922 19417
rect 17866 19343 17922 19352
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18340 19334 18368 19722
rect 18616 19514 18644 22200
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18878 19952 18934 19961
rect 18878 19887 18934 19896
rect 18786 19816 18842 19825
rect 18786 19751 18842 19760
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 16182 17448 18226
rect 17498 17640 17554 17649
rect 17498 17575 17554 17584
rect 17512 17542 17540 17575
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17512 16114 17540 16390
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17406 15464 17462 15473
rect 17406 15399 17462 15408
rect 17420 14074 17448 15399
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12918 17448 13330
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17236 11206 17356 11234
rect 17420 11218 17448 11698
rect 17512 11558 17540 15098
rect 17604 13870 17632 19110
rect 17972 18630 18000 19314
rect 18340 19306 18460 19334
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 18064 18306 18092 18702
rect 17972 18278 18092 18306
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17202 17724 17478
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17972 16998 18000 18278
rect 18052 18216 18104 18222
rect 18156 18204 18184 18770
rect 18432 18737 18460 19306
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18104 18176 18184 18204
rect 18052 18158 18104 18164
rect 18064 17882 18092 18158
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18064 17270 18092 17818
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 14521 17816 16050
rect 18156 15366 18184 17138
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18248 16425 18276 16458
rect 18234 16416 18290 16425
rect 18234 16351 18290 16360
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14929 18000 14962
rect 17958 14920 18014 14929
rect 17958 14855 18014 14864
rect 17774 14512 17830 14521
rect 17774 14447 17830 14456
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17696 12889 17724 14282
rect 17682 12880 17738 12889
rect 17682 12815 17738 12824
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17696 11801 17724 11834
rect 17682 11792 17738 11801
rect 17682 11727 17738 11736
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17696 11354 17724 11727
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17144 11082 17264 11098
rect 17144 11076 17276 11082
rect 17144 11070 17224 11076
rect 17224 11018 17276 11024
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 9450 16988 9930
rect 17052 9722 17080 10678
rect 17328 10470 17356 11206
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17144 9654 17172 9998
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 17880 9110 17908 12038
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10062 18092 10406
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9586 18092 9998
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18156 9489 18184 15302
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18248 14618 18276 14962
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18432 10810 18460 18663
rect 18694 17776 18750 17785
rect 18694 17711 18750 17720
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 14074 18552 14214
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18524 13938 18552 14010
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18142 9480 18198 9489
rect 18142 9415 18198 9424
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 18616 6866 18644 15302
rect 18708 9926 18736 17711
rect 18800 13802 18828 19751
rect 18892 19378 18920 19887
rect 18984 19854 19012 20742
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 19076 18970 19104 22200
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19536 18970 19564 22200
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19720 18698 19748 19110
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 18352 19668 18358
rect 19616 18294 19668 18300
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 18170 19472 18226
rect 19444 18142 19564 18170
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19432 17808 19484 17814
rect 19536 17762 19564 18142
rect 19628 17814 19656 18294
rect 19484 17756 19564 17762
rect 19432 17750 19564 17756
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 19444 17734 19564 17750
rect 19720 17746 19748 18634
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16182 19012 16934
rect 19076 16658 19104 17274
rect 19352 17066 19380 17478
rect 19444 17082 19472 17614
rect 19536 17542 19564 17734
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19812 17202 19840 20334
rect 19996 20074 20024 22200
rect 19904 20046 20024 20074
rect 19904 19718 19932 20046
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19996 19446 20024 19858
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19996 18766 20024 19382
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19996 18290 20024 18702
rect 20088 18426 20116 19654
rect 20456 18630 20484 22200
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20640 18290 20668 18566
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 19996 17882 20024 18226
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19996 17338 20024 17818
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19340 17060 19392 17066
rect 19444 17054 19564 17082
rect 19340 17002 19392 17008
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18892 15026 18920 15574
rect 18984 15366 19012 16118
rect 19076 16114 19104 16594
rect 19536 16561 19564 17054
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19720 16590 19748 16934
rect 19708 16584 19760 16590
rect 19522 16552 19578 16561
rect 19708 16526 19760 16532
rect 19522 16487 19578 16496
rect 19904 16114 19932 16934
rect 20088 16794 20116 18226
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20364 16250 20392 17002
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19076 15638 19104 16050
rect 19984 15904 20036 15910
rect 19904 15852 19984 15858
rect 19904 15846 20036 15852
rect 19904 15830 20024 15846
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 13938 18920 14962
rect 19444 14906 19472 15098
rect 19720 15094 19748 15302
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19444 14878 19564 14906
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18892 12986 18920 13874
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18892 12442 18920 12922
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18800 11762 18828 12038
rect 18892 11830 18920 12378
rect 18984 12102 19012 13738
rect 19076 13326 19104 14214
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19536 13530 19564 14878
rect 19720 14618 19748 15030
rect 19904 14822 19932 15830
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 15162 20024 15302
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19904 14414 19932 14758
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12986 19380 13194
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19628 12850 19656 13398
rect 19812 12986 19840 14282
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 19536 11898 19564 12582
rect 19628 12102 19656 12786
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 10266 18828 11698
rect 18892 11218 18920 11766
rect 19628 11665 19656 12038
rect 19614 11656 19670 11665
rect 19614 11591 19670 11600
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 19444 10742 19472 11290
rect 19720 11150 19748 11494
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19628 10742 19656 11086
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19444 10520 19472 10678
rect 19444 10492 19564 10520
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 19338 10160 19394 10169
rect 19338 10095 19394 10104
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18708 9110 18736 9862
rect 19352 9450 19380 10095
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19536 9382 19564 10492
rect 19720 9518 19748 11086
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19904 7818 19932 14350
rect 19996 13258 20024 14758
rect 20364 13938 20392 16186
rect 20732 15706 20760 20402
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20824 17610 20852 19314
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20916 16454 20944 22200
rect 21376 20482 21404 22200
rect 21836 20890 21864 22200
rect 21284 20454 21404 20482
rect 21652 20862 21864 20890
rect 21284 20330 21312 20454
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21376 19922 21404 20334
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21284 18850 21312 19722
rect 21376 19378 21404 19858
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21362 18864 21418 18873
rect 21284 18822 21362 18850
rect 21362 18799 21418 18808
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21008 17610 21036 18362
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 16522 21036 17206
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20824 15434 20852 16390
rect 21100 16153 21128 16526
rect 21086 16144 21142 16153
rect 21086 16079 21142 16088
rect 21086 16008 21142 16017
rect 21086 15943 21088 15952
rect 21140 15943 21142 15952
rect 21088 15914 21140 15920
rect 21100 15586 21128 15914
rect 20916 15558 21128 15586
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20916 14090 20944 15558
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20824 14062 20944 14090
rect 20996 14068 21048 14074
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20088 10810 20116 13194
rect 20364 13190 20392 13874
rect 20824 13258 20852 14062
rect 20996 14010 21048 14016
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20916 13394 20944 13874
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20916 12986 20944 13330
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20548 11830 20576 12038
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20548 9450 20576 11766
rect 21008 11354 21036 14010
rect 21100 14006 21128 15370
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21192 13841 21220 18702
rect 21376 18426 21404 18799
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21652 18358 21680 20862
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 22296 20466 22324 22200
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22756 19174 22784 22200
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21376 17202 21404 17614
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21376 15570 21404 17138
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21376 15026 21404 15506
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21376 14482 21404 14962
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14074 21404 14418
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21178 13832 21234 13841
rect 21178 13767 21234 13776
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21376 12306 21404 12786
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21284 11898 21312 12106
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21376 11762 21404 12242
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21376 11354 21404 11698
rect 21468 11529 21496 13262
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21454 11520 21510 11529
rect 21454 11455 21510 11464
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21086 10704 21142 10713
rect 21376 10674 21404 11290
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21086 10639 21088 10648
rect 21140 10639 21142 10648
rect 21364 10668 21416 10674
rect 21088 10610 21140 10616
rect 21364 10610 21416 10616
rect 21100 10266 21128 10610
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 21100 8634 21128 10202
rect 21376 10062 21404 10610
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21376 9722 21404 9998
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21376 9178 21404 9658
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8634 21404 9114
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 2240 1737 2268 2382
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 2145 2820 2314
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 2778 2136 2834 2145
rect 6148 2139 6456 2148
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 2778 2071 2834 2080
rect 2226 1728 2282 1737
rect 2226 1663 2282 1672
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 2246
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 11532 734 11744 762
<< via2 >>
rect 1490 18808 1546 18864
rect 2042 21256 2098 21312
rect 1490 18400 1546 18456
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15544 1546 15600
rect 1490 15136 1546 15192
rect 2134 19236 2190 19272
rect 2134 19216 2136 19236
rect 2136 19216 2188 19236
rect 2188 19216 2190 19236
rect 2778 20032 2834 20088
rect 2134 17584 2190 17640
rect 2778 19660 2780 19680
rect 2780 19660 2832 19680
rect 2832 19660 2834 19680
rect 2778 19624 2834 19660
rect 2042 15972 2098 16008
rect 2042 15952 2044 15972
rect 2044 15952 2096 15972
rect 2096 15952 2098 15972
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1490 13912 1546 13968
rect 1490 13504 1546 13560
rect 1398 13096 1454 13152
rect 1398 12708 1454 12744
rect 1398 12688 1400 12708
rect 1400 12688 1452 12708
rect 1452 12688 1454 12708
rect 1398 11872 1454 11928
rect 1398 11464 1454 11520
rect 1490 11056 1546 11112
rect 1398 10240 1454 10296
rect 1398 9832 1454 9888
rect 1398 9424 1454 9480
rect 1674 10784 1730 10840
rect 2042 14320 2098 14376
rect 2042 12280 2098 12336
rect 1950 12144 2006 12200
rect 1398 8744 1454 8800
rect 1858 8608 1914 8664
rect 1398 8200 1454 8256
rect 2134 9968 2190 10024
rect 3146 20440 3202 20496
rect 3974 20848 4030 20904
rect 2318 12280 2374 12336
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3422 19488 3478 19544
rect 3514 19216 3570 19272
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 4066 19760 4122 19816
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3790 17176 3846 17232
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3514 15000 3570 15056
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 4158 15428 4214 15464
rect 4158 15408 4160 15428
rect 4160 15408 4212 15428
rect 4212 15408 4214 15428
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3974 11736 4030 11792
rect 3606 11636 3608 11656
rect 3608 11636 3660 11656
rect 3660 11636 3662 11656
rect 3606 11600 3662 11636
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 4434 16088 4490 16144
rect 4434 14900 4436 14920
rect 4436 14900 4488 14920
rect 4488 14900 4490 14920
rect 4434 14864 4490 14900
rect 4802 16496 4858 16552
rect 5538 19352 5594 19408
rect 5170 17076 5172 17096
rect 5172 17076 5224 17096
rect 5224 17076 5226 17096
rect 5170 17040 5226 17076
rect 4894 15816 4950 15872
rect 4894 15408 4950 15464
rect 4618 13404 4620 13424
rect 4620 13404 4672 13424
rect 4672 13404 4674 13424
rect 4618 13368 4674 13404
rect 2778 10648 2834 10704
rect 2686 10548 2688 10568
rect 2688 10548 2740 10568
rect 2740 10548 2742 10568
rect 2686 10512 2742 10548
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6642 20440 6698 20496
rect 6550 19780 6606 19816
rect 6550 19760 6552 19780
rect 6552 19760 6604 19780
rect 6604 19760 6606 19780
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5998 19352 6054 19408
rect 6366 19388 6368 19408
rect 6368 19388 6420 19408
rect 6420 19388 6422 19408
rect 6366 19352 6422 19388
rect 6550 19352 6606 19408
rect 6458 18808 6514 18864
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5354 14864 5410 14920
rect 5262 12960 5318 13016
rect 5170 12824 5226 12880
rect 1858 7828 1860 7848
rect 1860 7828 1912 7848
rect 1912 7828 1914 7848
rect 1858 7792 1914 7828
rect 2778 9016 2834 9072
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 1398 7404 1454 7440
rect 1398 7384 1400 7404
rect 1400 7384 1452 7404
rect 1452 7384 1454 7404
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 1858 6976 1914 7032
rect 1398 6568 1454 6624
rect 1398 6160 1454 6216
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 1858 5752 1914 5808
rect 1398 5344 1454 5400
rect 2226 4936 2282 4992
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 2226 4564 2228 4584
rect 2228 4564 2280 4584
rect 2280 4564 2282 4584
rect 2226 4528 2282 4564
rect 1490 4140 1546 4176
rect 1490 4120 1492 4140
rect 1492 4120 1544 4140
rect 1544 4120 1546 4140
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 2042 3712 2098 3768
rect 5630 12416 5686 12472
rect 5354 11056 5410 11112
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 5814 13912 5870 13968
rect 6918 18828 6974 18864
rect 6918 18808 6920 18828
rect 6920 18808 6972 18828
rect 6972 18808 6974 18828
rect 6826 17740 6882 17776
rect 6826 17720 6828 17740
rect 6828 17720 6880 17740
rect 6880 17720 6882 17740
rect 7010 17992 7066 18048
rect 7194 17176 7250 17232
rect 6550 14184 6606 14240
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 7010 15988 7012 16008
rect 7012 15988 7064 16008
rect 7064 15988 7066 16008
rect 7010 15952 7066 15988
rect 6826 14612 6882 14648
rect 6826 14592 6828 14612
rect 6828 14592 6880 14612
rect 6880 14592 6882 14612
rect 6642 13232 6698 13288
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6642 12416 6698 12472
rect 5722 12144 5778 12200
rect 5262 10124 5318 10160
rect 5262 10104 5264 10124
rect 5264 10104 5316 10124
rect 5316 10104 5318 10124
rect 1490 3304 1546 3360
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6642 11872 6698 11928
rect 6182 11212 6238 11248
rect 6182 11192 6184 11212
rect 6184 11192 6236 11212
rect 6236 11192 6238 11212
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 7194 15564 7250 15600
rect 7194 15544 7196 15564
rect 7196 15544 7248 15564
rect 7248 15544 7250 15564
rect 7470 18164 7472 18184
rect 7472 18164 7524 18184
rect 7524 18164 7526 18184
rect 7470 18128 7526 18164
rect 7102 12180 7104 12200
rect 7104 12180 7156 12200
rect 7156 12180 7158 12200
rect 7102 12144 7158 12180
rect 7470 16088 7526 16144
rect 7838 16652 7894 16688
rect 7838 16632 7840 16652
rect 7840 16632 7892 16652
rect 7892 16632 7894 16652
rect 8206 17584 8262 17640
rect 7838 16088 7894 16144
rect 7838 15816 7894 15872
rect 7654 15020 7710 15056
rect 7654 15000 7656 15020
rect 7656 15000 7708 15020
rect 7708 15000 7710 15020
rect 7562 14864 7618 14920
rect 7746 14864 7802 14920
rect 7286 10240 7342 10296
rect 7102 9968 7158 10024
rect 6550 8472 6606 8528
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6826 8880 6882 8936
rect 5906 6740 5908 6760
rect 5908 6740 5960 6760
rect 5960 6740 5962 6760
rect 5906 6704 5962 6740
rect 7838 14728 7894 14784
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 1490 2896 1546 2952
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 2042 2488 2098 2544
rect 7746 7948 7802 7984
rect 7746 7928 7748 7948
rect 7748 7928 7800 7948
rect 7800 7928 7802 7948
rect 8482 19488 8538 19544
rect 8298 14728 8354 14784
rect 8206 14320 8262 14376
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8574 18264 8630 18320
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 9402 19508 9458 19544
rect 9402 19488 9404 19508
rect 9404 19488 9456 19508
rect 9456 19488 9458 19508
rect 9034 17040 9090 17096
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9402 18400 9458 18456
rect 9862 20304 9918 20360
rect 9770 20032 9826 20088
rect 9678 19932 9680 19952
rect 9680 19932 9732 19952
rect 9732 19932 9734 19952
rect 9678 19896 9734 19932
rect 9678 19760 9734 19816
rect 9126 13912 9182 13968
rect 9126 13776 9182 13832
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9034 9460 9036 9480
rect 9036 9460 9088 9480
rect 9088 9460 9090 9480
rect 9034 9424 9090 9460
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9402 12144 9458 12200
rect 9862 13912 9918 13968
rect 10046 18164 10048 18184
rect 10048 18164 10100 18184
rect 10100 18164 10102 18184
rect 10046 18128 10102 18164
rect 10414 19216 10470 19272
rect 10598 19080 10654 19136
rect 10598 18672 10654 18728
rect 10138 14456 10194 14512
rect 10046 11872 10102 11928
rect 10414 13252 10470 13288
rect 10414 13232 10416 13252
rect 10416 13232 10468 13252
rect 10468 13232 10470 13252
rect 10966 19352 11022 19408
rect 10966 17856 11022 17912
rect 10966 17312 11022 17368
rect 10966 14184 11022 14240
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11150 18400 11206 18456
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11978 18672 12034 18728
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11978 17856 12034 17912
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11702 15952 11758 16008
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10874 8628 10930 8664
rect 10874 8608 10876 8628
rect 10876 8608 10928 8628
rect 10928 8608 10930 8628
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 10966 8472 11022 8528
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11518 12280 11574 12336
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11978 16632 12034 16688
rect 12162 16668 12164 16688
rect 12164 16668 12216 16688
rect 12216 16668 12218 16688
rect 12162 16632 12218 16668
rect 11794 11056 11850 11112
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 12622 17312 12678 17368
rect 12898 20052 12954 20088
rect 12898 20032 12900 20052
rect 12900 20032 12952 20052
rect 12952 20032 12954 20052
rect 12898 19760 12954 19816
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13266 19624 13322 19680
rect 13542 19080 13598 19136
rect 12990 16108 13046 16144
rect 12990 16088 12992 16108
rect 12992 16088 13044 16108
rect 13044 16088 13046 16108
rect 13726 18264 13782 18320
rect 15198 20460 15254 20496
rect 15198 20440 15200 20460
rect 15200 20440 15252 20460
rect 15252 20440 15254 20460
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13910 17312 13966 17368
rect 13634 16496 13690 16552
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13358 13776 13414 13832
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 14554 18128 14610 18184
rect 14922 14320 14978 14376
rect 14462 13776 14518 13832
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13634 11872 13690 11928
rect 13266 11192 13322 11248
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 15198 10512 15254 10568
rect 14370 8472 14426 8528
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16302 16496 16358 16552
rect 16946 16360 17002 16416
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16118 15544 16174 15600
rect 15934 11892 15990 11928
rect 15934 11872 15936 11892
rect 15936 11872 15988 11892
rect 15988 11872 15990 11892
rect 15842 9560 15898 9616
rect 15750 9016 15806 9072
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 16946 15408 17002 15464
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 17130 16632 17186 16688
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16670 13912 16726 13968
rect 16486 13812 16488 13832
rect 16488 13812 16540 13832
rect 16540 13812 16542 13832
rect 16486 13776 16542 13812
rect 16486 13368 16542 13424
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 17774 20304 17830 20360
rect 17866 19352 17922 19408
rect 18878 19896 18934 19952
rect 18786 19760 18842 19816
rect 17498 17584 17554 17640
rect 17406 15408 17462 15464
rect 18418 18672 18474 18728
rect 18234 16360 18290 16416
rect 17958 14864 18014 14920
rect 17774 14456 17830 14512
rect 17682 12824 17738 12880
rect 17682 11736 17738 11792
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 18694 17720 18750 17776
rect 18142 9424 18198 9480
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19522 16496 19578 16552
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19614 11600 19670 11656
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19338 10104 19394 10160
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 21362 18808 21418 18864
rect 21086 16088 21142 16144
rect 21086 15972 21142 16008
rect 21086 15952 21088 15972
rect 21088 15952 21140 15972
rect 21140 15952 21142 15972
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21178 13776 21234 13832
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21454 11464 21510 11520
rect 21086 10668 21142 10704
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21086 10648 21088 10668
rect 21088 10648 21140 10668
rect 21140 10648 21142 10668
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 2778 2080 2834 2136
rect 2226 1672 2282 1728
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 2037 21314 2103 21317
rect 0 21312 2103 21314
rect 0 21256 2042 21312
rect 2098 21256 2103 21312
rect 0 21254 2103 21256
rect 0 21224 800 21254
rect 2037 21251 2103 21254
rect 0 20906 800 20936
rect 3969 20906 4035 20909
rect 0 20904 4035 20906
rect 0 20848 3974 20904
rect 4030 20848 4035 20904
rect 0 20846 4035 20848
rect 0 20816 800 20846
rect 3969 20843 4035 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 3141 20498 3207 20501
rect 0 20496 3207 20498
rect 0 20440 3146 20496
rect 3202 20440 3207 20496
rect 0 20438 3207 20440
rect 0 20408 800 20438
rect 3141 20435 3207 20438
rect 6637 20498 6703 20501
rect 15193 20498 15259 20501
rect 6637 20496 15259 20498
rect 6637 20440 6642 20496
rect 6698 20440 15198 20496
rect 15254 20440 15259 20496
rect 6637 20438 15259 20440
rect 6637 20435 6703 20438
rect 15193 20435 15259 20438
rect 9857 20362 9923 20365
rect 17769 20362 17835 20365
rect 9857 20360 17835 20362
rect 9857 20304 9862 20360
rect 9918 20304 17774 20360
rect 17830 20304 17835 20360
rect 9857 20302 17835 20304
rect 9857 20299 9923 20302
rect 17769 20299 17835 20302
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 2773 20090 2839 20093
rect 0 20088 2839 20090
rect 0 20032 2778 20088
rect 2834 20032 2839 20088
rect 0 20030 2839 20032
rect 0 20000 800 20030
rect 2773 20027 2839 20030
rect 9765 20090 9831 20093
rect 12893 20090 12959 20093
rect 9765 20088 12959 20090
rect 9765 20032 9770 20088
rect 9826 20032 12898 20088
rect 12954 20032 12959 20088
rect 9765 20030 12959 20032
rect 9765 20027 9831 20030
rect 12893 20027 12959 20030
rect 9673 19954 9739 19957
rect 18873 19954 18939 19957
rect 9673 19952 18939 19954
rect 9673 19896 9678 19952
rect 9734 19896 18878 19952
rect 18934 19896 18939 19952
rect 9673 19894 18939 19896
rect 9673 19891 9739 19894
rect 18873 19891 18939 19894
rect 4061 19818 4127 19821
rect 6545 19818 6611 19821
rect 4061 19816 6611 19818
rect 4061 19760 4066 19816
rect 4122 19760 6550 19816
rect 6606 19760 6611 19816
rect 4061 19758 6611 19760
rect 4061 19755 4127 19758
rect 6545 19755 6611 19758
rect 9673 19818 9739 19821
rect 12893 19818 12959 19821
rect 18781 19818 18847 19821
rect 9673 19816 12450 19818
rect 9673 19760 9678 19816
rect 9734 19760 12450 19816
rect 9673 19758 12450 19760
rect 9673 19755 9739 19758
rect 0 19682 800 19712
rect 2773 19682 2839 19685
rect 0 19680 2839 19682
rect 0 19624 2778 19680
rect 2834 19624 2839 19680
rect 0 19622 2839 19624
rect 12390 19682 12450 19758
rect 12893 19816 18847 19818
rect 12893 19760 12898 19816
rect 12954 19760 18786 19816
rect 18842 19760 18847 19816
rect 12893 19758 18847 19760
rect 12893 19755 12959 19758
rect 18781 19755 18847 19758
rect 13261 19682 13327 19685
rect 12390 19680 13327 19682
rect 12390 19624 13266 19680
rect 13322 19624 13327 19680
rect 12390 19622 13327 19624
rect 0 19592 800 19622
rect 2773 19619 2839 19622
rect 13261 19619 13327 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 3417 19546 3483 19549
rect 8477 19548 8543 19549
rect 3918 19546 3924 19548
rect 3417 19544 3924 19546
rect 3417 19488 3422 19544
rect 3478 19488 3924 19544
rect 3417 19486 3924 19488
rect 3417 19483 3483 19486
rect 3918 19484 3924 19486
rect 3988 19484 3994 19548
rect 8477 19544 8524 19548
rect 8588 19546 8594 19548
rect 9397 19546 9463 19549
rect 8477 19488 8482 19544
rect 8477 19484 8524 19488
rect 8588 19486 8634 19546
rect 9397 19544 11162 19546
rect 9397 19488 9402 19544
rect 9458 19488 11162 19544
rect 9397 19486 11162 19488
rect 8588 19484 8594 19486
rect 8477 19483 8543 19484
rect 9397 19483 9463 19486
rect 5533 19412 5599 19413
rect 5993 19412 6059 19413
rect 5533 19408 5580 19412
rect 5644 19410 5650 19412
rect 5942 19410 5948 19412
rect 5533 19352 5538 19408
rect 5533 19348 5580 19352
rect 5644 19350 5690 19410
rect 5902 19350 5948 19410
rect 6012 19408 6059 19412
rect 6054 19352 6059 19408
rect 5644 19348 5650 19350
rect 5942 19348 5948 19350
rect 6012 19348 6059 19352
rect 5533 19347 5599 19348
rect 5993 19347 6059 19348
rect 6361 19410 6427 19413
rect 6545 19410 6611 19413
rect 10961 19412 11027 19413
rect 10910 19410 10916 19412
rect 6361 19408 6611 19410
rect 6361 19352 6366 19408
rect 6422 19352 6550 19408
rect 6606 19352 6611 19408
rect 6361 19350 6611 19352
rect 10870 19350 10916 19410
rect 10980 19408 11027 19412
rect 11022 19352 11027 19408
rect 6361 19347 6427 19350
rect 6545 19347 6611 19350
rect 10910 19348 10916 19350
rect 10980 19348 11027 19352
rect 11102 19410 11162 19486
rect 17861 19410 17927 19413
rect 11102 19408 17927 19410
rect 11102 19352 17866 19408
rect 17922 19352 17927 19408
rect 11102 19350 17927 19352
rect 10961 19347 11027 19348
rect 17861 19347 17927 19350
rect 0 19274 800 19304
rect 2129 19274 2195 19277
rect 0 19272 2195 19274
rect 0 19216 2134 19272
rect 2190 19216 2195 19272
rect 0 19214 2195 19216
rect 0 19184 800 19214
rect 2129 19211 2195 19214
rect 3509 19274 3575 19277
rect 10409 19274 10475 19277
rect 3509 19272 10475 19274
rect 3509 19216 3514 19272
rect 3570 19216 10414 19272
rect 10470 19216 10475 19272
rect 3509 19214 10475 19216
rect 3509 19211 3575 19214
rect 10409 19211 10475 19214
rect 10593 19138 10659 19141
rect 13537 19138 13603 19141
rect 10593 19136 13603 19138
rect 10593 19080 10598 19136
rect 10654 19080 13542 19136
rect 13598 19080 13603 19136
rect 10593 19078 13603 19080
rect 10593 19075 10659 19078
rect 13537 19075 13603 19078
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 6453 18866 6519 18869
rect 6678 18866 6684 18868
rect 6453 18864 6684 18866
rect 6453 18808 6458 18864
rect 6514 18808 6684 18864
rect 6453 18806 6684 18808
rect 6453 18803 6519 18806
rect 6678 18804 6684 18806
rect 6748 18804 6754 18868
rect 6913 18866 6979 18869
rect 21357 18866 21423 18869
rect 6913 18864 21423 18866
rect 6913 18808 6918 18864
rect 6974 18808 21362 18864
rect 21418 18808 21423 18864
rect 6913 18806 21423 18808
rect 6913 18803 6979 18806
rect 21357 18803 21423 18806
rect 5390 18668 5396 18732
rect 5460 18730 5466 18732
rect 10593 18730 10659 18733
rect 5460 18728 10659 18730
rect 5460 18672 10598 18728
rect 10654 18672 10659 18728
rect 5460 18670 10659 18672
rect 5460 18668 5466 18670
rect 10593 18667 10659 18670
rect 11973 18730 12039 18733
rect 18413 18730 18479 18733
rect 11973 18728 18479 18730
rect 11973 18672 11978 18728
rect 12034 18672 18418 18728
rect 18474 18672 18479 18728
rect 11973 18670 18479 18672
rect 11973 18667 12039 18670
rect 18413 18667 18479 18670
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 9397 18458 9463 18461
rect 11145 18458 11211 18461
rect 9397 18456 11211 18458
rect 9397 18400 9402 18456
rect 9458 18400 11150 18456
rect 11206 18400 11211 18456
rect 9397 18398 11211 18400
rect 9397 18395 9463 18398
rect 11145 18395 11211 18398
rect 8569 18322 8635 18325
rect 13721 18322 13787 18325
rect 8569 18320 13787 18322
rect 8569 18264 8574 18320
rect 8630 18264 13726 18320
rect 13782 18264 13787 18320
rect 8569 18262 13787 18264
rect 8569 18259 8635 18262
rect 13721 18259 13787 18262
rect 7465 18186 7531 18189
rect 10041 18186 10107 18189
rect 14549 18186 14615 18189
rect 7465 18184 14615 18186
rect 7465 18128 7470 18184
rect 7526 18128 10046 18184
rect 10102 18128 14554 18184
rect 14610 18128 14615 18184
rect 7465 18126 14615 18128
rect 7465 18123 7531 18126
rect 10041 18123 10107 18126
rect 14549 18123 14615 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 7005 18052 7071 18053
rect 7005 18048 7052 18052
rect 7116 18050 7122 18052
rect 7005 17992 7010 18048
rect 7005 17988 7052 17992
rect 7116 17990 7162 18050
rect 7116 17988 7122 17990
rect 7005 17987 7071 17988
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 10961 17914 11027 17917
rect 11973 17914 12039 17917
rect 10961 17912 12039 17914
rect 10961 17856 10966 17912
rect 11022 17856 11978 17912
rect 12034 17856 12039 17912
rect 10961 17854 12039 17856
rect 10961 17851 11027 17854
rect 11973 17851 12039 17854
rect 6821 17778 6887 17781
rect 18689 17778 18755 17781
rect 6821 17776 18755 17778
rect 6821 17720 6826 17776
rect 6882 17720 18694 17776
rect 18750 17720 18755 17776
rect 6821 17718 18755 17720
rect 6821 17715 6887 17718
rect 18689 17715 18755 17718
rect 0 17642 800 17672
rect 2129 17642 2195 17645
rect 0 17640 2195 17642
rect 0 17584 2134 17640
rect 2190 17584 2195 17640
rect 0 17582 2195 17584
rect 0 17552 800 17582
rect 2129 17579 2195 17582
rect 8201 17642 8267 17645
rect 17493 17642 17559 17645
rect 8201 17640 17559 17642
rect 8201 17584 8206 17640
rect 8262 17584 17498 17640
rect 17554 17584 17559 17640
rect 8201 17582 17559 17584
rect 8201 17579 8267 17582
rect 17493 17579 17559 17582
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 10961 17370 11027 17373
rect 7054 17368 11027 17370
rect 7054 17312 10966 17368
rect 11022 17312 11027 17368
rect 7054 17310 11027 17312
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 3785 17234 3851 17237
rect 7054 17234 7114 17310
rect 10961 17307 11027 17310
rect 12617 17370 12683 17373
rect 13905 17370 13971 17373
rect 12617 17368 13971 17370
rect 12617 17312 12622 17368
rect 12678 17312 13910 17368
rect 13966 17312 13971 17368
rect 12617 17310 13971 17312
rect 12617 17307 12683 17310
rect 13905 17307 13971 17310
rect 3785 17232 7114 17234
rect 3785 17176 3790 17232
rect 3846 17176 7114 17232
rect 3785 17174 7114 17176
rect 7189 17234 7255 17237
rect 13118 17234 13124 17236
rect 7189 17232 13124 17234
rect 7189 17176 7194 17232
rect 7250 17176 13124 17232
rect 7189 17174 13124 17176
rect 3785 17171 3851 17174
rect 7189 17171 7255 17174
rect 13118 17172 13124 17174
rect 13188 17172 13194 17236
rect 5165 17098 5231 17101
rect 6862 17098 6868 17100
rect 5165 17096 6868 17098
rect 5165 17040 5170 17096
rect 5226 17040 6868 17096
rect 5165 17038 6868 17040
rect 5165 17035 5231 17038
rect 6862 17036 6868 17038
rect 6932 17036 6938 17100
rect 8334 17036 8340 17100
rect 8404 17098 8410 17100
rect 9029 17098 9095 17101
rect 8404 17096 9095 17098
rect 8404 17040 9034 17096
rect 9090 17040 9095 17096
rect 8404 17038 9095 17040
rect 8404 17036 8410 17038
rect 9029 17035 9095 17038
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 7833 16690 7899 16693
rect 11973 16690 12039 16693
rect 7833 16688 12039 16690
rect 7833 16632 7838 16688
rect 7894 16632 11978 16688
rect 12034 16632 12039 16688
rect 7833 16630 12039 16632
rect 7833 16627 7899 16630
rect 11973 16627 12039 16630
rect 12157 16690 12223 16693
rect 17125 16690 17191 16693
rect 12157 16688 17191 16690
rect 12157 16632 12162 16688
rect 12218 16632 17130 16688
rect 17186 16632 17191 16688
rect 12157 16630 17191 16632
rect 12157 16627 12223 16630
rect 17125 16627 17191 16630
rect 4797 16554 4863 16557
rect 13629 16554 13695 16557
rect 4797 16552 13695 16554
rect 4797 16496 4802 16552
rect 4858 16496 13634 16552
rect 13690 16496 13695 16552
rect 4797 16494 13695 16496
rect 4797 16491 4863 16494
rect 13629 16491 13695 16494
rect 16297 16554 16363 16557
rect 19517 16554 19583 16557
rect 16297 16552 19583 16554
rect 16297 16496 16302 16552
rect 16358 16496 19522 16552
rect 19578 16496 19583 16552
rect 16297 16494 19583 16496
rect 16297 16491 16363 16494
rect 19517 16491 19583 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 16941 16418 17007 16421
rect 18229 16418 18295 16421
rect 16941 16416 18295 16418
rect 16941 16360 16946 16416
rect 17002 16360 18234 16416
rect 18290 16360 18295 16416
rect 16941 16358 18295 16360
rect 16941 16355 17007 16358
rect 18229 16355 18295 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 4429 16146 4495 16149
rect 7465 16146 7531 16149
rect 4429 16144 7531 16146
rect 4429 16088 4434 16144
rect 4490 16088 7470 16144
rect 7526 16088 7531 16144
rect 4429 16086 7531 16088
rect 4429 16083 4495 16086
rect 7465 16083 7531 16086
rect 7833 16146 7899 16149
rect 12985 16148 13051 16149
rect 12934 16146 12940 16148
rect 7833 16144 12450 16146
rect 7833 16088 7838 16144
rect 7894 16088 12450 16144
rect 7833 16086 12450 16088
rect 12858 16086 12940 16146
rect 13004 16146 13051 16148
rect 21081 16146 21147 16149
rect 13004 16144 21147 16146
rect 13046 16088 21086 16144
rect 21142 16088 21147 16144
rect 7833 16083 7899 16086
rect 0 16010 800 16040
rect 2037 16010 2103 16013
rect 0 16008 2103 16010
rect 0 15952 2042 16008
rect 2098 15952 2103 16008
rect 0 15950 2103 15952
rect 0 15920 800 15950
rect 2037 15947 2103 15950
rect 7005 16010 7071 16013
rect 11697 16010 11763 16013
rect 7005 16008 11763 16010
rect 7005 15952 7010 16008
rect 7066 15952 11702 16008
rect 11758 15952 11763 16008
rect 7005 15950 11763 15952
rect 12390 16010 12450 16086
rect 12934 16084 12940 16086
rect 13004 16086 21147 16088
rect 13004 16084 13051 16086
rect 12985 16083 13051 16084
rect 21081 16083 21147 16086
rect 21081 16010 21147 16013
rect 12390 16008 21147 16010
rect 12390 15952 21086 16008
rect 21142 15952 21147 16008
rect 12390 15950 21147 15952
rect 7005 15947 7071 15950
rect 11697 15947 11763 15950
rect 21081 15947 21147 15950
rect 4889 15874 4955 15877
rect 7833 15874 7899 15877
rect 4889 15872 7899 15874
rect 4889 15816 4894 15872
rect 4950 15816 7838 15872
rect 7894 15816 7899 15872
rect 4889 15814 7899 15816
rect 4889 15811 4955 15814
rect 7833 15811 7899 15814
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 7189 15602 7255 15605
rect 16113 15602 16179 15605
rect 7189 15600 16179 15602
rect 7189 15544 7194 15600
rect 7250 15544 16118 15600
rect 16174 15544 16179 15600
rect 7189 15542 16179 15544
rect 7189 15539 7255 15542
rect 16113 15539 16179 15542
rect 4153 15466 4219 15469
rect 4889 15466 4955 15469
rect 16941 15466 17007 15469
rect 17401 15466 17467 15469
rect 4153 15464 17467 15466
rect 4153 15408 4158 15464
rect 4214 15408 4894 15464
rect 4950 15408 16946 15464
rect 17002 15408 17406 15464
rect 17462 15408 17467 15464
rect 4153 15406 17467 15408
rect 4153 15403 4219 15406
rect 4889 15403 4955 15406
rect 16941 15403 17007 15406
rect 17401 15403 17467 15406
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 3509 15058 3575 15061
rect 7649 15058 7715 15061
rect 3509 15056 7715 15058
rect 3509 15000 3514 15056
rect 3570 15000 7654 15056
rect 7710 15000 7715 15056
rect 3509 14998 7715 15000
rect 3509 14995 3575 14998
rect 7649 14995 7715 14998
rect 4429 14922 4495 14925
rect 5349 14922 5415 14925
rect 7557 14922 7623 14925
rect 4429 14920 7623 14922
rect 4429 14864 4434 14920
rect 4490 14864 5354 14920
rect 5410 14864 7562 14920
rect 7618 14864 7623 14920
rect 4429 14862 7623 14864
rect 4429 14859 4495 14862
rect 5349 14859 5415 14862
rect 7557 14859 7623 14862
rect 7741 14922 7807 14925
rect 17953 14922 18019 14925
rect 7741 14920 18019 14922
rect 7741 14864 7746 14920
rect 7802 14864 17958 14920
rect 18014 14864 18019 14920
rect 7741 14862 18019 14864
rect 7741 14859 7807 14862
rect 17953 14859 18019 14862
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 7833 14786 7899 14789
rect 8293 14786 8359 14789
rect 7833 14784 8359 14786
rect 7833 14728 7838 14784
rect 7894 14728 8298 14784
rect 8354 14728 8359 14784
rect 7833 14726 8359 14728
rect 7833 14723 7899 14726
rect 8293 14723 8359 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 6678 14588 6684 14652
rect 6748 14650 6754 14652
rect 6821 14650 6887 14653
rect 6748 14648 6887 14650
rect 6748 14592 6826 14648
rect 6882 14592 6887 14648
rect 6748 14590 6887 14592
rect 6748 14588 6754 14590
rect 6821 14587 6887 14590
rect 10133 14514 10199 14517
rect 17769 14514 17835 14517
rect 10133 14512 17835 14514
rect 10133 14456 10138 14512
rect 10194 14456 17774 14512
rect 17830 14456 17835 14512
rect 10133 14454 17835 14456
rect 10133 14451 10199 14454
rect 17769 14451 17835 14454
rect 0 14378 800 14408
rect 2037 14378 2103 14381
rect 0 14376 2103 14378
rect 0 14320 2042 14376
rect 2098 14320 2103 14376
rect 0 14318 2103 14320
rect 0 14288 800 14318
rect 2037 14315 2103 14318
rect 8201 14378 8267 14381
rect 14917 14378 14983 14381
rect 8201 14376 14983 14378
rect 8201 14320 8206 14376
rect 8262 14320 14922 14376
rect 14978 14320 14983 14376
rect 8201 14318 14983 14320
rect 8201 14315 8267 14318
rect 14917 14315 14983 14318
rect 6545 14242 6611 14245
rect 10961 14242 11027 14245
rect 6545 14240 11027 14242
rect 6545 14184 6550 14240
rect 6606 14184 10966 14240
rect 11022 14184 11027 14240
rect 6545 14182 11027 14184
rect 6545 14179 6611 14182
rect 10961 14179 11027 14182
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 2078 13908 2084 13972
rect 2148 13970 2154 13972
rect 5809 13970 5875 13973
rect 9121 13970 9187 13973
rect 2148 13910 2790 13970
rect 2148 13908 2154 13910
rect 2730 13834 2790 13910
rect 5809 13968 9187 13970
rect 5809 13912 5814 13968
rect 5870 13912 9126 13968
rect 9182 13912 9187 13968
rect 5809 13910 9187 13912
rect 5809 13907 5875 13910
rect 9121 13907 9187 13910
rect 9857 13970 9923 13973
rect 16665 13970 16731 13973
rect 9857 13968 16731 13970
rect 9857 13912 9862 13968
rect 9918 13912 16670 13968
rect 16726 13912 16731 13968
rect 9857 13910 16731 13912
rect 9857 13907 9923 13910
rect 16665 13907 16731 13910
rect 8334 13834 8340 13836
rect 2730 13774 8340 13834
rect 8334 13772 8340 13774
rect 8404 13772 8410 13836
rect 8518 13772 8524 13836
rect 8588 13834 8594 13836
rect 9121 13834 9187 13837
rect 8588 13832 9187 13834
rect 8588 13776 9126 13832
rect 9182 13776 9187 13832
rect 8588 13774 9187 13776
rect 8588 13772 8594 13774
rect 9121 13771 9187 13774
rect 13353 13834 13419 13837
rect 14457 13834 14523 13837
rect 13353 13832 14523 13834
rect 13353 13776 13358 13832
rect 13414 13776 14462 13832
rect 14518 13776 14523 13832
rect 13353 13774 14523 13776
rect 13353 13771 13419 13774
rect 14457 13771 14523 13774
rect 16481 13834 16547 13837
rect 21173 13834 21239 13837
rect 16481 13832 21239 13834
rect 16481 13776 16486 13832
rect 16542 13776 21178 13832
rect 21234 13776 21239 13832
rect 16481 13774 21239 13776
rect 16481 13771 16547 13774
rect 21173 13771 21239 13774
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 4613 13426 4679 13429
rect 16481 13426 16547 13429
rect 4613 13424 16547 13426
rect 4613 13368 4618 13424
rect 4674 13368 16486 13424
rect 16542 13368 16547 13424
rect 4613 13366 16547 13368
rect 4613 13363 4679 13366
rect 16481 13363 16547 13366
rect 6637 13290 6703 13293
rect 10409 13290 10475 13293
rect 6637 13288 10475 13290
rect 6637 13232 6642 13288
rect 6698 13232 10414 13288
rect 10470 13232 10475 13288
rect 6637 13230 10475 13232
rect 6637 13227 6703 13230
rect 10409 13227 10475 13230
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 5257 13018 5323 13021
rect 5390 13018 5396 13020
rect 5257 13016 5396 13018
rect 5257 12960 5262 13016
rect 5318 12960 5396 13016
rect 5257 12958 5396 12960
rect 5257 12955 5323 12958
rect 5390 12956 5396 12958
rect 5460 12956 5466 13020
rect 5165 12882 5231 12885
rect 17677 12882 17743 12885
rect 5165 12880 17743 12882
rect 5165 12824 5170 12880
rect 5226 12824 17682 12880
rect 17738 12824 17743 12880
rect 5165 12822 17743 12824
rect 5165 12819 5231 12822
rect 17677 12819 17743 12822
rect 0 12746 800 12776
rect 1393 12746 1459 12749
rect 0 12744 1459 12746
rect 0 12688 1398 12744
rect 1454 12688 1459 12744
rect 0 12686 1459 12688
rect 0 12656 800 12686
rect 1393 12683 1459 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 5625 12474 5691 12477
rect 6637 12474 6703 12477
rect 5625 12472 6703 12474
rect 5625 12416 5630 12472
rect 5686 12416 6642 12472
rect 6698 12416 6703 12472
rect 5625 12414 6703 12416
rect 5625 12411 5691 12414
rect 6637 12411 6703 12414
rect 0 12338 800 12368
rect 2037 12338 2103 12341
rect 0 12336 2103 12338
rect 0 12280 2042 12336
rect 2098 12280 2103 12336
rect 0 12278 2103 12280
rect 0 12248 800 12278
rect 2037 12275 2103 12278
rect 2313 12338 2379 12341
rect 11513 12338 11579 12341
rect 2313 12336 11579 12338
rect 2313 12280 2318 12336
rect 2374 12280 11518 12336
rect 11574 12280 11579 12336
rect 2313 12278 11579 12280
rect 2313 12275 2379 12278
rect 11513 12275 11579 12278
rect 1945 12202 2011 12205
rect 2078 12202 2084 12204
rect 1945 12200 2084 12202
rect 1945 12144 1950 12200
rect 2006 12144 2084 12200
rect 1945 12142 2084 12144
rect 1945 12139 2011 12142
rect 2078 12140 2084 12142
rect 2148 12140 2154 12204
rect 5717 12202 5783 12205
rect 7097 12202 7163 12205
rect 9397 12202 9463 12205
rect 5717 12200 6700 12202
rect 5717 12144 5722 12200
rect 5778 12144 6700 12200
rect 5717 12142 6700 12144
rect 5717 12139 5783 12142
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 6640 11933 6700 12142
rect 7097 12200 9463 12202
rect 7097 12144 7102 12200
rect 7158 12144 9402 12200
rect 9458 12144 9463 12200
rect 7097 12142 9463 12144
rect 7097 12139 7163 12142
rect 9397 12139 9463 12142
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 1393 11930 1459 11933
rect 0 11928 1459 11930
rect 0 11872 1398 11928
rect 1454 11872 1459 11928
rect 0 11870 1459 11872
rect 0 11840 800 11870
rect 1393 11867 1459 11870
rect 6637 11930 6703 11933
rect 10041 11930 10107 11933
rect 6637 11928 10107 11930
rect 6637 11872 6642 11928
rect 6698 11872 10046 11928
rect 10102 11872 10107 11928
rect 6637 11870 10107 11872
rect 6637 11867 6703 11870
rect 10041 11867 10107 11870
rect 13629 11930 13695 11933
rect 15929 11930 15995 11933
rect 13629 11928 15995 11930
rect 13629 11872 13634 11928
rect 13690 11872 15934 11928
rect 15990 11872 15995 11928
rect 13629 11870 15995 11872
rect 13629 11867 13695 11870
rect 15929 11867 15995 11870
rect 3969 11794 4035 11797
rect 17677 11794 17743 11797
rect 3969 11792 17743 11794
rect 3969 11736 3974 11792
rect 4030 11736 17682 11792
rect 17738 11736 17743 11792
rect 3969 11734 17743 11736
rect 3969 11731 4035 11734
rect 17677 11731 17743 11734
rect 3601 11658 3667 11661
rect 19609 11658 19675 11661
rect 3601 11656 19675 11658
rect 3601 11600 3606 11656
rect 3662 11600 19614 11656
rect 19670 11600 19675 11656
rect 3601 11598 19675 11600
rect 3601 11595 3667 11598
rect 19609 11595 19675 11598
rect 0 11522 800 11552
rect 1393 11522 1459 11525
rect 0 11520 1459 11522
rect 0 11464 1398 11520
rect 1454 11464 1459 11520
rect 0 11462 1459 11464
rect 0 11432 800 11462
rect 1393 11459 1459 11462
rect 21449 11522 21515 11525
rect 22200 11522 23000 11552
rect 21449 11520 23000 11522
rect 21449 11464 21454 11520
rect 21510 11464 23000 11520
rect 21449 11462 23000 11464
rect 21449 11459 21515 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 6177 11250 6243 11253
rect 13261 11250 13327 11253
rect 6177 11248 13327 11250
rect 6177 11192 6182 11248
rect 6238 11192 13266 11248
rect 13322 11192 13327 11248
rect 6177 11190 13327 11192
rect 6177 11187 6243 11190
rect 13261 11187 13327 11190
rect 0 11114 800 11144
rect 1485 11114 1551 11117
rect 0 11112 1551 11114
rect 0 11056 1490 11112
rect 1546 11056 1551 11112
rect 0 11054 1551 11056
rect 0 11024 800 11054
rect 1485 11051 1551 11054
rect 5349 11114 5415 11117
rect 11789 11114 11855 11117
rect 5349 11112 11855 11114
rect 5349 11056 5354 11112
rect 5410 11056 11794 11112
rect 11850 11056 11855 11112
rect 5349 11054 11855 11056
rect 5349 11051 5415 11054
rect 11789 11051 11855 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 1669 10842 1735 10845
rect 1669 10840 4906 10842
rect 1669 10784 1674 10840
rect 1730 10784 4906 10840
rect 1669 10782 4906 10784
rect 1669 10779 1735 10782
rect 0 10706 800 10736
rect 2773 10706 2839 10709
rect 0 10704 2839 10706
rect 0 10648 2778 10704
rect 2834 10648 2839 10704
rect 0 10646 2839 10648
rect 4846 10706 4906 10782
rect 6862 10780 6868 10844
rect 6932 10842 6938 10844
rect 6932 10782 7298 10842
rect 6932 10780 6938 10782
rect 7046 10706 7052 10708
rect 4846 10646 7052 10706
rect 0 10616 800 10646
rect 2773 10643 2839 10646
rect 7046 10644 7052 10646
rect 7116 10644 7122 10708
rect 7238 10706 7298 10782
rect 21081 10706 21147 10709
rect 7238 10704 21147 10706
rect 7238 10648 21086 10704
rect 21142 10648 21147 10704
rect 7238 10646 21147 10648
rect 21081 10643 21147 10646
rect 2681 10570 2747 10573
rect 15193 10570 15259 10573
rect 2681 10568 15259 10570
rect 2681 10512 2686 10568
rect 2742 10512 15198 10568
rect 15254 10512 15259 10568
rect 2681 10510 15259 10512
rect 2681 10507 2747 10510
rect 15193 10507 15259 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 5942 10236 5948 10300
rect 6012 10298 6018 10300
rect 7281 10298 7347 10301
rect 6012 10296 7347 10298
rect 6012 10240 7286 10296
rect 7342 10240 7347 10296
rect 6012 10238 7347 10240
rect 6012 10236 6018 10238
rect 7281 10235 7347 10238
rect 5257 10162 5323 10165
rect 19333 10162 19399 10165
rect 5257 10160 19399 10162
rect 5257 10104 5262 10160
rect 5318 10104 19338 10160
rect 19394 10104 19399 10160
rect 5257 10102 19399 10104
rect 5257 10099 5323 10102
rect 19333 10099 19399 10102
rect 2129 10026 2195 10029
rect 7097 10026 7163 10029
rect 2129 10024 7163 10026
rect 2129 9968 2134 10024
rect 2190 9968 7102 10024
rect 7158 9968 7163 10024
rect 2129 9966 7163 9968
rect 2129 9963 2195 9966
rect 7097 9963 7163 9966
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 13118 9556 13124 9620
rect 13188 9618 13194 9620
rect 15837 9618 15903 9621
rect 13188 9616 15903 9618
rect 13188 9560 15842 9616
rect 15898 9560 15903 9616
rect 13188 9558 15903 9560
rect 13188 9556 13194 9558
rect 15837 9555 15903 9558
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 9029 9482 9095 9485
rect 18137 9482 18203 9485
rect 9029 9480 18203 9482
rect 9029 9424 9034 9480
rect 9090 9424 18142 9480
rect 18198 9424 18203 9480
rect 9029 9422 18203 9424
rect 9029 9419 9095 9422
rect 18137 9419 18203 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 2773 9074 2839 9077
rect 15745 9074 15811 9077
rect 0 9014 1410 9074
rect 0 8984 800 9014
rect 1350 8805 1410 9014
rect 2773 9072 15811 9074
rect 2773 9016 2778 9072
rect 2834 9016 15750 9072
rect 15806 9016 15811 9072
rect 2773 9014 15811 9016
rect 2773 9011 2839 9014
rect 15745 9011 15811 9014
rect 3918 8876 3924 8940
rect 3988 8938 3994 8940
rect 6821 8938 6887 8941
rect 3988 8936 6887 8938
rect 3988 8880 6826 8936
rect 6882 8880 6887 8936
rect 3988 8878 6887 8880
rect 3988 8876 3994 8878
rect 6821 8875 6887 8878
rect 1350 8800 1459 8805
rect 1350 8744 1398 8800
rect 1454 8744 1459 8800
rect 1350 8742 1459 8744
rect 1393 8739 1459 8742
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 1853 8666 1919 8669
rect 10869 8668 10935 8669
rect 10869 8666 10916 8668
rect 0 8664 1919 8666
rect 0 8608 1858 8664
rect 1914 8608 1919 8664
rect 0 8606 1919 8608
rect 10824 8664 10916 8666
rect 10824 8608 10874 8664
rect 10824 8606 10916 8608
rect 0 8576 800 8606
rect 1853 8603 1919 8606
rect 10869 8604 10916 8606
rect 10980 8604 10986 8668
rect 10869 8603 10935 8604
rect 6545 8530 6611 8533
rect 10961 8530 11027 8533
rect 14365 8530 14431 8533
rect 6545 8528 14431 8530
rect 6545 8472 6550 8528
rect 6606 8472 10966 8528
rect 11022 8472 14370 8528
rect 14426 8472 14431 8528
rect 6545 8470 14431 8472
rect 6545 8467 6611 8470
rect 10961 8467 11027 8470
rect 14365 8467 14431 8470
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 5574 7924 5580 7988
rect 5644 7986 5650 7988
rect 7741 7986 7807 7989
rect 5644 7984 7807 7986
rect 5644 7928 7746 7984
rect 7802 7928 7807 7984
rect 5644 7926 7807 7928
rect 5644 7924 5650 7926
rect 7741 7923 7807 7926
rect 0 7850 800 7880
rect 1853 7850 1919 7853
rect 0 7848 1919 7850
rect 0 7792 1858 7848
rect 1914 7792 1919 7848
rect 0 7790 1919 7792
rect 0 7760 800 7790
rect 1853 7787 1919 7790
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 1853 7034 1919 7037
rect 0 7032 1919 7034
rect 0 6976 1858 7032
rect 1914 6976 1919 7032
rect 0 6974 1919 6976
rect 0 6944 800 6974
rect 1853 6971 1919 6974
rect 5901 6762 5967 6765
rect 12934 6762 12940 6764
rect 5901 6760 12940 6762
rect 5901 6704 5906 6760
rect 5962 6704 12940 6760
rect 5901 6702 12940 6704
rect 5901 6699 5967 6702
rect 12934 6700 12940 6702
rect 13004 6700 13010 6764
rect 0 6626 800 6656
rect 1393 6626 1459 6629
rect 0 6624 1459 6626
rect 0 6568 1398 6624
rect 1454 6568 1459 6624
rect 0 6566 1459 6568
rect 0 6536 800 6566
rect 1393 6563 1459 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 0 5810 800 5840
rect 1853 5810 1919 5813
rect 0 5808 1919 5810
rect 0 5752 1858 5808
rect 1914 5752 1919 5808
rect 0 5750 1919 5752
rect 0 5720 800 5750
rect 1853 5747 1919 5750
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 1393 5402 1459 5405
rect 0 5400 1459 5402
rect 0 5344 1398 5400
rect 1454 5344 1459 5400
rect 0 5342 1459 5344
rect 0 5312 800 5342
rect 1393 5339 1459 5342
rect 0 4994 800 5024
rect 2221 4994 2287 4997
rect 0 4992 2287 4994
rect 0 4936 2226 4992
rect 2282 4936 2287 4992
rect 0 4934 2287 4936
rect 0 4904 800 4934
rect 2221 4931 2287 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 0 4586 800 4616
rect 2221 4586 2287 4589
rect 0 4584 2287 4586
rect 0 4528 2226 4584
rect 2282 4528 2287 4584
rect 0 4526 2287 4528
rect 0 4496 800 4526
rect 2221 4523 2287 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 2037 3770 2103 3773
rect 0 3768 2103 3770
rect 0 3712 2042 3768
rect 2098 3712 2103 3768
rect 0 3710 2103 3712
rect 0 3680 800 3710
rect 2037 3707 2103 3710
rect 0 3362 800 3392
rect 1485 3362 1551 3365
rect 0 3360 1551 3362
rect 0 3304 1490 3360
rect 1546 3304 1551 3360
rect 0 3302 1551 3304
rect 0 3272 800 3302
rect 1485 3299 1551 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 0 2954 800 2984
rect 1485 2954 1551 2957
rect 0 2952 1551 2954
rect 0 2896 1490 2952
rect 1546 2896 1551 2952
rect 0 2894 1551 2896
rect 0 2864 800 2894
rect 1485 2891 1551 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 0 2546 800 2576
rect 2037 2546 2103 2549
rect 0 2544 2103 2546
rect 0 2488 2042 2544
rect 2098 2488 2103 2544
rect 0 2486 2103 2488
rect 0 2456 800 2486
rect 2037 2483 2103 2486
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 800 2078
rect 2773 2075 2839 2078
rect 0 1730 800 1760
rect 2221 1730 2287 1733
rect 0 1728 2287 1730
rect 0 1672 2226 1728
rect 2282 1672 2287 1728
rect 0 1670 2287 1672
rect 0 1640 800 1670
rect 2221 1667 2287 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3924 19484 3988 19548
rect 8524 19544 8588 19548
rect 8524 19488 8538 19544
rect 8538 19488 8588 19544
rect 8524 19484 8588 19488
rect 5580 19408 5644 19412
rect 5580 19352 5594 19408
rect 5594 19352 5644 19408
rect 5580 19348 5644 19352
rect 5948 19408 6012 19412
rect 5948 19352 5998 19408
rect 5998 19352 6012 19408
rect 5948 19348 6012 19352
rect 10916 19408 10980 19412
rect 10916 19352 10966 19408
rect 10966 19352 10980 19408
rect 10916 19348 10980 19352
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6684 18804 6748 18868
rect 5396 18668 5460 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 7052 18048 7116 18052
rect 7052 17992 7066 18048
rect 7066 17992 7116 18048
rect 7052 17988 7116 17992
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 13124 17172 13188 17236
rect 6868 17036 6932 17100
rect 8340 17036 8404 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 12940 16144 13004 16148
rect 12940 16088 12990 16144
rect 12990 16088 13004 16144
rect 12940 16084 13004 16088
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6684 14588 6748 14652
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 2084 13908 2148 13972
rect 8340 13772 8404 13836
rect 8524 13772 8588 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 5396 12956 5460 13020
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 2084 12140 2148 12204
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 6868 10780 6932 10844
rect 7052 10644 7116 10708
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5948 10236 6012 10300
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 13124 9556 13188 9620
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 3924 8876 3988 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 10916 8664 10980 8668
rect 10916 8608 10930 8664
rect 10930 8608 10980 8664
rect 10916 8604 10980 8608
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 5580 7924 5644 7988
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 12940 6700 13004 6764
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 3923 19548 3989 19549
rect 3923 19484 3924 19548
rect 3988 19484 3989 19548
rect 3923 19483 3989 19484
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 2083 13972 2149 13973
rect 2083 13908 2084 13972
rect 2148 13908 2149 13972
rect 2083 13907 2149 13908
rect 2086 12205 2146 13907
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 2083 12204 2149 12205
rect 2083 12140 2084 12204
rect 2148 12140 2149 12204
rect 2083 12139 2149 12140
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3926 8941 3986 19483
rect 5579 19412 5645 19413
rect 5579 19348 5580 19412
rect 5644 19348 5645 19412
rect 5579 19347 5645 19348
rect 5947 19412 6013 19413
rect 5947 19348 5948 19412
rect 6012 19348 6013 19412
rect 5947 19347 6013 19348
rect 5395 18732 5461 18733
rect 5395 18668 5396 18732
rect 5460 18668 5461 18732
rect 5395 18667 5461 18668
rect 5398 13021 5458 18667
rect 5395 13020 5461 13021
rect 5395 12956 5396 13020
rect 5460 12956 5461 13020
rect 5395 12955 5461 12956
rect 3923 8940 3989 8941
rect 3923 8876 3924 8940
rect 3988 8876 3989 8940
rect 3923 8875 3989 8876
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 5582 7989 5642 19347
rect 5950 10301 6010 19347
rect 6142 18528 6462 19552
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8523 19548 8589 19549
rect 8523 19484 8524 19548
rect 8588 19484 8589 19548
rect 8523 19483 8589 19484
rect 6683 18868 6749 18869
rect 6683 18804 6684 18868
rect 6748 18804 6749 18868
rect 6683 18803 6749 18804
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6686 14653 6746 18803
rect 7051 18052 7117 18053
rect 7051 17988 7052 18052
rect 7116 17988 7117 18052
rect 7051 17987 7117 17988
rect 6867 17100 6933 17101
rect 6867 17036 6868 17100
rect 6932 17036 6933 17100
rect 6867 17035 6933 17036
rect 6683 14652 6749 14653
rect 6683 14588 6684 14652
rect 6748 14588 6749 14652
rect 6683 14587 6749 14588
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5947 10300 6013 10301
rect 5947 10236 5948 10300
rect 6012 10236 6013 10300
rect 5947 10235 6013 10236
rect 6142 9824 6462 10848
rect 6870 10845 6930 17035
rect 6867 10844 6933 10845
rect 6867 10780 6868 10844
rect 6932 10780 6933 10844
rect 6867 10779 6933 10780
rect 7054 10709 7114 17987
rect 8339 17100 8405 17101
rect 8339 17036 8340 17100
rect 8404 17036 8405 17100
rect 8339 17035 8405 17036
rect 8342 13837 8402 17035
rect 8526 13837 8586 19483
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 10915 19412 10981 19413
rect 10915 19348 10916 19412
rect 10980 19348 10981 19412
rect 10915 19347 10981 19348
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8339 13836 8405 13837
rect 8339 13772 8340 13836
rect 8404 13772 8405 13836
rect 8339 13771 8405 13772
rect 8523 13836 8589 13837
rect 8523 13772 8524 13836
rect 8588 13772 8589 13836
rect 8523 13771 8589 13772
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 7051 10708 7117 10709
rect 7051 10644 7052 10708
rect 7116 10644 7117 10708
rect 7051 10643 7117 10644
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 5579 7988 5645 7989
rect 5579 7924 5580 7988
rect 5644 7924 5645 7988
rect 5579 7923 5645 7924
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 10918 8669 10978 19347
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13123 17236 13189 17237
rect 13123 17172 13124 17236
rect 13188 17172 13189 17236
rect 13123 17171 13189 17172
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 12939 16148 13005 16149
rect 12939 16084 12940 16148
rect 13004 16084 13005 16148
rect 12939 16083 13005 16084
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 10915 8668 10981 8669
rect 10915 8604 10916 8668
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 12942 6765 13002 16083
rect 13126 9621 13186 17171
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13123 9620 13189 9621
rect 13123 9556 13124 9620
rect 13188 9556 13189 9620
rect 13123 9555 13189 9556
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 12939 6764 13005 6765
rect 12939 6700 12940 6764
rect 13004 6700 13005 6764
rect 12939 6699 13005 6700
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 2024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 12052 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 8280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 11040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 11132 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19964 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 21160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 20700 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9844 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7360 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 3036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 4048 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform -1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform -1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 13064 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43
timestamp 1649977179
transform 1 0 5060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1649977179
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp 1649977179
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1649977179
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_17
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_29
timestamp 1649977179
transform 1 0 3772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_41
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_14
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1649977179
transform 1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_72
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_14
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_113
timestamp 1649977179
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_88
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_92
timestamp 1649977179
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_102
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_132
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_123
timestamp 1649977179
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_199
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_205
timestamp 1649977179
transform 1 0 19964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_211
timestamp 1649977179
transform 1 0 20516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1649977179
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_13
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_31
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_40
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_187
timestamp 1649977179
transform 1 0 18308 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_213
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_12
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_46
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_51
timestamp 1649977179
transform 1 0 5796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_200
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_204
timestamp 1649977179
transform 1 0 19872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1649977179
transform 1 0 3036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1649977179
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1649977179
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_6
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_17
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1649977179
transform 1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1649977179
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_12
timestamp 1649977179
transform 1 0 2208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1649977179
transform 1 0 3312 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_32
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_60
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1649977179
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_177
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_10
timestamp 1649977179
transform 1 0 2024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_14
timestamp 1649977179
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_68
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_76
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_99
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_171
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_5
timestamp 1649977179
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1649977179
transform 1 0 2024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1649977179
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1649977179
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_6
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_10
timestamp 1649977179
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_40
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_52
timestamp 1649977179
transform 1 0 5888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1649977179
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_216
timestamp 1649977179
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_34
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1649977179
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1649977179
transform 1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_94
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_116
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_188
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_17
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1649977179
transform 1 0 3036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_59
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_103
timestamp 1649977179
transform 1 0 10580 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1649977179
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1649977179
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1649977179
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1649977179
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_102
timestamp 1649977179
transform 1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_119
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1649977179
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1649977179
transform 1 0 13064 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_101
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_126
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1649977179
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_31
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1649977179
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1649977179
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1649977179
transform 1 0 2576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1649977179
transform 1 0 9200 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_119
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1649977179
transform 1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_163
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1649977179
transform 1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1649977179
transform 1 0 6256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1649977179
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1649977179
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_94
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1649977179
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1649977179
transform 1 0 10856 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1649977179
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_191
timestamp 1649977179
transform 1 0 18676 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_203
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1649977179
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_22
timestamp 1649977179
transform 1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1649977179
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1649977179
transform 1 0 4784 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_50
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_63
timestamp 1649977179
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1649977179
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1649977179
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1649977179
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1649977179
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_13
timestamp 1649977179
transform 1 0 2300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_18
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1649977179
transform 1 0 4048 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_51
timestamp 1649977179
transform 1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_56
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1649977179
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_89
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1649977179
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1649977179
transform 1 0 11592 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_183
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_28
timestamp 1649977179
transform 1 0 3680 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_32
timestamp 1649977179
transform 1 0 4048 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1649977179
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_45
timestamp 1649977179
transform 1 0 5244 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_88
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_103
timestamp 1649977179
transform 1 0 10580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1649977179
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1649977179
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_201
timestamp 1649977179
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_34
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_44
timestamp 1649977179
transform 1 0 5152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_94
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_108
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1649977179
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_154
timestamp 1649977179
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_160
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_25
timestamp 1649977179
transform 1 0 3404 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_33
timestamp 1649977179
transform 1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_44
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_66
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_89
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_100
timestamp 1649977179
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_119
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_124
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1649977179
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _068_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform -1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 8740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 6900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 6072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 9292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 11500 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 21160 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 3496 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 8188 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 8648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 9292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 12696 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 5152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 3312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18308 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16744 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17572 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21344 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14628 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13616 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16100 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13616 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17204 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14996 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17204 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20976 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20516 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19136 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18676 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18032 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16100 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13892 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_1__124 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_1__101
timestamp 1649977179
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_1__107
timestamp 1649977179
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l2_in_1__108
timestamp 1649977179
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l1_in_1__109
timestamp 1649977179
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_0__125
timestamp 1649977179
transform -1 0 11224 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_0__126
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_0__127
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_0__128
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l2_in_0__129
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l2_in_0__130
timestamp 1649977179
transform -1 0 6348 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__132
timestamp 1649977179
transform -1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_27.mux_l2_in_0__133
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__134
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__102
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__103
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__104
timestamp 1649977179
transform -1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__105
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__106
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_1__110
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7636 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2852 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_1__116
timestamp 1649977179
transform 1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5704 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_1__121
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8096 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_6.mux_l2_in_1__122
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l1_in_1__123
timestamp 1649977179
transform -1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5888 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_10.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7452 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_12.mux_l2_in_0__112
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10304 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5060 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_14.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7452 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_0__114
timestamp 1649977179
transform -1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_18.mux_l2_in_0__115
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11316 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_20.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9568 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6808 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_22.mux_l2_in_0__118
timestamp 1649977179
transform 1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l1_in_1__119
timestamp 1649977179
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_26.mux_l2_in_0__120
timestamp 1649977179
transform -1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 1932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 3404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 4 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 5 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 6 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 7 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 8 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 9 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 10 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 11 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 12 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 13 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 14 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 15 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 16 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 17 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 18 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 19 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 20 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 21 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 22 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 23 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 24 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 25 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 26 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 27 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 28 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 29 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 30 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 31 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 32 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 33 nsew signal tristate
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 34 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 44 nsew signal input
flabel metal2 s 8482 22200 8538 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 45 nsew signal input
flabel metal2 s 8942 22200 8998 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 46 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 47 nsew signal input
flabel metal2 s 9862 22200 9918 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 48 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 49 nsew signal input
flabel metal2 s 10782 22200 10838 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 50 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 51 nsew signal input
flabel metal2 s 11702 22200 11758 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 52 nsew signal input
flabel metal2 s 12162 22200 12218 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 53 nsew signal input
flabel metal2 s 12622 22200 12678 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 54 nsew signal input
flabel metal2 s 4342 22200 4398 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 55 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 56 nsew signal input
flabel metal2 s 5262 22200 5318 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 57 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 58 nsew signal input
flabel metal2 s 6182 22200 6238 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 59 nsew signal input
flabel metal2 s 6642 22200 6698 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 60 nsew signal input
flabel metal2 s 7102 22200 7158 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 61 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 62 nsew signal input
flabel metal2 s 8022 22200 8078 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 63 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 64 nsew signal tristate
flabel metal2 s 17682 22200 17738 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 65 nsew signal tristate
flabel metal2 s 18142 22200 18198 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 66 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 67 nsew signal tristate
flabel metal2 s 19062 22200 19118 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 68 nsew signal tristate
flabel metal2 s 19522 22200 19578 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 69 nsew signal tristate
flabel metal2 s 19982 22200 20038 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 70 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 71 nsew signal tristate
flabel metal2 s 20902 22200 20958 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 72 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 73 nsew signal tristate
flabel metal2 s 21822 22200 21878 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 74 nsew signal tristate
flabel metal2 s 13542 22200 13598 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 75 nsew signal tristate
flabel metal2 s 14002 22200 14058 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 76 nsew signal tristate
flabel metal2 s 14462 22200 14518 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 77 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 78 nsew signal tristate
flabel metal2 s 15382 22200 15438 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 79 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 80 nsew signal tristate
flabel metal2 s 16302 22200 16358 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 81 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 82 nsew signal tristate
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 83 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_11_
port 84 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_13_
port 85 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_15_
port 86 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 left_bottom_grid_pin_17_
port 87 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_1_
port 88 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_3_
port 89 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_5_
port 90 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_7_
port 91 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_9_
port 92 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 93 nsew signal input
flabel metal2 s 202 22200 258 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 94 nsew signal input
flabel metal2 s 662 22200 718 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 95 nsew signal input
flabel metal2 s 1122 22200 1178 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 96 nsew signal input
flabel metal2 s 1582 22200 1638 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 97 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 98 nsew signal input
flabel metal2 s 2502 22200 2558 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 99 nsew signal input
flabel metal2 s 2962 22200 3018 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 100 nsew signal input
flabel metal2 s 3422 22200 3478 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 101 nsew signal input
flabel metal2 s 22742 22200 22798 23000 0 FreeSans 224 90 0 0 top_right_grid_pin_1_
port 102 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
