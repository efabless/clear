magic
tech sky130A
magscale 1 2
timestamp 1656943210
<< obsli1 >>
rect 1104 2159 16008 17425
<< obsm1 >>
rect 1026 1436 16178 18012
<< metal2 >>
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11702 19200 11758 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
<< obsm2 >>
rect 1142 19144 1342 19258
rect 1510 19144 1710 19258
rect 1878 19144 2078 19258
rect 2246 19144 2446 19258
rect 2614 19144 2814 19258
rect 2982 19144 3182 19258
rect 3350 19144 3550 19258
rect 3718 19144 3918 19258
rect 4086 19144 4286 19258
rect 4454 19144 4654 19258
rect 4822 19144 5022 19258
rect 5190 19144 5390 19258
rect 5558 19144 5758 19258
rect 5926 19144 6126 19258
rect 6294 19144 6494 19258
rect 6662 19144 6862 19258
rect 7030 19144 7230 19258
rect 7398 19144 7598 19258
rect 7766 19144 7966 19258
rect 8134 19144 8334 19258
rect 8502 19144 8702 19258
rect 8870 19144 9070 19258
rect 9238 19144 9438 19258
rect 9606 19144 9806 19258
rect 9974 19144 10174 19258
rect 10342 19144 10542 19258
rect 10710 19144 10910 19258
rect 11078 19144 11278 19258
rect 11446 19144 11646 19258
rect 11814 19144 12014 19258
rect 12182 19144 12382 19258
rect 12550 19144 12750 19258
rect 12918 19144 13118 19258
rect 13286 19144 13486 19258
rect 13654 19144 13854 19258
rect 14022 19144 14222 19258
rect 14390 19144 14590 19258
rect 14758 19144 14958 19258
rect 15126 19144 15326 19258
rect 15494 19144 15694 19258
rect 15862 19144 16062 19258
rect 1032 856 16172 19144
rect 1032 734 1158 856
rect 1326 734 1526 856
rect 1694 734 1894 856
rect 2062 734 2262 856
rect 2430 734 2630 856
rect 2798 734 2998 856
rect 3166 734 3366 856
rect 3534 734 3734 856
rect 3902 734 4102 856
rect 4270 734 4470 856
rect 4638 734 4838 856
rect 5006 734 5206 856
rect 5374 734 5574 856
rect 5742 734 5942 856
rect 6110 734 6310 856
rect 6478 734 6678 856
rect 6846 734 7046 856
rect 7214 734 7414 856
rect 7582 734 7782 856
rect 7950 734 8150 856
rect 8318 734 8518 856
rect 8686 734 8886 856
rect 9054 734 9254 856
rect 9422 734 9622 856
rect 9790 734 9990 856
rect 10158 734 10358 856
rect 10526 734 10726 856
rect 10894 734 11094 856
rect 11262 734 11462 856
rect 11630 734 11830 856
rect 11998 734 12198 856
rect 12366 734 12566 856
rect 12734 734 12934 856
rect 13102 734 13302 856
rect 13470 734 13670 856
rect 13838 734 14038 856
rect 14206 734 14406 856
rect 14574 734 14774 856
rect 14942 734 15142 856
rect 15310 734 15510 856
rect 15678 734 15878 856
rect 16046 734 16172 856
<< metal3 >>
rect 0 19456 800 19576
rect 0 18504 800 18624
rect 16400 17824 17200 17944
rect 0 17552 800 17672
rect 0 16600 800 16720
rect 0 15648 800 15768
rect 0 14696 800 14816
rect 0 13744 800 13864
rect 16400 13880 17200 14000
rect 0 12792 800 12912
rect 0 11840 800 11960
rect 0 10888 800 11008
rect 0 9936 800 10056
rect 16400 9936 17200 10056
rect 0 8984 800 9104
rect 0 8032 800 8152
rect 0 7080 800 7200
rect 0 6128 800 6248
rect 16400 5992 17200 6112
rect 0 5176 800 5296
rect 0 4224 800 4344
rect 0 3272 800 3392
rect 0 2320 800 2440
rect 16400 2048 17200 2168
rect 0 1368 800 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 19376 16400 19546
rect 800 18704 16400 19376
rect 880 18424 16400 18704
rect 800 18024 16400 18424
rect 800 17752 16320 18024
rect 880 17744 16320 17752
rect 880 17472 16400 17744
rect 800 16800 16400 17472
rect 880 16520 16400 16800
rect 800 15848 16400 16520
rect 880 15568 16400 15848
rect 800 14896 16400 15568
rect 880 14616 16400 14896
rect 800 14080 16400 14616
rect 800 13944 16320 14080
rect 880 13800 16320 13944
rect 880 13664 16400 13800
rect 800 12992 16400 13664
rect 880 12712 16400 12992
rect 800 12040 16400 12712
rect 880 11760 16400 12040
rect 800 11088 16400 11760
rect 880 10808 16400 11088
rect 800 10136 16400 10808
rect 880 9856 16320 10136
rect 800 9184 16400 9856
rect 880 8904 16400 9184
rect 800 8232 16400 8904
rect 880 7952 16400 8232
rect 800 7280 16400 7952
rect 880 7000 16400 7280
rect 800 6328 16400 7000
rect 880 6192 16400 6328
rect 880 6048 16320 6192
rect 800 5912 16320 6048
rect 800 5376 16400 5912
rect 880 5096 16400 5376
rect 800 4424 16400 5096
rect 880 4144 16400 4424
rect 800 3472 16400 4144
rect 880 3192 16400 3472
rect 800 2520 16400 3192
rect 880 2248 16400 2520
rect 880 2240 16320 2248
rect 800 1968 16320 2240
rect 800 1568 16400 1968
rect 880 1288 16400 1568
rect 800 616 16400 1288
rect 880 446 16400 616
<< metal4 >>
rect 2818 2128 3138 17456
rect 4692 2128 5012 17456
rect 6566 2128 6886 17456
rect 8440 2128 8760 17456
rect 10314 2128 10634 17456
rect 12188 2128 12508 17456
rect 14062 2128 14382 17456
<< obsm4 >>
rect 3371 2211 4612 17237
rect 5092 2211 6486 17237
rect 6966 2211 8360 17237
rect 8840 2211 10234 17237
rect 10714 2211 12108 17237
rect 12588 2211 13982 17237
rect 14462 2211 15029 17237
<< labels >>
rlabel metal2 s 1030 19200 1086 20000 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 3 nsew power bidirectional
rlabel metal3 s 0 1368 800 1488 6 ccff_head
port 4 nsew signal input
rlabel metal3 s 16400 2048 17200 2168 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[0]
port 6 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[10]
port 7 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[11]
port 8 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_in[12]
port 9 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 chany_bottom_in[13]
port 10 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_in[14]
port 11 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_in[15]
port 12 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_in[16]
port 13 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_in[17]
port 14 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_in[18]
port 15 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 chany_bottom_in[19]
port 16 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[1]
port 17 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 chany_bottom_in[2]
port 18 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[3]
port 19 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[4]
port 20 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[5]
port 21 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[6]
port 22 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[7]
port 23 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 chany_bottom_in[8]
port 24 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[9]
port 25 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 chany_bottom_out[0]
port 26 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[10]
port 27 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_out[11]
port 28 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_out[12]
port 29 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_out[13]
port 30 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_out[14]
port 31 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_out[15]
port 32 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 chany_bottom_out[16]
port 33 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_out[17]
port 34 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_out[18]
port 35 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_out[19]
port 36 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 chany_bottom_out[1]
port 37 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 chany_bottom_out[2]
port 38 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[3]
port 39 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[4]
port 40 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_out[5]
port 41 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_out[6]
port 42 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_out[7]
port 43 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_out[8]
port 44 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[9]
port 45 nsew signal output
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_in[0]
port 46 nsew signal input
rlabel metal2 s 12438 19200 12494 20000 6 chany_top_in[10]
port 47 nsew signal input
rlabel metal2 s 12806 19200 12862 20000 6 chany_top_in[11]
port 48 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[12]
port 49 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[13]
port 50 nsew signal input
rlabel metal2 s 13910 19200 13966 20000 6 chany_top_in[14]
port 51 nsew signal input
rlabel metal2 s 14278 19200 14334 20000 6 chany_top_in[15]
port 52 nsew signal input
rlabel metal2 s 14646 19200 14702 20000 6 chany_top_in[16]
port 53 nsew signal input
rlabel metal2 s 15014 19200 15070 20000 6 chany_top_in[17]
port 54 nsew signal input
rlabel metal2 s 15382 19200 15438 20000 6 chany_top_in[18]
port 55 nsew signal input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[19]
port 56 nsew signal input
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_in[1]
port 57 nsew signal input
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_in[2]
port 58 nsew signal input
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[3]
port 59 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[4]
port 60 nsew signal input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[5]
port 61 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[6]
port 62 nsew signal input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[7]
port 63 nsew signal input
rlabel metal2 s 11702 19200 11758 20000 6 chany_top_in[8]
port 64 nsew signal input
rlabel metal2 s 12070 19200 12126 20000 6 chany_top_in[9]
port 65 nsew signal input
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[0]
port 66 nsew signal output
rlabel metal2 s 5078 19200 5134 20000 6 chany_top_out[10]
port 67 nsew signal output
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[11]
port 68 nsew signal output
rlabel metal2 s 5814 19200 5870 20000 6 chany_top_out[12]
port 69 nsew signal output
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[13]
port 70 nsew signal output
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[14]
port 71 nsew signal output
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[15]
port 72 nsew signal output
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[16]
port 73 nsew signal output
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[17]
port 74 nsew signal output
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[18]
port 75 nsew signal output
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[19]
port 76 nsew signal output
rlabel metal2 s 1766 19200 1822 20000 6 chany_top_out[1]
port 77 nsew signal output
rlabel metal2 s 2134 19200 2190 20000 6 chany_top_out[2]
port 78 nsew signal output
rlabel metal2 s 2502 19200 2558 20000 6 chany_top_out[3]
port 79 nsew signal output
rlabel metal2 s 2870 19200 2926 20000 6 chany_top_out[4]
port 80 nsew signal output
rlabel metal2 s 3238 19200 3294 20000 6 chany_top_out[5]
port 81 nsew signal output
rlabel metal2 s 3606 19200 3662 20000 6 chany_top_out[6]
port 82 nsew signal output
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[7]
port 83 nsew signal output
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[8]
port 84 nsew signal output
rlabel metal2 s 4710 19200 4766 20000 6 chany_top_out[9]
port 85 nsew signal output
rlabel metal3 s 16400 9936 17200 10056 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 86 nsew signal output
rlabel metal3 s 16400 13880 17200 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 87 nsew signal input
rlabel metal3 s 16400 17824 17200 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 88 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 left_grid_pin_16_
port 89 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 left_grid_pin_17_
port 90 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 left_grid_pin_18_
port 91 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 left_grid_pin_19_
port 92 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 left_grid_pin_20_
port 93 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 left_grid_pin_21_
port 94 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 left_grid_pin_22_
port 95 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 left_grid_pin_23_
port 96 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 left_grid_pin_24_
port 97 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 left_grid_pin_25_
port 98 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 left_grid_pin_26_
port 99 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 left_grid_pin_27_
port 100 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 left_grid_pin_28_
port 101 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 left_grid_pin_29_
port 102 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 left_grid_pin_30_
port 103 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 left_grid_pin_31_
port 104 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 left_width_0_height_0__pin_0_
port 105 nsew signal input
rlabel metal3 s 0 416 800 536 6 left_width_0_height_0__pin_1_lower
port 106 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 left_width_0_height_0__pin_1_upper
port 107 nsew signal output
rlabel metal2 s 16118 19200 16174 20000 6 prog_clk_0_N_out
port 108 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 prog_clk_0_S_out
port 109 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 prog_clk_0_W_in
port 110 nsew signal input
rlabel metal3 s 16400 5992 17200 6112 6 right_grid_pin_0_
port 111 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 17200 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1123424
string GDS_FILE /home/marwan/clear_signoff_final/openlane/cby_2__1_/runs/cby_2__1_/results/signoff/cby_2__1_.magic.gds
string GDS_START 84912
<< end >>

