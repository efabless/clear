magic
tech sky130A
magscale 1 2
timestamp 1681041682
<< viali >>
rect 3985 24361 4019 24395
rect 9137 24361 9171 24395
rect 21281 24361 21315 24395
rect 3249 24225 3283 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 14473 24225 14507 24259
rect 17325 24225 17359 24259
rect 17509 24225 17543 24259
rect 18521 24225 18555 24259
rect 18705 24225 18739 24259
rect 20085 24225 20119 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7297 24157 7331 24191
rect 9321 24157 9355 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14197 24157 14231 24191
rect 14749 24157 14783 24191
rect 15945 24157 15979 24191
rect 21465 24157 21499 24191
rect 22293 24157 22327 24191
rect 24961 24157 24995 24191
rect 25053 24157 25087 24191
rect 1593 24089 1627 24123
rect 5825 24089 5859 24123
rect 18429 24089 18463 24123
rect 19901 24089 19935 24123
rect 22569 24089 22603 24123
rect 1777 24021 1811 24055
rect 6561 24021 6595 24055
rect 11713 24021 11747 24055
rect 15761 24021 15795 24055
rect 16221 24021 16255 24055
rect 16405 24021 16439 24055
rect 16865 24021 16899 24055
rect 17233 24021 17267 24055
rect 18061 24021 18095 24055
rect 19349 24021 19383 24055
rect 19441 24021 19475 24055
rect 19809 24021 19843 24055
rect 20637 24021 20671 24055
rect 21925 24021 21959 24055
rect 24041 24021 24075 24055
rect 24593 24021 24627 24055
rect 2329 23817 2363 23851
rect 2513 23817 2547 23851
rect 11621 23817 11655 23851
rect 11805 23817 11839 23851
rect 13829 23817 13863 23851
rect 14105 23817 14139 23851
rect 14473 23817 14507 23851
rect 24041 23817 24075 23851
rect 3985 23749 4019 23783
rect 5825 23749 5859 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 15209 23749 15243 23783
rect 15393 23749 15427 23783
rect 15945 23749 15979 23783
rect 16037 23749 16071 23783
rect 17233 23749 17267 23783
rect 24317 23749 24351 23783
rect 25145 23749 25179 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6653 23681 6687 23715
rect 6929 23681 6963 23715
rect 7941 23681 7975 23715
rect 9965 23681 9999 23715
rect 12081 23681 12115 23715
rect 17325 23681 17359 23715
rect 12541 23613 12575 23647
rect 14565 23613 14599 23647
rect 14749 23613 14783 23647
rect 16221 23613 16255 23647
rect 17509 23613 17543 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 20269 23613 20303 23647
rect 20637 23613 20671 23647
rect 20913 23613 20947 23647
rect 22293 23613 22327 23647
rect 22569 23613 22603 23647
rect 24685 23613 24719 23647
rect 1869 23545 1903 23579
rect 24593 23545 24627 23579
rect 15577 23477 15611 23511
rect 16865 23477 16899 23511
rect 19809 23477 19843 23511
rect 20085 23477 20119 23511
rect 21833 23477 21867 23511
rect 25237 23477 25271 23511
rect 1593 23273 1627 23307
rect 1777 23205 1811 23239
rect 23397 23205 23431 23239
rect 3249 23137 3283 23171
rect 6561 23137 6595 23171
rect 8217 23137 8251 23171
rect 10517 23137 10551 23171
rect 12173 23137 12207 23171
rect 15301 23137 15335 23171
rect 17785 23137 17819 23171
rect 18705 23137 18739 23171
rect 19717 23137 19751 23171
rect 21649 23137 21683 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 4077 23069 4111 23103
rect 4353 23069 4387 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 9413 23069 9447 23103
rect 9873 23069 9907 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 14381 23001 14415 23035
rect 17693 23001 17727 23035
rect 18521 23001 18555 23035
rect 21925 23001 21959 23035
rect 9229 22933 9263 22967
rect 13553 22933 13587 22967
rect 14473 22933 14507 22967
rect 16773 22933 16807 22967
rect 17233 22933 17267 22967
rect 18981 22933 19015 22967
rect 21189 22933 21223 22967
rect 23857 22933 23891 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 1685 22729 1719 22763
rect 7205 22729 7239 22763
rect 13093 22729 13127 22763
rect 15393 22729 15427 22763
rect 18613 22729 18647 22763
rect 19257 22729 19291 22763
rect 2145 22661 2179 22695
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 6653 22661 6687 22695
rect 8769 22661 8803 22695
rect 12173 22661 12207 22695
rect 15945 22661 15979 22695
rect 17141 22661 17175 22695
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6837 22593 6871 22627
rect 7573 22593 7607 22627
rect 12081 22593 12115 22627
rect 13001 22593 13035 22627
rect 13645 22593 13679 22627
rect 16865 22593 16899 22627
rect 19165 22593 19199 22627
rect 20085 22593 20119 22627
rect 22017 22593 22051 22627
rect 1593 22525 1627 22559
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 12265 22525 12299 22559
rect 13921 22525 13955 22559
rect 20545 22525 20579 22559
rect 22293 22525 22327 22559
rect 23305 22525 23339 22559
rect 23581 22525 23615 22559
rect 11161 22457 11195 22491
rect 16129 22457 16163 22491
rect 16497 22457 16531 22491
rect 2237 22389 2271 22423
rect 11713 22389 11747 22423
rect 19625 22389 19659 22423
rect 25053 22389 25087 22423
rect 25421 22389 25455 22423
rect 14552 22185 14586 22219
rect 18797 22185 18831 22219
rect 19625 22185 19659 22219
rect 20624 22185 20658 22219
rect 16497 22117 16531 22151
rect 18981 22117 19015 22151
rect 1685 22049 1719 22083
rect 2881 22049 2915 22083
rect 6101 22049 6135 22083
rect 8125 22049 8159 22083
rect 10701 22049 10735 22083
rect 12449 22049 12483 22083
rect 17049 22049 17083 22083
rect 18153 22049 18187 22083
rect 18245 22049 18279 22083
rect 22569 22049 22603 22083
rect 23443 22049 23477 22083
rect 25237 22049 25271 22083
rect 2237 21981 2271 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 5549 21981 5583 22015
rect 7389 21981 7423 22015
rect 8953 21981 8987 22015
rect 9505 21981 9539 22015
rect 13093 21981 13127 22015
rect 14289 21981 14323 22015
rect 20361 21981 20395 22015
rect 23213 21981 23247 22015
rect 24961 21981 24995 22015
rect 10977 21913 11011 21947
rect 12909 21913 12943 21947
rect 13553 21913 13587 21947
rect 19533 21913 19567 21947
rect 9321 21845 9355 21879
rect 10057 21845 10091 21879
rect 13645 21845 13679 21879
rect 16037 21845 16071 21879
rect 16865 21845 16899 21879
rect 16957 21845 16991 21879
rect 17693 21845 17727 21879
rect 18061 21845 18095 21879
rect 19993 21845 20027 21879
rect 22109 21845 22143 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 11161 21641 11195 21675
rect 11345 21641 11379 21675
rect 11989 21641 12023 21675
rect 12265 21641 12299 21675
rect 12633 21641 12667 21675
rect 12725 21641 12759 21675
rect 13829 21641 13863 21675
rect 15025 21641 15059 21675
rect 20453 21641 20487 21675
rect 20913 21641 20947 21675
rect 22477 21641 22511 21675
rect 1685 21573 1719 21607
rect 2145 21573 2179 21607
rect 11621 21573 11655 21607
rect 14197 21573 14231 21607
rect 18245 21573 18279 21607
rect 21465 21573 21499 21607
rect 23673 21573 23707 21607
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 6745 21505 6779 21539
rect 7389 21505 7423 21539
rect 9045 21505 9079 21539
rect 15393 21505 15427 21539
rect 15485 21505 15519 21539
rect 17417 21505 17451 21539
rect 20821 21505 20855 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 7665 21437 7699 21471
rect 9321 21437 9355 21471
rect 12817 21437 12851 21471
rect 14289 21437 14323 21471
rect 14473 21437 14507 21471
rect 15669 21437 15703 21471
rect 16037 21437 16071 21471
rect 17509 21437 17543 21471
rect 17693 21437 17727 21471
rect 21005 21437 21039 21471
rect 22569 21437 22603 21471
rect 1869 21369 1903 21403
rect 11805 21369 11839 21403
rect 13369 21369 13403 21403
rect 22017 21369 22051 21403
rect 6561 21301 6595 21335
rect 10793 21301 10827 21335
rect 13461 21301 13495 21335
rect 16313 21301 16347 21335
rect 16405 21301 16439 21335
rect 16681 21301 16715 21335
rect 17049 21301 17083 21335
rect 19533 21301 19567 21335
rect 23029 21301 23063 21335
rect 25145 21301 25179 21335
rect 25421 21301 25455 21335
rect 5825 21097 5859 21131
rect 8677 21097 8711 21131
rect 13645 21097 13679 21131
rect 16681 21097 16715 21131
rect 17877 21097 17911 21131
rect 22845 21097 22879 21131
rect 6285 21029 6319 21063
rect 9965 21029 9999 21063
rect 12909 21029 12943 21063
rect 15485 21029 15519 21063
rect 18889 21029 18923 21063
rect 21189 21029 21223 21063
rect 23949 21029 23983 21063
rect 24041 21029 24075 21063
rect 2881 20961 2915 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 10425 20961 10459 20995
rect 10517 20961 10551 20995
rect 11161 20961 11195 20995
rect 11437 20961 11471 20995
rect 16037 20961 16071 20995
rect 17233 20961 17267 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 22201 20961 22235 20995
rect 23305 20961 23339 20995
rect 23397 20961 23431 20995
rect 25145 20961 25179 20995
rect 2237 20893 2271 20927
rect 4077 20893 4111 20927
rect 6469 20893 6503 20927
rect 7113 20893 7147 20927
rect 10333 20893 10367 20927
rect 14381 20893 14415 20927
rect 15945 20893 15979 20927
rect 18245 20893 18279 20927
rect 19441 20893 19475 20927
rect 22017 20893 22051 20927
rect 22109 20893 22143 20927
rect 23213 20893 23247 20927
rect 25053 20893 25087 20927
rect 8953 20825 8987 20859
rect 9321 20825 9355 20859
rect 13553 20825 13587 20859
rect 17049 20825 17083 20859
rect 24409 20825 24443 20859
rect 24961 20825 24995 20859
rect 5733 20757 5767 20791
rect 14473 20757 14507 20791
rect 14841 20757 14875 20791
rect 15025 20757 15059 20791
rect 15853 20757 15887 20791
rect 17141 20757 17175 20791
rect 21649 20757 21683 20791
rect 24593 20757 24627 20791
rect 6469 20553 6503 20587
rect 7757 20553 7791 20587
rect 12081 20553 12115 20587
rect 12449 20553 12483 20587
rect 13185 20553 13219 20587
rect 18705 20553 18739 20587
rect 21005 20553 21039 20587
rect 22109 20553 22143 20587
rect 22569 20553 22603 20587
rect 1685 20485 1719 20519
rect 2145 20485 2179 20519
rect 4905 20485 4939 20519
rect 5089 20485 5123 20519
rect 5181 20485 5215 20519
rect 11805 20485 11839 20519
rect 12541 20485 12575 20519
rect 23765 20485 23799 20519
rect 3065 20417 3099 20451
rect 6009 20417 6043 20451
rect 7297 20417 7331 20451
rect 8585 20417 8619 20451
rect 9045 20417 9079 20451
rect 13553 20417 13587 20451
rect 15853 20417 15887 20451
rect 16957 20417 16991 20451
rect 22477 20417 22511 20451
rect 23489 20417 23523 20451
rect 3341 20349 3375 20383
rect 6653 20349 6687 20383
rect 9321 20349 9355 20383
rect 12725 20349 12759 20383
rect 13829 20349 13863 20383
rect 17233 20349 17267 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 22661 20349 22695 20383
rect 1869 20281 1903 20315
rect 5825 20281 5859 20315
rect 6837 20281 6871 20315
rect 15301 20281 15335 20315
rect 21465 20281 21499 20315
rect 23121 20281 23155 20315
rect 7113 20213 7147 20247
rect 8401 20213 8435 20247
rect 10793 20213 10827 20247
rect 11161 20213 11195 20247
rect 11345 20213 11379 20247
rect 11621 20213 11655 20247
rect 15945 20213 15979 20247
rect 16405 20213 16439 20247
rect 21281 20213 21315 20247
rect 25237 20213 25271 20247
rect 10425 20009 10459 20043
rect 14933 20009 14967 20043
rect 17693 20009 17727 20043
rect 21360 20009 21394 20043
rect 4537 19941 4571 19975
rect 13369 19941 13403 19975
rect 18889 19941 18923 19975
rect 20637 19941 20671 19975
rect 2513 19873 2547 19907
rect 5181 19873 5215 19907
rect 5457 19873 5491 19907
rect 7389 19873 7423 19907
rect 10977 19873 11011 19907
rect 15485 19873 15519 19907
rect 17233 19873 17267 19907
rect 18153 19873 18187 19907
rect 18245 19873 18279 19907
rect 18705 19873 18739 19907
rect 20085 19873 20119 19907
rect 21097 19873 21131 19907
rect 23949 19873 23983 19907
rect 25053 19873 25087 19907
rect 25145 19873 25179 19907
rect 2237 19805 2271 19839
rect 4721 19805 4755 19839
rect 6653 19805 6687 19839
rect 7113 19805 7147 19839
rect 11621 19805 11655 19839
rect 14289 19805 14323 19839
rect 18061 19805 18095 19839
rect 19809 19805 19843 19839
rect 23673 19805 23707 19839
rect 8401 19737 8435 19771
rect 10793 19737 10827 19771
rect 10885 19737 10919 19771
rect 11897 19737 11931 19771
rect 15393 19737 15427 19771
rect 16185 19737 16219 19771
rect 17049 19737 17083 19771
rect 20453 19737 20487 19771
rect 6469 19669 6503 19703
rect 9137 19669 9171 19703
rect 9781 19669 9815 19703
rect 13645 19669 13679 19703
rect 13921 19669 13955 19703
rect 15301 19669 15335 19703
rect 16313 19669 16347 19703
rect 19441 19669 19475 19703
rect 19901 19669 19935 19703
rect 22845 19669 22879 19703
rect 23305 19669 23339 19703
rect 23765 19669 23799 19703
rect 24593 19669 24627 19703
rect 24961 19669 24995 19703
rect 3893 19465 3927 19499
rect 5825 19465 5859 19499
rect 7113 19465 7147 19499
rect 8401 19465 8435 19499
rect 11069 19465 11103 19499
rect 11529 19465 11563 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 18797 19465 18831 19499
rect 19625 19465 19659 19499
rect 20453 19465 20487 19499
rect 20913 19465 20947 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 25053 19465 25087 19499
rect 15393 19397 15427 19431
rect 19717 19397 19751 19431
rect 20821 19397 20855 19431
rect 1961 19329 1995 19363
rect 4077 19329 4111 19363
rect 4813 19329 4847 19363
rect 6009 19329 6043 19363
rect 7297 19329 7331 19363
rect 7941 19329 7975 19363
rect 8585 19329 8619 19363
rect 9045 19329 9079 19363
rect 12725 19329 12759 19363
rect 16313 19329 16347 19363
rect 17038 19329 17072 19363
rect 23305 19329 23339 19363
rect 2237 19261 2271 19295
rect 4537 19261 4571 19295
rect 6469 19261 6503 19295
rect 6653 19261 6687 19295
rect 6745 19261 6779 19295
rect 9321 19261 9355 19295
rect 12081 19261 12115 19295
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 17325 19261 17359 19295
rect 19901 19261 19935 19295
rect 21005 19261 21039 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 23581 19261 23615 19295
rect 7757 19193 7791 19227
rect 16681 19193 16715 19227
rect 19257 19193 19291 19227
rect 21465 19193 21499 19227
rect 25329 19193 25363 19227
rect 10793 19125 10827 19159
rect 11345 19125 11379 19159
rect 11805 19125 11839 19159
rect 16129 19125 16163 19159
rect 1961 18921 1995 18955
rect 3893 18921 3927 18955
rect 8401 18921 8435 18955
rect 12541 18921 12575 18955
rect 14289 18921 14323 18955
rect 2605 18853 2639 18887
rect 9229 18853 9263 18887
rect 13001 18853 13035 18887
rect 17233 18853 17267 18887
rect 18061 18853 18095 18887
rect 22569 18853 22603 18887
rect 4077 18785 4111 18819
rect 5825 18785 5859 18819
rect 7113 18785 7147 18819
rect 7389 18785 7423 18819
rect 9781 18785 9815 18819
rect 13645 18785 13679 18819
rect 14841 18785 14875 18819
rect 18613 18785 18647 18819
rect 20637 18785 20671 18819
rect 23121 18785 23155 18819
rect 25053 18785 25087 18819
rect 25237 18785 25271 18819
rect 2145 18717 2179 18751
rect 2789 18717 2823 18751
rect 3433 18717 3467 18751
rect 4169 18717 4203 18751
rect 4721 18717 4755 18751
rect 5365 18717 5399 18751
rect 6101 18717 6135 18751
rect 8585 18717 8619 18751
rect 9597 18717 9631 18751
rect 10425 18717 10459 18751
rect 15485 18717 15519 18751
rect 18429 18717 18463 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 23029 18717 23063 18751
rect 23857 18717 23891 18751
rect 9689 18649 9723 18683
rect 13369 18649 13403 18683
rect 14657 18649 14691 18683
rect 15761 18649 15795 18683
rect 24041 18649 24075 18683
rect 3249 18581 3283 18615
rect 4537 18581 4571 18615
rect 5181 18581 5215 18615
rect 11713 18581 11747 18615
rect 12725 18581 12759 18615
rect 13461 18581 13495 18615
rect 14749 18581 14783 18615
rect 17509 18581 17543 18615
rect 17693 18581 17727 18615
rect 18521 18581 18555 18615
rect 19441 18581 19475 18615
rect 19901 18581 19935 18615
rect 22109 18581 22143 18615
rect 22937 18581 22971 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 2237 18377 2271 18411
rect 2605 18377 2639 18411
rect 3249 18377 3283 18411
rect 4537 18377 4571 18411
rect 5825 18377 5859 18411
rect 7665 18377 7699 18411
rect 8309 18377 8343 18411
rect 12173 18377 12207 18411
rect 14289 18377 14323 18411
rect 15209 18377 15243 18411
rect 15669 18377 15703 18411
rect 16313 18377 16347 18411
rect 19625 18377 19659 18411
rect 23305 18377 23339 18411
rect 24225 18377 24259 18411
rect 9229 18309 9263 18343
rect 11253 18309 11287 18343
rect 13001 18309 13035 18343
rect 22017 18309 22051 18343
rect 24041 18309 24075 18343
rect 24501 18309 24535 18343
rect 24961 18309 24995 18343
rect 1777 18241 1811 18275
rect 2145 18241 2179 18275
rect 2789 18241 2823 18275
rect 3433 18241 3467 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 6009 18241 6043 18275
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 15577 18241 15611 18275
rect 16405 18241 16439 18275
rect 17233 18241 17267 18275
rect 18429 18241 18463 18275
rect 20821 18241 20855 18275
rect 3801 18173 3835 18207
rect 3893 18173 3927 18207
rect 6561 18173 6595 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 15761 18173 15795 18207
rect 17325 18173 17359 18207
rect 17417 18173 17451 18207
rect 18521 18173 18555 18207
rect 18705 18173 18739 18207
rect 19717 18173 19751 18207
rect 19809 18173 19843 18207
rect 20913 18173 20947 18207
rect 21005 18173 21039 18207
rect 25053 18173 25087 18207
rect 25237 18173 25271 18207
rect 1593 18105 1627 18139
rect 5181 18105 5215 18139
rect 7021 18105 7055 18139
rect 10701 18105 10735 18139
rect 11805 18105 11839 18139
rect 16865 18105 16899 18139
rect 20453 18105 20487 18139
rect 21465 18105 21499 18139
rect 24593 18105 24627 18139
rect 6745 18037 6779 18071
rect 11161 18037 11195 18071
rect 18061 18037 18095 18071
rect 19257 18037 19291 18071
rect 2789 17833 2823 17867
rect 6469 17833 6503 17867
rect 7113 17833 7147 17867
rect 7757 17833 7791 17867
rect 17141 17833 17175 17867
rect 18245 17833 18279 17867
rect 20992 17833 21026 17867
rect 22477 17833 22511 17867
rect 24593 17833 24627 17867
rect 1593 17765 1627 17799
rect 16681 17765 16715 17799
rect 23305 17765 23339 17799
rect 2237 17697 2271 17731
rect 5181 17697 5215 17731
rect 5457 17697 5491 17731
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14289 17697 14323 17731
rect 14933 17697 14967 17731
rect 17693 17697 17727 17731
rect 19901 17697 19935 17731
rect 20085 17697 20119 17731
rect 20729 17697 20763 17731
rect 23949 17697 23983 17731
rect 25053 17697 25087 17731
rect 25237 17697 25271 17731
rect 1777 17629 1811 17663
rect 3433 17629 3467 17663
rect 4261 17629 4295 17663
rect 4721 17629 4755 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 9781 17629 9815 17663
rect 18797 17629 18831 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 10057 17561 10091 17595
rect 15209 17561 15243 17595
rect 17509 17561 17543 17595
rect 19809 17561 19843 17595
rect 3249 17493 3283 17527
rect 3893 17493 3927 17527
rect 4537 17493 4571 17527
rect 8401 17493 8435 17527
rect 9137 17493 9171 17527
rect 11529 17493 11563 17527
rect 13737 17493 13771 17527
rect 17601 17493 17635 17527
rect 18613 17493 18647 17527
rect 19441 17493 19475 17527
rect 22845 17493 22879 17527
rect 23029 17493 23063 17527
rect 24961 17493 24995 17527
rect 5825 17289 5859 17323
rect 15853 17289 15887 17323
rect 15945 17289 15979 17323
rect 24317 17289 24351 17323
rect 9505 17221 9539 17255
rect 11345 17221 11379 17255
rect 11989 17221 12023 17255
rect 21465 17221 21499 17255
rect 4077 17153 4111 17187
rect 4813 17153 4847 17187
rect 6009 17153 6043 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 11713 17153 11747 17187
rect 14381 17153 14415 17187
rect 15025 17153 15059 17187
rect 17233 17153 17267 17187
rect 17325 17153 17359 17187
rect 18337 17153 18371 17187
rect 20821 17153 20855 17187
rect 22569 17153 22603 17187
rect 24869 17153 24903 17187
rect 4537 17085 4571 17119
rect 10977 17085 11011 17119
rect 13461 17085 13495 17119
rect 13921 17085 13955 17119
rect 16037 17085 16071 17119
rect 17417 17085 17451 17119
rect 17877 17085 17911 17119
rect 18613 17085 18647 17119
rect 20085 17085 20119 17119
rect 20453 17085 20487 17119
rect 22845 17085 22879 17119
rect 3893 17017 3927 17051
rect 7849 17017 7883 17051
rect 8585 17017 8619 17051
rect 14841 17017 14875 17051
rect 25053 17017 25087 17051
rect 6561 16949 6595 16983
rect 7205 16949 7239 16983
rect 15485 16949 15519 16983
rect 16865 16949 16899 16983
rect 21833 16949 21867 16983
rect 22017 16949 22051 16983
rect 22293 16949 22327 16983
rect 25329 16949 25363 16983
rect 4261 16745 4295 16779
rect 8401 16745 8435 16779
rect 9045 16745 9079 16779
rect 16037 16745 16071 16779
rect 19704 16745 19738 16779
rect 25237 16745 25271 16779
rect 6929 16677 6963 16711
rect 7297 16609 7331 16643
rect 7481 16609 7515 16643
rect 9229 16609 9263 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 14289 16609 14323 16643
rect 17141 16609 17175 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 7941 16541 7975 16575
rect 8585 16541 8619 16575
rect 9689 16541 9723 16575
rect 11161 16541 11195 16575
rect 11989 16541 12023 16575
rect 16681 16541 16715 16575
rect 21649 16541 21683 16575
rect 24593 16541 24627 16575
rect 5365 16473 5399 16507
rect 12265 16473 12299 16507
rect 14565 16473 14599 16507
rect 4721 16405 4755 16439
rect 7757 16405 7791 16439
rect 9505 16405 9539 16439
rect 10149 16405 10183 16439
rect 10793 16405 10827 16439
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18889 16405 18923 16439
rect 21189 16405 21223 16439
rect 24041 16405 24075 16439
rect 8033 16201 8067 16235
rect 9781 16201 9815 16235
rect 10793 16201 10827 16235
rect 13461 16201 13495 16235
rect 15025 16201 15059 16235
rect 16681 16201 16715 16235
rect 18429 16201 18463 16235
rect 19349 16201 19383 16235
rect 20545 16201 20579 16235
rect 20913 16201 20947 16235
rect 22477 16201 22511 16235
rect 23857 16201 23891 16235
rect 25237 16201 25271 16235
rect 14381 16133 14415 16167
rect 8217 16065 8251 16099
rect 8677 16065 8711 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 14289 16065 14323 16099
rect 15209 16065 15243 16099
rect 15853 16065 15887 16099
rect 17141 16065 17175 16099
rect 19717 16065 19751 16099
rect 21005 16065 21039 16099
rect 22385 16065 22419 16099
rect 23765 16065 23799 16099
rect 24593 16065 24627 16099
rect 10885 15997 10919 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 14565 15997 14599 16031
rect 15945 15997 15979 16031
rect 16037 15997 16071 16031
rect 19809 15997 19843 16031
rect 19901 15997 19935 16031
rect 21189 15997 21223 16031
rect 22569 15997 22603 16031
rect 23949 15997 23983 16031
rect 10425 15929 10459 15963
rect 15485 15929 15519 15963
rect 23029 15929 23063 15963
rect 8493 15861 8527 15895
rect 9137 15861 9171 15895
rect 13921 15861 13955 15895
rect 21557 15861 21591 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 8769 15657 8803 15691
rect 9873 15657 9907 15691
rect 13829 15657 13863 15691
rect 16037 15657 16071 15691
rect 16681 15657 16715 15691
rect 18705 15657 18739 15691
rect 22845 15657 22879 15691
rect 24133 15657 24167 15691
rect 25329 15657 25363 15691
rect 9229 15589 9263 15623
rect 10793 15521 10827 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 20085 15521 20119 15555
rect 21189 15521 21223 15555
rect 21281 15521 21315 15555
rect 25145 15521 25179 15555
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10517 15453 10551 15487
rect 13093 15453 13127 15487
rect 21097 15453 21131 15487
rect 23397 15453 23431 15487
rect 24685 15453 24719 15487
rect 13185 15385 13219 15419
rect 14565 15385 14599 15419
rect 19901 15385 19935 15419
rect 22017 15385 22051 15419
rect 22753 15385 22787 15419
rect 23857 15385 23891 15419
rect 24869 15385 24903 15419
rect 12265 15317 12299 15351
rect 12725 15317 12759 15351
rect 16313 15317 16347 15351
rect 19073 15317 19107 15351
rect 19533 15317 19567 15351
rect 19993 15317 20027 15351
rect 20729 15317 20763 15351
rect 22109 15317 22143 15351
rect 9413 15113 9447 15147
rect 9689 15113 9723 15147
rect 13921 15113 13955 15147
rect 16129 15113 16163 15147
rect 18981 15113 19015 15147
rect 21373 15113 21407 15147
rect 24593 15113 24627 15147
rect 9873 15045 9907 15079
rect 22109 15045 22143 15079
rect 23121 15045 23155 15079
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 22845 14977 22879 15011
rect 25145 14977 25179 15011
rect 10057 14909 10091 14943
rect 11713 14909 11747 14943
rect 11989 14909 12023 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 16865 14909 16899 14943
rect 17141 14909 17175 14943
rect 19349 14909 19383 14943
rect 19625 14909 19659 14943
rect 21097 14909 21131 14943
rect 10333 14841 10367 14875
rect 25329 14841 25363 14875
rect 10977 14773 11011 14807
rect 13461 14773 13495 14807
rect 14841 14773 14875 14807
rect 18613 14773 18647 14807
rect 21557 14773 21591 14807
rect 22201 14773 22235 14807
rect 10425 14569 10459 14603
rect 12449 14569 12483 14603
rect 25329 14569 25363 14603
rect 18245 14501 18279 14535
rect 19441 14501 19475 14535
rect 23305 14501 23339 14535
rect 25237 14501 25271 14535
rect 10977 14433 11011 14467
rect 13553 14433 13587 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16773 14433 16807 14467
rect 19993 14433 20027 14467
rect 22385 14433 22419 14467
rect 22937 14433 22971 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 10701 14365 10735 14399
rect 13093 14365 13127 14399
rect 16497 14365 16531 14399
rect 19901 14365 19935 14399
rect 20821 14365 20855 14399
rect 24685 14365 24719 14399
rect 18705 14297 18739 14331
rect 19809 14297 19843 14331
rect 24869 14297 24903 14331
rect 12909 14229 12943 14263
rect 16037 14229 16071 14263
rect 20545 14229 20579 14263
rect 23673 14229 23707 14263
rect 11161 14025 11195 14059
rect 11805 14025 11839 14059
rect 12449 14025 12483 14059
rect 13093 14025 13127 14059
rect 15485 14025 15519 14059
rect 16129 14025 16163 14059
rect 17049 14025 17083 14059
rect 17509 14025 17543 14059
rect 21189 14025 21223 14059
rect 18245 13957 18279 13991
rect 21097 13957 21131 13991
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 13277 13889 13311 13923
rect 13737 13889 13771 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 22109 13889 22143 13923
rect 22845 13889 22879 13923
rect 25145 13889 25179 13923
rect 11345 13821 11379 13855
rect 17601 13821 17635 13855
rect 21281 13821 21315 13855
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 25329 13821 25363 13855
rect 22293 13753 22327 13787
rect 14000 13685 14034 13719
rect 15853 13685 15887 13719
rect 16681 13685 16715 13719
rect 19717 13685 19751 13719
rect 20361 13685 20395 13719
rect 20729 13685 20763 13719
rect 16037 13481 16071 13515
rect 18705 13481 18739 13515
rect 19980 13481 20014 13515
rect 21465 13481 21499 13515
rect 23949 13481 23983 13515
rect 13553 13413 13587 13447
rect 19349 13413 19383 13447
rect 24133 13413 24167 13447
rect 12081 13345 12115 13379
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 16773 13345 16807 13379
rect 21925 13345 21959 13379
rect 23673 13345 23707 13379
rect 25053 13345 25087 13379
rect 25145 13345 25179 13379
rect 11805 13277 11839 13311
rect 18889 13277 18923 13311
rect 19717 13277 19751 13311
rect 9597 13209 9631 13243
rect 14565 13209 14599 13243
rect 22201 13209 22235 13243
rect 24961 13209 24995 13243
rect 10885 13141 10919 13175
rect 13921 13141 13955 13175
rect 18245 13141 18279 13175
rect 24593 13141 24627 13175
rect 11529 12937 11563 12971
rect 12633 12937 12667 12971
rect 14289 12937 14323 12971
rect 19533 12937 19567 12971
rect 20729 12937 20763 12971
rect 21373 12937 21407 12971
rect 23765 12937 23799 12971
rect 13001 12869 13035 12903
rect 24225 12869 24259 12903
rect 25329 12869 25363 12903
rect 16865 12801 16899 12835
rect 19441 12801 19475 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 25053 12801 25087 12835
rect 15209 12733 15243 12767
rect 15485 12733 15519 12767
rect 17141 12733 17175 12767
rect 19625 12733 19659 12767
rect 20821 12733 20855 12767
rect 22293 12733 22327 12767
rect 18613 12665 18647 12699
rect 16405 12597 16439 12631
rect 19073 12597 19107 12631
rect 20269 12597 20303 12631
rect 21465 12597 21499 12631
rect 24869 12597 24903 12631
rect 13921 12393 13955 12427
rect 15485 12393 15519 12427
rect 17509 12393 17543 12427
rect 24041 12393 24075 12427
rect 24501 12393 24535 12427
rect 24685 12393 24719 12427
rect 14565 12257 14599 12291
rect 15761 12257 15795 12291
rect 17969 12257 18003 12291
rect 19441 12257 19475 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 25053 12257 25087 12291
rect 14289 12189 14323 12223
rect 21833 12189 21867 12223
rect 16037 12121 16071 12155
rect 18669 12121 18703 12155
rect 18889 12121 18923 12155
rect 19717 12121 19751 12155
rect 13461 12053 13495 12087
rect 13737 12053 13771 12087
rect 21189 12053 21223 12087
rect 21649 12053 21683 12087
rect 14565 11849 14599 11883
rect 16129 11849 16163 11883
rect 16773 11849 16807 11883
rect 18889 11849 18923 11883
rect 21189 11849 21223 11883
rect 13093 11781 13127 11815
rect 23305 11781 23339 11815
rect 12817 11713 12851 11747
rect 15301 11713 15335 11747
rect 15853 11713 15887 11747
rect 16313 11713 16347 11747
rect 17141 11713 17175 11747
rect 19441 11713 19475 11747
rect 22109 11713 22143 11747
rect 23949 11713 23983 11747
rect 15669 11645 15703 11679
rect 17417 11645 17451 11679
rect 19717 11645 19751 11679
rect 24777 11645 24811 11679
rect 15117 11509 15151 11543
rect 21465 11509 21499 11543
rect 15485 11305 15519 11339
rect 16129 11305 16163 11339
rect 16773 11305 16807 11339
rect 17417 11305 17451 11339
rect 21005 11305 21039 11339
rect 25329 11305 25363 11339
rect 14749 11237 14783 11271
rect 20453 11237 20487 11271
rect 24593 11237 24627 11271
rect 25145 11237 25179 11271
rect 18061 11169 18095 11203
rect 21649 11169 21683 11203
rect 22201 11169 22235 11203
rect 23857 11169 23891 11203
rect 15669 11101 15703 11135
rect 16313 11101 16347 11135
rect 16957 11101 16991 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 19349 11101 19383 11135
rect 19533 11101 19567 11135
rect 19993 11101 20027 11135
rect 21189 11101 21223 11135
rect 22661 11101 22695 11135
rect 24777 11101 24811 11135
rect 20177 11033 20211 11067
rect 25421 11033 25455 11067
rect 18705 10965 18739 10999
rect 20729 10965 20763 10999
rect 22293 10965 22327 10999
rect 15761 10761 15795 10795
rect 16405 10761 16439 10795
rect 17141 10761 17175 10795
rect 18061 10761 18095 10795
rect 23305 10693 23339 10727
rect 16957 10625 16991 10659
rect 18245 10625 18279 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 20177 10649 20211 10683
rect 20821 10625 20855 10659
rect 21465 10625 21499 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 17417 10557 17451 10591
rect 24685 10557 24719 10591
rect 18705 10489 18739 10523
rect 19993 10489 20027 10523
rect 19349 10421 19383 10455
rect 20637 10421 20671 10455
rect 21281 10421 21315 10455
rect 17417 10217 17451 10251
rect 24593 10217 24627 10251
rect 20729 10149 20763 10183
rect 23121 10149 23155 10183
rect 18061 10081 18095 10115
rect 21373 10081 21407 10115
rect 23581 10081 23615 10115
rect 25145 10081 25179 10115
rect 17601 10013 17635 10047
rect 18337 10013 18371 10047
rect 19625 10013 19659 10047
rect 20913 10013 20947 10047
rect 24041 10013 24075 10047
rect 25053 10013 25087 10047
rect 20085 9945 20119 9979
rect 21649 9945 21683 9979
rect 24961 9945 24995 9979
rect 19441 9877 19475 9911
rect 23857 9877 23891 9911
rect 21281 9673 21315 9707
rect 23305 9605 23339 9639
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19533 9537 19567 9571
rect 20177 9537 20211 9571
rect 20913 9537 20947 9571
rect 21465 9537 21499 9571
rect 21649 9537 21683 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 24777 9469 24811 9503
rect 18061 9401 18095 9435
rect 19349 9401 19383 9435
rect 20729 9401 20763 9435
rect 18705 9333 18739 9367
rect 19993 9333 20027 9367
rect 11805 9129 11839 9163
rect 20913 9129 20947 9163
rect 25145 9129 25179 9163
rect 25421 9129 25455 9163
rect 21281 9061 21315 9095
rect 10057 8993 10091 9027
rect 19441 8993 19475 9027
rect 22017 8993 22051 9027
rect 23857 8993 23891 9027
rect 19073 8925 19107 8959
rect 19717 8925 19751 8959
rect 20545 8925 20579 8959
rect 21465 8925 21499 8959
rect 22661 8925 22695 8959
rect 10333 8857 10367 8891
rect 12081 8857 12115 8891
rect 24685 8857 24719 8891
rect 24869 8857 24903 8891
rect 19441 8585 19475 8619
rect 21373 8585 21407 8619
rect 23305 8517 23339 8551
rect 19625 8449 19659 8483
rect 20269 8449 20303 8483
rect 20913 8449 20947 8483
rect 21281 8449 21315 8483
rect 22109 8449 22143 8483
rect 23949 8449 23983 8483
rect 24593 8381 24627 8415
rect 20085 8313 20119 8347
rect 20729 8313 20763 8347
rect 22017 8041 22051 8075
rect 21373 7973 21407 8007
rect 23857 7905 23891 7939
rect 20913 7837 20947 7871
rect 21557 7837 21591 7871
rect 22201 7837 22235 7871
rect 22845 7837 22879 7871
rect 24869 7837 24903 7871
rect 20085 7769 20119 7803
rect 20729 7701 20763 7735
rect 24685 7701 24719 7735
rect 21281 7497 21315 7531
rect 23305 7429 23339 7463
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 24685 7293 24719 7327
rect 20637 7225 20671 7259
rect 22017 6817 22051 6851
rect 23857 6817 23891 6851
rect 20821 6749 20855 6783
rect 21465 6749 21499 6783
rect 22661 6749 22695 6783
rect 24685 6749 24719 6783
rect 24869 6681 24903 6715
rect 20637 6613 20671 6647
rect 21281 6613 21315 6647
rect 9321 6409 9355 6443
rect 21557 6409 21591 6443
rect 23305 6341 23339 6375
rect 8677 6273 8711 6307
rect 22293 6273 22327 6307
rect 24133 6273 24167 6307
rect 24777 6205 24811 6239
rect 22017 5865 22051 5899
rect 21373 5797 21407 5831
rect 21557 5661 21591 5695
rect 22201 5661 22235 5695
rect 22845 5661 22879 5695
rect 24869 5661 24903 5695
rect 23857 5593 23891 5627
rect 24685 5525 24719 5559
rect 23305 5253 23339 5287
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 24685 5117 24719 5151
rect 22017 4777 22051 4811
rect 21741 4573 21775 4607
rect 22201 4573 22235 4607
rect 22661 4573 22695 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 24685 4437 24719 4471
rect 20085 4097 20119 4131
rect 22293 4097 22327 4131
rect 23949 4097 23983 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 6837 3485 6871 3519
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 24777 3485 24811 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 7481 3349 7515 3383
rect 24593 3349 24627 3383
rect 7481 3145 7515 3179
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 6837 3009 6871 3043
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 24133 3009 24167 3043
rect 19441 2941 19475 2975
rect 21281 2941 21315 2975
rect 6561 2805 6595 2839
rect 6561 2601 6595 2635
rect 19809 2601 19843 2635
rect 7849 2465 7883 2499
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 20269 2397 20303 2431
rect 22845 2397 22879 2431
rect 21281 2329 21315 2363
rect 23857 2329 23891 2363
<< metal1 >>
rect 3050 26392 3056 26444
rect 3108 26432 3114 26444
rect 3326 26432 3332 26444
rect 3108 26404 3332 26432
rect 3108 26392 3114 26404
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 2498 26188 2504 26240
rect 2556 26228 2562 26240
rect 12618 26228 12624 26240
rect 2556 26200 12624 26228
rect 2556 26188 2562 26200
rect 12618 26188 12624 26200
rect 12676 26188 12682 26240
rect 9122 25032 9128 25084
rect 9180 25072 9186 25084
rect 20898 25072 20904 25084
rect 9180 25044 20904 25072
rect 9180 25032 9186 25044
rect 20898 25032 20904 25044
rect 20956 25032 20962 25084
rect 4798 24964 4804 25016
rect 4856 25004 4862 25016
rect 18690 25004 18696 25016
rect 4856 24976 18696 25004
rect 4856 24964 4862 24976
rect 18690 24964 18696 24976
rect 18748 24964 18754 25016
rect 10226 24896 10232 24948
rect 10284 24936 10290 24948
rect 22370 24936 22376 24948
rect 10284 24908 22376 24936
rect 10284 24896 10290 24908
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 7742 24828 7748 24880
rect 7800 24868 7806 24880
rect 18414 24868 18420 24880
rect 7800 24840 18420 24868
rect 7800 24828 7806 24840
rect 18414 24828 18420 24840
rect 18472 24828 18478 24880
rect 20530 24828 20536 24880
rect 20588 24868 20594 24880
rect 23382 24868 23388 24880
rect 20588 24840 23388 24868
rect 20588 24828 20594 24840
rect 23382 24828 23388 24840
rect 23440 24828 23446 24880
rect 2406 24760 2412 24812
rect 2464 24800 2470 24812
rect 15194 24800 15200 24812
rect 2464 24772 15200 24800
rect 2464 24760 2470 24772
rect 15194 24760 15200 24772
rect 15252 24800 15258 24812
rect 17402 24800 17408 24812
rect 15252 24772 17408 24800
rect 15252 24760 15258 24772
rect 17402 24760 17408 24772
rect 17460 24760 17466 24812
rect 17770 24760 17776 24812
rect 17828 24800 17834 24812
rect 24118 24800 24124 24812
rect 17828 24772 24124 24800
rect 17828 24760 17834 24772
rect 24118 24760 24124 24772
rect 24176 24760 24182 24812
rect 5810 24692 5816 24744
rect 5868 24732 5874 24744
rect 7282 24732 7288 24744
rect 5868 24704 7288 24732
rect 5868 24692 5874 24704
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 10410 24692 10416 24744
rect 10468 24732 10474 24744
rect 19242 24732 19248 24744
rect 10468 24704 19248 24732
rect 10468 24692 10474 24704
rect 19242 24692 19248 24704
rect 19300 24692 19306 24744
rect 2314 24624 2320 24676
rect 2372 24664 2378 24676
rect 7098 24664 7104 24676
rect 2372 24636 7104 24664
rect 2372 24624 2378 24636
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 14826 24624 14832 24676
rect 14884 24664 14890 24676
rect 22830 24664 22836 24676
rect 14884 24636 22836 24664
rect 14884 24624 14890 24636
rect 22830 24624 22836 24636
rect 22888 24624 22894 24676
rect 5902 24556 5908 24608
rect 5960 24596 5966 24608
rect 10318 24596 10324 24608
rect 5960 24568 10324 24596
rect 5960 24556 5966 24568
rect 10318 24556 10324 24568
rect 10376 24556 10382 24608
rect 11698 24556 11704 24608
rect 11756 24596 11762 24608
rect 14550 24596 14556 24608
rect 11756 24568 14556 24596
rect 11756 24556 11762 24568
rect 14550 24556 14556 24568
rect 14608 24556 14614 24608
rect 22646 24556 22652 24608
rect 22704 24596 22710 24608
rect 23106 24596 23112 24608
rect 22704 24568 23112 24596
rect 22704 24556 22710 24568
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 3970 24352 3976 24404
rect 4028 24352 4034 24404
rect 6730 24352 6736 24404
rect 6788 24392 6794 24404
rect 6788 24364 8524 24392
rect 6788 24352 6794 24364
rect 8496 24324 8524 24364
rect 9122 24352 9128 24404
rect 9180 24352 9186 24404
rect 17310 24392 17316 24404
rect 11348 24364 17316 24392
rect 11054 24324 11060 24336
rect 8496 24296 11060 24324
rect 11054 24284 11060 24296
rect 11112 24284 11118 24336
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11238 24256 11244 24268
rect 11011 24228 11244 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3878 24188 3884 24200
rect 2271 24160 3884 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 6730 24148 6736 24200
rect 6788 24148 6794 24200
rect 7282 24148 7288 24200
rect 7340 24148 7346 24200
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 9416 24160 9781 24188
rect 1578 24080 1584 24132
rect 1636 24080 1642 24132
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8662 24120 8668 24132
rect 5859 24092 8668 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 1765 24055 1823 24061
rect 1765 24021 1777 24055
rect 1811 24052 1823 24055
rect 2314 24052 2320 24064
rect 1811 24024 2320 24052
rect 1811 24021 1823 24024
rect 1765 24015 1823 24021
rect 2314 24012 2320 24024
rect 2372 24012 2378 24064
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 6549 24055 6607 24061
rect 6549 24052 6561 24055
rect 6420 24024 6561 24052
rect 6420 24012 6426 24024
rect 6549 24021 6561 24024
rect 6595 24021 6607 24055
rect 6549 24015 6607 24021
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 9416 24052 9444 24160
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 11348 24188 11376 24364
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 21269 24395 21327 24401
rect 21269 24392 21281 24395
rect 17420 24364 21281 24392
rect 12342 24284 12348 24336
rect 12400 24324 12406 24336
rect 17420 24324 17448 24364
rect 21269 24361 21281 24364
rect 21315 24361 21327 24395
rect 21269 24355 21327 24361
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 22152 24364 23612 24392
rect 22152 24352 22158 24364
rect 12400 24296 12664 24324
rect 12400 24284 12406 24296
rect 12434 24256 12440 24268
rect 12406 24216 12440 24256
rect 12492 24216 12498 24268
rect 12636 24256 12664 24296
rect 17236 24296 17448 24324
rect 18708 24296 22094 24324
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12636 24228 12817 24256
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 14461 24259 14519 24265
rect 14461 24225 14473 24259
rect 14507 24256 14519 24259
rect 17236 24256 17264 24296
rect 14507 24228 17264 24256
rect 17313 24259 17371 24265
rect 14507 24225 14519 24228
rect 14461 24219 14519 24225
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 17402 24256 17408 24268
rect 17359 24228 17408 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 17494 24216 17500 24268
rect 17552 24216 17558 24268
rect 18506 24216 18512 24268
rect 18564 24216 18570 24268
rect 18708 24265 18736 24296
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24225 18751 24259
rect 18693 24219 18751 24225
rect 20073 24259 20131 24265
rect 20073 24225 20085 24259
rect 20119 24256 20131 24259
rect 20714 24256 20720 24268
rect 20119 24228 20720 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 20714 24216 20720 24228
rect 20772 24216 20778 24268
rect 22066 24256 22094 24296
rect 22554 24256 22560 24268
rect 22066 24228 22560 24256
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 23584 24256 23612 24364
rect 23584 24228 23796 24256
rect 10008 24160 11376 24188
rect 11885 24191 11943 24197
rect 10008 24148 10014 24160
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12406 24188 12434 24216
rect 11931 24160 12434 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12526 24148 12532 24200
rect 12584 24148 12590 24200
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14185 24191 14243 24197
rect 14185 24188 14197 24191
rect 14056 24160 14197 24188
rect 14056 24148 14062 24160
rect 14185 24157 14197 24160
rect 14231 24188 14243 24191
rect 14737 24191 14795 24197
rect 14231 24160 14320 24188
rect 14231 24157 14243 24160
rect 14185 24151 14243 24157
rect 9582 24080 9588 24132
rect 9640 24120 9646 24132
rect 14292 24120 14320 24160
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 15838 24188 15844 24200
rect 14783 24160 15844 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 15979 24160 19472 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 9640 24092 12434 24120
rect 9640 24080 9646 24092
rect 7524 24024 9444 24052
rect 7524 24012 7530 24024
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 11701 24055 11759 24061
rect 11701 24052 11713 24055
rect 9916 24024 11713 24052
rect 9916 24012 9922 24024
rect 11701 24021 11713 24024
rect 11747 24021 11759 24055
rect 12406 24052 12434 24092
rect 12544 24092 14228 24120
rect 14292 24092 16436 24120
rect 12544 24052 12572 24092
rect 12406 24024 12572 24052
rect 14200 24052 14228 24092
rect 16408 24064 16436 24092
rect 17586 24080 17592 24132
rect 17644 24120 17650 24132
rect 18230 24120 18236 24132
rect 17644 24092 18236 24120
rect 17644 24080 17650 24092
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 18417 24123 18475 24129
rect 18417 24089 18429 24123
rect 18463 24120 18475 24123
rect 19150 24120 19156 24132
rect 18463 24092 19156 24120
rect 18463 24089 18475 24092
rect 18417 24083 18475 24089
rect 19150 24080 19156 24092
rect 19208 24080 19214 24132
rect 15749 24055 15807 24061
rect 15749 24052 15761 24055
rect 14200 24024 15761 24052
rect 11701 24015 11759 24021
rect 15749 24021 15761 24024
rect 15795 24021 15807 24055
rect 15749 24015 15807 24021
rect 16206 24012 16212 24064
rect 16264 24012 16270 24064
rect 16390 24012 16396 24064
rect 16448 24012 16454 24064
rect 16850 24012 16856 24064
rect 16908 24012 16914 24064
rect 17218 24012 17224 24064
rect 17276 24012 17282 24064
rect 18049 24055 18107 24061
rect 18049 24021 18061 24055
rect 18095 24052 18107 24055
rect 18966 24052 18972 24064
rect 18095 24024 18972 24052
rect 18095 24021 18107 24024
rect 18049 24015 18107 24021
rect 18966 24012 18972 24024
rect 19024 24012 19030 24064
rect 19334 24012 19340 24064
rect 19392 24012 19398 24064
rect 19444 24061 19472 24160
rect 21450 24148 21456 24200
rect 21508 24148 21514 24200
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 23768 24188 23796 24228
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 25133 24259 25191 24265
rect 25133 24256 25145 24259
rect 23900 24228 25145 24256
rect 23900 24216 23906 24228
rect 25133 24225 25145 24228
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 23768 24160 24961 24188
rect 24949 24157 24961 24160
rect 24995 24157 25007 24191
rect 24949 24151 25007 24157
rect 25038 24148 25044 24200
rect 25096 24148 25102 24200
rect 19889 24123 19947 24129
rect 19889 24089 19901 24123
rect 19935 24120 19947 24123
rect 22462 24120 22468 24132
rect 19935 24092 22468 24120
rect 19935 24089 19947 24092
rect 19889 24083 19947 24089
rect 22462 24080 22468 24092
rect 22520 24080 22526 24132
rect 22557 24123 22615 24129
rect 22557 24089 22569 24123
rect 22603 24120 22615 24123
rect 23934 24120 23940 24132
rect 22603 24092 22968 24120
rect 23782 24092 23940 24120
rect 22603 24089 22615 24092
rect 22557 24083 22615 24089
rect 22940 24064 22968 24092
rect 23934 24080 23940 24092
rect 23992 24080 23998 24132
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 19797 24055 19855 24061
rect 19797 24052 19809 24055
rect 19576 24024 19809 24052
rect 19576 24012 19582 24024
rect 19797 24021 19809 24024
rect 19843 24021 19855 24055
rect 19797 24015 19855 24021
rect 20622 24012 20628 24064
rect 20680 24012 20686 24064
rect 21913 24055 21971 24061
rect 21913 24021 21925 24055
rect 21959 24052 21971 24055
rect 22002 24052 22008 24064
rect 21959 24024 22008 24052
rect 21959 24021 21971 24024
rect 21913 24015 21971 24021
rect 22002 24012 22008 24024
rect 22060 24012 22066 24064
rect 22922 24012 22928 24064
rect 22980 24012 22986 24064
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24118 24052 24124 24064
rect 24075 24024 24124 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 24854 24052 24860 24064
rect 24627 24024 24860 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 2501 23851 2559 23857
rect 2501 23817 2513 23851
rect 2547 23848 2559 23851
rect 6822 23848 6828 23860
rect 2547 23820 6828 23848
rect 2547 23817 2559 23820
rect 2501 23811 2559 23817
rect 6822 23808 6828 23820
rect 6880 23808 6886 23860
rect 8018 23848 8024 23860
rect 6932 23820 8024 23848
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5350 23780 5356 23792
rect 4019 23752 5356 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 5810 23740 5816 23792
rect 5868 23740 5874 23792
rect 6932 23780 6960 23820
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 9306 23808 9312 23860
rect 9364 23848 9370 23860
rect 11609 23851 11667 23857
rect 11609 23848 11621 23851
rect 9364 23820 11621 23848
rect 9364 23808 9370 23820
rect 11609 23817 11621 23820
rect 11655 23848 11667 23851
rect 11698 23848 11704 23860
rect 11655 23820 11704 23848
rect 11655 23817 11667 23820
rect 11609 23811 11667 23817
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 11793 23851 11851 23857
rect 11793 23817 11805 23851
rect 11839 23848 11851 23851
rect 13817 23851 13875 23857
rect 13817 23848 13829 23851
rect 11839 23820 13829 23848
rect 11839 23817 11851 23820
rect 11793 23811 11851 23817
rect 13817 23817 13829 23820
rect 13863 23848 13875 23851
rect 13998 23848 14004 23860
rect 13863 23820 14004 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23817 14151 23851
rect 14093 23811 14151 23817
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 20622 23848 20628 23860
rect 14507 23820 20628 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 9125 23783 9183 23789
rect 6564 23752 6960 23780
rect 7024 23752 8064 23780
rect 1670 23672 1676 23724
rect 1728 23672 1734 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3602 23712 3608 23724
rect 3007 23684 3608 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3602 23672 3608 23684
rect 3660 23672 3666 23724
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 6564 23712 6592 23752
rect 4847 23684 6592 23712
rect 6641 23715 6699 23721
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 6641 23681 6653 23715
rect 6687 23712 6699 23715
rect 6730 23712 6736 23724
rect 6687 23684 6736 23712
rect 6687 23681 6699 23684
rect 6641 23675 6699 23681
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 6914 23672 6920 23724
rect 6972 23672 6978 23724
rect 5994 23604 6000 23656
rect 6052 23644 6058 23656
rect 7024 23644 7052 23752
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 8036 23712 8064 23752
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 10134 23780 10140 23792
rect 9171 23752 10140 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 10962 23740 10968 23792
rect 11020 23780 11026 23792
rect 14108 23780 14136 23811
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 22922 23808 22928 23860
rect 22980 23848 22986 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 22980 23820 24041 23848
rect 22980 23808 22986 23820
rect 24029 23817 24041 23820
rect 24075 23848 24087 23851
rect 25498 23848 25504 23860
rect 24075 23820 25504 23848
rect 24075 23817 24087 23820
rect 24029 23811 24087 23817
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 11020 23752 14136 23780
rect 11020 23740 11026 23752
rect 15194 23740 15200 23792
rect 15252 23740 15258 23792
rect 15378 23740 15384 23792
rect 15436 23780 15442 23792
rect 15933 23783 15991 23789
rect 15933 23780 15945 23783
rect 15436 23752 15945 23780
rect 15436 23740 15442 23752
rect 15933 23749 15945 23752
rect 15979 23749 15991 23783
rect 15933 23743 15991 23749
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23780 16083 23783
rect 16114 23780 16120 23792
rect 16071 23752 16120 23780
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 16114 23740 16120 23752
rect 16172 23740 16178 23792
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23780 17279 23783
rect 17402 23780 17408 23792
rect 17267 23752 17408 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 17402 23740 17408 23752
rect 17460 23740 17466 23792
rect 18414 23780 18420 23792
rect 18064 23752 18420 23780
rect 9766 23712 9772 23724
rect 8036 23684 9772 23712
rect 7929 23675 7987 23681
rect 6052 23616 7052 23644
rect 6052 23604 6058 23616
rect 1857 23579 1915 23585
rect 1857 23545 1869 23579
rect 1903 23576 1915 23579
rect 5902 23576 5908 23588
rect 1903 23548 5908 23576
rect 1903 23545 1915 23548
rect 1857 23539 1915 23545
rect 5902 23536 5908 23548
rect 5960 23536 5966 23588
rect 5442 23468 5448 23520
rect 5500 23508 5506 23520
rect 7944 23508 7972 23675
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 8018 23604 8024 23656
rect 8076 23644 8082 23656
rect 9968 23644 9996 23675
rect 12066 23672 12072 23724
rect 12124 23672 12130 23724
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 15896 23684 17264 23712
rect 15896 23672 15902 23684
rect 10042 23644 10048 23656
rect 8076 23616 9904 23644
rect 9968 23616 10048 23644
rect 8076 23604 8082 23616
rect 9876 23576 9904 23616
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 12710 23576 12716 23588
rect 9876 23548 12716 23576
rect 12710 23536 12716 23548
rect 12768 23536 12774 23588
rect 14568 23576 14596 23607
rect 14734 23604 14740 23656
rect 14792 23604 14798 23656
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16298 23644 16304 23656
rect 16255 23616 16304 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16298 23604 16304 23616
rect 16356 23604 16362 23656
rect 17236 23644 17264 23684
rect 17310 23672 17316 23724
rect 17368 23672 17374 23724
rect 18064 23712 18092 23752
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 18874 23740 18880 23792
rect 18932 23740 18938 23792
rect 23934 23780 23940 23792
rect 23782 23752 23940 23780
rect 23934 23740 23940 23752
rect 23992 23780 23998 23792
rect 24305 23783 24363 23789
rect 24305 23780 24317 23783
rect 23992 23752 24317 23780
rect 23992 23740 23998 23752
rect 24305 23749 24317 23752
rect 24351 23749 24363 23783
rect 24305 23743 24363 23749
rect 25130 23740 25136 23792
rect 25188 23740 25194 23792
rect 20714 23712 20720 23724
rect 17420 23684 18092 23712
rect 19812 23684 20720 23712
rect 17420 23644 17448 23684
rect 17236 23616 17448 23644
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23644 17555 23647
rect 17770 23644 17776 23656
rect 17543 23616 17776 23644
rect 17543 23613 17555 23616
rect 17497 23607 17555 23613
rect 17770 23604 17776 23616
rect 17828 23604 17834 23656
rect 18046 23604 18052 23656
rect 18104 23604 18110 23656
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23644 18383 23647
rect 19812 23644 19840 23684
rect 20714 23672 20720 23684
rect 20772 23672 20778 23724
rect 18371 23616 19840 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20036 23616 20269 23644
rect 20036 23604 20042 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 20622 23604 20628 23656
rect 20680 23604 20686 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 22094 23644 22100 23656
rect 20947 23616 22100 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 17954 23576 17960 23588
rect 14568 23548 17960 23576
rect 17954 23536 17960 23548
rect 18012 23536 18018 23588
rect 20916 23576 20944 23607
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 22554 23604 22560 23656
rect 22612 23644 22618 23656
rect 23290 23644 23296 23656
rect 22612 23616 23296 23644
rect 22612 23604 22618 23616
rect 23290 23604 23296 23616
rect 23348 23604 23354 23656
rect 24302 23604 24308 23656
rect 24360 23644 24366 23656
rect 24673 23647 24731 23653
rect 24673 23644 24685 23647
rect 24360 23616 24685 23644
rect 24360 23604 24366 23616
rect 24673 23613 24685 23616
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 19720 23548 20944 23576
rect 5500 23480 7972 23508
rect 5500 23468 5506 23480
rect 9214 23468 9220 23520
rect 9272 23508 9278 23520
rect 10962 23508 10968 23520
rect 9272 23480 10968 23508
rect 9272 23468 9278 23480
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 12618 23468 12624 23520
rect 12676 23508 12682 23520
rect 13354 23508 13360 23520
rect 12676 23480 13360 23508
rect 12676 23468 12682 23480
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 15565 23511 15623 23517
rect 15565 23477 15577 23511
rect 15611 23508 15623 23511
rect 16666 23508 16672 23520
rect 15611 23480 16672 23508
rect 15611 23477 15623 23480
rect 15565 23471 15623 23477
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 17218 23468 17224 23520
rect 17276 23508 17282 23520
rect 19720 23508 19748 23548
rect 17276 23480 19748 23508
rect 17276 23468 17282 23480
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 20070 23468 20076 23520
rect 20128 23468 20134 23520
rect 21358 23468 21364 23520
rect 21416 23508 21422 23520
rect 21821 23511 21879 23517
rect 21821 23508 21833 23511
rect 21416 23480 21833 23508
rect 21416 23468 21422 23480
rect 21821 23477 21833 23480
rect 21867 23477 21879 23511
rect 22112 23508 22140 23604
rect 24581 23579 24639 23585
rect 24581 23545 24593 23579
rect 24627 23576 24639 23579
rect 25866 23576 25872 23588
rect 24627 23548 25872 23576
rect 24627 23545 24639 23548
rect 24581 23539 24639 23545
rect 25866 23536 25872 23548
rect 25924 23536 25930 23588
rect 22370 23508 22376 23520
rect 22112 23480 22376 23508
rect 21821 23471 21879 23477
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 22554 23468 22560 23520
rect 22612 23508 22618 23520
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 22612 23480 25237 23508
rect 22612 23468 22618 23480
rect 25225 23477 25237 23480
rect 25271 23477 25283 23511
rect 25225 23471 25283 23477
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 3602 23304 3608 23316
rect 1627 23276 3608 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 3602 23264 3608 23276
rect 3660 23304 3666 23316
rect 3970 23304 3976 23316
rect 3660 23276 3976 23304
rect 3660 23264 3666 23276
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 6730 23264 6736 23316
rect 6788 23304 6794 23316
rect 9122 23304 9128 23316
rect 6788 23276 9128 23304
rect 6788 23264 6794 23276
rect 9122 23264 9128 23276
rect 9180 23304 9186 23316
rect 13262 23304 13268 23316
rect 9180 23276 13268 23304
rect 9180 23264 9186 23276
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 15654 23304 15660 23316
rect 14016 23276 15660 23304
rect 1765 23239 1823 23245
rect 1765 23205 1777 23239
rect 1811 23236 1823 23239
rect 1946 23236 1952 23248
rect 1811 23208 1952 23236
rect 1811 23205 1823 23208
rect 1765 23199 1823 23205
rect 1946 23196 1952 23208
rect 2004 23196 2010 23248
rect 7006 23236 7012 23248
rect 2746 23208 7012 23236
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2746 23100 2774 23208
rect 7006 23196 7012 23208
rect 7064 23196 7070 23248
rect 9398 23236 9404 23248
rect 8220 23208 9404 23236
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 4614 23168 4620 23180
rect 3283 23140 4620 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23168 6607 23171
rect 7650 23168 7656 23180
rect 6595 23140 7656 23168
rect 6595 23137 6607 23140
rect 6549 23131 6607 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 8220 23177 8248 23208
rect 9398 23196 9404 23208
rect 9456 23196 9462 23248
rect 14016 23236 14044 23276
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16850 23264 16856 23316
rect 16908 23304 16914 23316
rect 16908 23276 25084 23304
rect 16908 23264 16914 23276
rect 9508 23208 14044 23236
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23137 8263 23171
rect 8205 23131 8263 23137
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 9508 23168 9536 23208
rect 16298 23196 16304 23248
rect 16356 23236 16362 23248
rect 17034 23236 17040 23248
rect 16356 23208 17040 23236
rect 16356 23196 16362 23208
rect 17034 23196 17040 23208
rect 17092 23236 17098 23248
rect 19426 23236 19432 23248
rect 17092 23208 19432 23236
rect 17092 23196 17098 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 23382 23196 23388 23248
rect 23440 23196 23446 23248
rect 8720 23140 9536 23168
rect 8720 23128 8726 23140
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11664 23140 12173 23168
rect 11664 23128 11670 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 12161 23131 12219 23137
rect 12250 23128 12256 23180
rect 12308 23168 12314 23180
rect 14918 23168 14924 23180
rect 12308 23140 14924 23168
rect 12308 23128 12314 23140
rect 14918 23128 14924 23140
rect 14976 23128 14982 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 15335 23140 17785 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 17773 23137 17785 23140
rect 17819 23168 17831 23171
rect 18506 23168 18512 23180
rect 17819 23140 18512 23168
rect 17819 23137 17831 23140
rect 17773 23131 17831 23137
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 18690 23128 18696 23180
rect 18748 23128 18754 23180
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 21174 23168 21180 23180
rect 19751 23140 21180 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 22278 23168 22284 23180
rect 21683 23140 22284 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22278 23128 22284 23140
rect 22336 23168 22342 23180
rect 23290 23168 23296 23180
rect 22336 23140 23296 23168
rect 22336 23128 22342 23140
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 25056 23177 25084 23276
rect 25041 23171 25099 23177
rect 25041 23137 25053 23171
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 2271 23072 2774 23100
rect 4065 23103 4123 23109
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 4065 23069 4077 23103
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 4080 23032 4108 23063
rect 4338 23060 4344 23112
rect 4396 23060 4402 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 5534 23100 5540 23112
rect 5491 23072 5540 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 6270 23060 6276 23112
rect 6328 23100 6334 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6328 23072 7205 23100
rect 6328 23060 6334 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23100 9459 23103
rect 9582 23100 9588 23112
rect 9447 23072 9588 23100
rect 9447 23069 9459 23072
rect 9401 23063 9459 23069
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23069 9919 23103
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 9861 23063 9919 23069
rect 9968 23072 11713 23100
rect 5810 23032 5816 23044
rect 4080 23004 5816 23032
rect 5810 22992 5816 23004
rect 5868 22992 5874 23044
rect 7558 22992 7564 23044
rect 7616 23032 7622 23044
rect 9876 23032 9904 23063
rect 7616 23004 9904 23032
rect 7616 22992 7622 23004
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 9968 22964 9996 23072
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 11701 23063 11759 23069
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14240 23072 15025 23100
rect 14240 23060 14246 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 16390 23060 16396 23112
rect 16448 23060 16454 23112
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 17589 23103 17647 23109
rect 17589 23100 17601 23103
rect 16724 23072 17601 23100
rect 16724 23060 16730 23072
rect 17589 23069 17601 23072
rect 17635 23069 17647 23103
rect 17862 23100 17868 23112
rect 17589 23063 17647 23069
rect 17696 23072 17868 23100
rect 10042 22992 10048 23044
rect 10100 23032 10106 23044
rect 13906 23032 13912 23044
rect 10100 23004 13912 23032
rect 10100 22992 10106 23004
rect 13906 22992 13912 23004
rect 13964 22992 13970 23044
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 14056 23004 14381 23032
rect 14056 22992 14062 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 14550 22992 14556 23044
rect 14608 23032 14614 23044
rect 15378 23032 15384 23044
rect 14608 23004 15384 23032
rect 14608 22992 14614 23004
rect 15378 22992 15384 23004
rect 15436 22992 15442 23044
rect 17696 23041 17724 23072
rect 17862 23060 17868 23072
rect 17920 23060 17926 23112
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 19334 23100 19340 23112
rect 18104 23072 19340 23100
rect 18104 23060 18110 23072
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 24762 23060 24768 23112
rect 24820 23100 24826 23112
rect 25148 23100 25176 23131
rect 24820 23072 25176 23100
rect 24820 23060 24826 23072
rect 17681 23035 17739 23041
rect 16776 23004 17356 23032
rect 9263 22936 9996 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 12526 22924 12532 22976
rect 12584 22964 12590 22976
rect 12802 22964 12808 22976
rect 12584 22936 12808 22964
rect 12584 22924 12590 22936
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 13538 22924 13544 22976
rect 13596 22924 13602 22976
rect 14458 22924 14464 22976
rect 14516 22924 14522 22976
rect 15654 22924 15660 22976
rect 15712 22964 15718 22976
rect 16298 22964 16304 22976
rect 15712 22936 16304 22964
rect 15712 22924 15718 22936
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 16574 22924 16580 22976
rect 16632 22964 16638 22976
rect 16776 22973 16804 23004
rect 16761 22967 16819 22973
rect 16761 22964 16773 22967
rect 16632 22936 16773 22964
rect 16632 22924 16638 22936
rect 16761 22933 16773 22936
rect 16807 22933 16819 22967
rect 16761 22927 16819 22933
rect 17218 22924 17224 22976
rect 17276 22924 17282 22976
rect 17328 22964 17356 23004
rect 17681 23001 17693 23035
rect 17727 23001 17739 23035
rect 17681 22995 17739 23001
rect 18509 23035 18567 23041
rect 18509 23001 18521 23035
rect 18555 23032 18567 23035
rect 18782 23032 18788 23044
rect 18555 23004 18788 23032
rect 18555 23001 18567 23004
rect 18509 22995 18567 23001
rect 18782 22992 18788 23004
rect 18840 23032 18846 23044
rect 19978 23032 19984 23044
rect 18840 23004 19984 23032
rect 18840 22992 18846 23004
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 20162 22992 20168 23044
rect 20220 22992 20226 23044
rect 21910 22992 21916 23044
rect 21968 22992 21974 23044
rect 22066 23004 22402 23032
rect 17770 22964 17776 22976
rect 17328 22936 17776 22964
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 18690 22924 18696 22976
rect 18748 22964 18754 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18748 22936 18981 22964
rect 18748 22924 18754 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 20714 22924 20720 22976
rect 20772 22964 20778 22976
rect 21177 22967 21235 22973
rect 21177 22964 21189 22967
rect 20772 22936 21189 22964
rect 20772 22924 20778 22936
rect 21177 22933 21189 22936
rect 21223 22933 21235 22967
rect 21177 22927 21235 22933
rect 21818 22924 21824 22976
rect 21876 22964 21882 22976
rect 22066 22964 22094 23004
rect 23750 22992 23756 23044
rect 23808 23032 23814 23044
rect 25314 23032 25320 23044
rect 23808 23004 25320 23032
rect 23808 22992 23814 23004
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 21876 22936 22094 22964
rect 21876 22924 21882 22936
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 23845 22967 23903 22973
rect 23845 22964 23857 22967
rect 23624 22936 23857 22964
rect 23624 22924 23630 22936
rect 23845 22933 23857 22936
rect 23891 22933 23903 22967
rect 23845 22927 23903 22933
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 24946 22924 24952 22976
rect 25004 22924 25010 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1486 22720 1492 22772
rect 1544 22760 1550 22772
rect 1673 22763 1731 22769
rect 1673 22760 1685 22763
rect 1544 22732 1685 22760
rect 1544 22720 1550 22732
rect 1673 22729 1685 22732
rect 1719 22760 1731 22763
rect 1719 22732 2176 22760
rect 1719 22729 1731 22732
rect 1673 22723 1731 22729
rect 2148 22701 2176 22732
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7098 22760 7104 22772
rect 6972 22732 7104 22760
rect 6972 22720 6978 22732
rect 7098 22720 7104 22732
rect 7156 22760 7162 22772
rect 7193 22763 7251 22769
rect 7193 22760 7205 22763
rect 7156 22732 7205 22760
rect 7156 22720 7162 22732
rect 7193 22729 7205 22732
rect 7239 22729 7251 22763
rect 12250 22760 12256 22772
rect 7193 22723 7251 22729
rect 8496 22732 12256 22760
rect 2133 22695 2191 22701
rect 2133 22661 2145 22695
rect 2179 22661 2191 22695
rect 2133 22655 2191 22661
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 8386 22692 8392 22704
rect 6687 22664 8392 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 8386 22652 8392 22664
rect 8444 22652 8450 22704
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 4522 22624 4528 22636
rect 3007 22596 4528 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 4522 22584 4528 22596
rect 4580 22584 4586 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22624 4859 22627
rect 5626 22624 5632 22636
rect 4847 22596 5632 22624
rect 4847 22593 4859 22596
rect 4801 22587 4859 22593
rect 5626 22584 5632 22596
rect 5684 22584 5690 22636
rect 6730 22584 6736 22636
rect 6788 22624 6794 22636
rect 6825 22627 6883 22633
rect 6825 22624 6837 22627
rect 6788 22596 6837 22624
rect 6788 22584 6794 22596
rect 6825 22593 6837 22596
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 1581 22559 1639 22565
rect 1581 22525 1593 22559
rect 1627 22556 1639 22559
rect 1627 22528 2774 22556
rect 1627 22525 1639 22528
rect 1581 22519 1639 22525
rect 2746 22488 2774 22528
rect 3602 22516 3608 22568
rect 3660 22556 3666 22568
rect 7576 22556 7604 22587
rect 3660 22528 7604 22556
rect 3660 22516 3666 22528
rect 4154 22488 4160 22500
rect 2746 22460 4160 22488
rect 4154 22448 4160 22460
rect 4212 22488 4218 22500
rect 8496 22488 8524 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12768 22732 13093 22760
rect 12768 22720 12774 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 14550 22760 14556 22772
rect 13320 22732 14556 22760
rect 13320 22720 13326 22732
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15381 22763 15439 22769
rect 15381 22760 15393 22763
rect 14792 22732 15393 22760
rect 14792 22720 14798 22732
rect 15381 22729 15393 22732
rect 15427 22729 15439 22763
rect 16482 22760 16488 22772
rect 15381 22723 15439 22729
rect 15856 22732 16488 22760
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 11146 22652 11152 22704
rect 11204 22692 11210 22704
rect 12161 22695 12219 22701
rect 11204 22664 12112 22692
rect 11204 22652 11210 22664
rect 10778 22584 10784 22636
rect 10836 22584 10842 22636
rect 12084 22633 12112 22664
rect 12161 22661 12173 22695
rect 12207 22692 12219 22695
rect 14182 22692 14188 22704
rect 12207 22664 13584 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 12069 22627 12127 22633
rect 10888 22596 11192 22624
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 10888 22556 10916 22596
rect 9723 22528 10916 22556
rect 11164 22556 11192 22596
rect 12069 22593 12081 22627
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12986 22584 12992 22636
rect 13044 22584 13050 22636
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 11164 22528 12265 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 12253 22525 12265 22528
rect 12299 22556 12311 22559
rect 12434 22556 12440 22568
rect 12299 22528 12440 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12434 22516 12440 22528
rect 12492 22516 12498 22568
rect 4212 22460 8524 22488
rect 4212 22448 4218 22460
rect 10870 22448 10876 22500
rect 10928 22488 10934 22500
rect 11149 22491 11207 22497
rect 11149 22488 11161 22491
rect 10928 22460 11161 22488
rect 10928 22448 10934 22460
rect 11149 22457 11161 22460
rect 11195 22488 11207 22491
rect 13354 22488 13360 22500
rect 11195 22460 13360 22488
rect 11195 22457 11207 22460
rect 11149 22451 11207 22457
rect 13354 22448 13360 22460
rect 13412 22448 13418 22500
rect 2222 22380 2228 22432
rect 2280 22380 2286 22432
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 10042 22420 10048 22432
rect 5868 22392 10048 22420
rect 5868 22380 5874 22392
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11296 22392 11713 22420
rect 11296 22380 11302 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 12250 22380 12256 22432
rect 12308 22420 12314 22432
rect 12986 22420 12992 22432
rect 12308 22392 12992 22420
rect 12308 22380 12314 22392
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 13556 22420 13584 22664
rect 13648 22664 14188 22692
rect 13648 22633 13676 22664
rect 14182 22652 14188 22664
rect 14240 22652 14246 22704
rect 15286 22652 15292 22704
rect 15344 22692 15350 22704
rect 15856 22692 15884 22732
rect 16482 22720 16488 22732
rect 16540 22720 16546 22772
rect 17862 22760 17868 22772
rect 16960 22732 17868 22760
rect 15344 22664 15884 22692
rect 15933 22695 15991 22701
rect 15344 22652 15350 22664
rect 15933 22661 15945 22695
rect 15979 22692 15991 22695
rect 16022 22692 16028 22704
rect 15979 22664 16028 22692
rect 15979 22661 15991 22664
rect 15933 22655 15991 22661
rect 16022 22652 16028 22664
rect 16080 22692 16086 22704
rect 16206 22692 16212 22704
rect 16080 22664 16212 22692
rect 16080 22652 16086 22664
rect 16206 22652 16212 22664
rect 16264 22652 16270 22704
rect 16960 22692 16988 22732
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 18564 22732 18613 22760
rect 18564 22720 18570 22732
rect 18601 22729 18613 22732
rect 18647 22729 18659 22763
rect 18601 22723 18659 22729
rect 19242 22720 19248 22772
rect 19300 22720 19306 22772
rect 23750 22760 23756 22772
rect 22112 22732 23756 22760
rect 16868 22664 16988 22692
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 15562 22624 15568 22636
rect 15042 22596 15568 22624
rect 13633 22587 13691 22593
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 16574 22624 16580 22636
rect 15672 22596 16580 22624
rect 13909 22559 13967 22565
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 15672 22556 15700 22596
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 16868 22633 16896 22664
rect 17034 22652 17040 22704
rect 17092 22692 17098 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 17092 22664 17141 22692
rect 17092 22652 17098 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 18414 22652 18420 22704
rect 18472 22692 18478 22704
rect 18472 22664 20116 22692
rect 18472 22652 18478 22664
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 18874 22624 18880 22636
rect 18262 22596 18880 22624
rect 16853 22587 16911 22593
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 20088 22633 20116 22664
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 13955 22528 15700 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 15746 22516 15752 22568
rect 15804 22556 15810 22568
rect 19168 22556 19196 22587
rect 20622 22584 20628 22636
rect 20680 22624 20686 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 20680 22596 22017 22624
rect 20680 22584 20686 22596
rect 22005 22593 22017 22596
rect 22051 22624 22063 22627
rect 22112 22624 22140 22732
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 23934 22720 23940 22772
rect 23992 22720 23998 22772
rect 23952 22692 23980 22720
rect 22051 22596 22140 22624
rect 22204 22664 24058 22692
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 15804 22528 19196 22556
rect 15804 22516 15810 22528
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 20533 22559 20591 22565
rect 20533 22556 20545 22559
rect 20220 22528 20545 22556
rect 20220 22516 20226 22528
rect 20533 22525 20545 22528
rect 20579 22556 20591 22559
rect 21082 22556 21088 22568
rect 20579 22528 21088 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 21082 22516 21088 22528
rect 21140 22556 21146 22568
rect 21818 22556 21824 22568
rect 21140 22528 21824 22556
rect 21140 22516 21146 22528
rect 21818 22516 21824 22528
rect 21876 22556 21882 22568
rect 22204 22556 22232 22664
rect 21876 22528 22232 22556
rect 22281 22559 22339 22565
rect 21876 22516 21882 22528
rect 22281 22525 22293 22559
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 15194 22448 15200 22500
rect 15252 22488 15258 22500
rect 16117 22491 16175 22497
rect 16117 22488 16129 22491
rect 15252 22460 16129 22488
rect 15252 22448 15258 22460
rect 16117 22457 16129 22460
rect 16163 22457 16175 22491
rect 16117 22451 16175 22457
rect 16390 22448 16396 22500
rect 16448 22488 16454 22500
rect 16485 22491 16543 22497
rect 16485 22488 16497 22491
rect 16448 22460 16497 22488
rect 16448 22448 16454 22460
rect 16485 22457 16497 22460
rect 16531 22488 16543 22491
rect 16850 22488 16856 22500
rect 16531 22460 16856 22488
rect 16531 22457 16543 22460
rect 16485 22451 16543 22457
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 20990 22488 20996 22500
rect 18156 22460 20996 22488
rect 16298 22420 16304 22432
rect 13556 22392 16304 22420
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 17678 22420 17684 22432
rect 16724 22392 17684 22420
rect 16724 22380 16730 22392
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18156 22420 18184 22460
rect 20990 22448 20996 22460
rect 21048 22448 21054 22500
rect 22094 22448 22100 22500
rect 22152 22488 22158 22500
rect 22296 22488 22324 22519
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 23569 22559 23627 22565
rect 23569 22525 23581 22559
rect 23615 22556 23627 22559
rect 24118 22556 24124 22568
rect 23615 22528 24124 22556
rect 23615 22525 23627 22528
rect 23569 22519 23627 22525
rect 24118 22516 24124 22528
rect 24176 22556 24182 22568
rect 25774 22556 25780 22568
rect 24176 22528 25780 22556
rect 24176 22516 24182 22528
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 22152 22460 22324 22488
rect 22152 22448 22158 22460
rect 17828 22392 18184 22420
rect 17828 22380 17834 22392
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 18932 22392 19625 22420
rect 18932 22380 18938 22392
rect 19613 22389 19625 22392
rect 19659 22420 19671 22423
rect 20070 22420 20076 22432
rect 19659 22392 20076 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20254 22380 20260 22432
rect 20312 22420 20318 22432
rect 22646 22420 22652 22432
rect 20312 22392 22652 22420
rect 20312 22380 20318 22392
rect 22646 22380 22652 22392
rect 22704 22380 22710 22432
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24762 22420 24768 22432
rect 23716 22392 24768 22420
rect 23716 22380 23722 22392
rect 24762 22380 24768 22392
rect 24820 22420 24826 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24820 22392 25053 22420
rect 24820 22380 24826 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 25041 22383 25099 22389
rect 25409 22423 25467 22429
rect 25409 22389 25421 22423
rect 25455 22420 25467 22423
rect 25682 22420 25688 22432
rect 25455 22392 25688 22420
rect 25455 22389 25467 22392
rect 25409 22383 25467 22389
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 2280 22188 8432 22216
rect 2280 22176 2286 22188
rect 8294 22148 8300 22160
rect 8220 22120 8300 22148
rect 1670 22040 1676 22092
rect 1728 22040 1734 22092
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8113 22083 8171 22089
rect 8113 22049 8125 22083
rect 8159 22080 8171 22083
rect 8220 22080 8248 22120
rect 8294 22108 8300 22120
rect 8352 22108 8358 22160
rect 8404 22148 8432 22188
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 13446 22216 13452 22228
rect 9548 22188 13452 22216
rect 9548 22176 9554 22188
rect 13446 22176 13452 22188
rect 13504 22176 13510 22228
rect 14540 22219 14598 22225
rect 14540 22185 14552 22219
rect 14586 22216 14598 22219
rect 14734 22216 14740 22228
rect 14586 22188 14740 22216
rect 14586 22185 14598 22188
rect 14540 22179 14598 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 18785 22219 18843 22225
rect 15580 22188 16988 22216
rect 10594 22148 10600 22160
rect 8404 22120 10600 22148
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 12768 22120 14412 22148
rect 12768 22108 12774 22120
rect 8159 22052 8248 22080
rect 8159 22049 8171 22052
rect 8113 22043 8171 22049
rect 9030 22040 9036 22092
rect 9088 22080 9094 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 9088 22052 10701 22080
rect 9088 22040 9094 22052
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 11054 22080 11060 22092
rect 10735 22052 11060 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 12434 22040 12440 22092
rect 12492 22040 12498 22092
rect 14384 22080 14412 22120
rect 15580 22080 15608 22188
rect 16298 22108 16304 22160
rect 16356 22148 16362 22160
rect 16485 22151 16543 22157
rect 16485 22148 16497 22151
rect 16356 22120 16497 22148
rect 16356 22108 16362 22120
rect 16485 22117 16497 22120
rect 16531 22117 16543 22151
rect 16485 22111 16543 22117
rect 16960 22094 16988 22188
rect 18785 22185 18797 22219
rect 18831 22216 18843 22219
rect 18874 22216 18880 22228
rect 18831 22188 18880 22216
rect 18831 22185 18843 22188
rect 18785 22179 18843 22185
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 19613 22219 19671 22225
rect 19613 22216 19625 22219
rect 19484 22188 19625 22216
rect 19484 22176 19490 22188
rect 19613 22185 19625 22188
rect 19659 22185 19671 22219
rect 19613 22179 19671 22185
rect 20612 22219 20670 22225
rect 20612 22185 20624 22219
rect 20658 22216 20670 22219
rect 21266 22216 21272 22228
rect 20658 22188 21272 22216
rect 20658 22185 20670 22188
rect 20612 22179 20670 22185
rect 21266 22176 21272 22188
rect 21324 22216 21330 22228
rect 23842 22216 23848 22228
rect 21324 22188 23848 22216
rect 21324 22176 21330 22188
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 17678 22108 17684 22160
rect 17736 22148 17742 22160
rect 18969 22151 19027 22157
rect 18969 22148 18981 22151
rect 17736 22120 18981 22148
rect 17736 22108 17742 22120
rect 18969 22117 18981 22120
rect 19015 22117 19027 22151
rect 18969 22111 19027 22117
rect 22370 22108 22376 22160
rect 22428 22148 22434 22160
rect 22646 22148 22652 22160
rect 22428 22120 22652 22148
rect 22428 22108 22434 22120
rect 22646 22108 22652 22120
rect 22704 22108 22710 22160
rect 25406 22148 25412 22160
rect 25240 22120 25412 22148
rect 16390 22080 16396 22092
rect 14384 22052 15608 22080
rect 15672 22052 16396 22080
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2682 22012 2688 22024
rect 2271 21984 2688 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4430 22012 4436 22024
rect 4295 21984 4436 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 4430 21972 4436 21984
rect 4488 21972 4494 22024
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 22012 5595 22015
rect 6454 22012 6460 22024
rect 5583 21984 6460 22012
rect 5583 21981 5595 21984
rect 5537 21975 5595 21981
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 8941 22015 8999 22021
rect 8941 21981 8953 22015
rect 8987 22012 8999 22015
rect 9490 22012 9496 22024
rect 8987 21984 9496 22012
rect 8987 21981 8999 21984
rect 8941 21975 8999 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 12066 21972 12072 22024
rect 12124 22012 12130 22024
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12124 21984 13093 22012
rect 12124 21972 12130 21984
rect 13081 21981 13093 21984
rect 13127 22012 13139 22015
rect 13446 22012 13452 22024
rect 13127 21984 13452 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 13446 21972 13452 21984
rect 13504 21972 13510 22024
rect 14182 21972 14188 22024
rect 14240 22012 14246 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14240 21984 14289 22012
rect 14240 21972 14246 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 15672 22012 15700 22052
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 16960 22089 17080 22094
rect 16960 22083 17095 22089
rect 16960 22066 17049 22083
rect 17037 22049 17049 22066
rect 17083 22080 17095 22083
rect 17083 22052 17117 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 18138 22080 18144 22092
rect 17276 22052 18144 22080
rect 17276 22040 17282 22052
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 18233 22043 18291 22049
rect 18248 22012 18276 22043
rect 18414 22040 18420 22092
rect 18472 22080 18478 22092
rect 23474 22089 23480 22092
rect 22557 22083 22615 22089
rect 22557 22080 22569 22083
rect 18472 22052 22569 22080
rect 18472 22040 18478 22052
rect 22557 22049 22569 22052
rect 22603 22049 22615 22083
rect 23431 22083 23480 22089
rect 23431 22080 23443 22083
rect 22557 22043 22615 22049
rect 22940 22052 23443 22080
rect 15620 21998 15700 22012
rect 15620 21984 15686 21998
rect 16040 21984 18276 22012
rect 15620 21972 15626 21984
rect 9398 21904 9404 21956
rect 9456 21944 9462 21956
rect 10410 21944 10416 21956
rect 9456 21916 10416 21944
rect 9456 21904 9462 21916
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 10965 21947 11023 21953
rect 10965 21913 10977 21947
rect 11011 21913 11023 21947
rect 10965 21907 11023 21913
rect 12897 21947 12955 21953
rect 12897 21913 12909 21947
rect 12943 21944 12955 21947
rect 13538 21944 13544 21956
rect 12943 21916 13544 21944
rect 12943 21913 12955 21916
rect 12897 21907 12955 21913
rect 2130 21836 2136 21888
rect 2188 21876 2194 21888
rect 8202 21876 8208 21888
rect 2188 21848 8208 21876
rect 2188 21836 2194 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 10502 21876 10508 21888
rect 10091 21848 10508 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10980 21876 11008 21907
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 12710 21876 12716 21888
rect 10980 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 13354 21836 13360 21888
rect 13412 21876 13418 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 13412 21848 13645 21876
rect 13412 21836 13418 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 14550 21836 14556 21888
rect 14608 21876 14614 21888
rect 16040 21885 16068 21984
rect 18598 21972 18604 22024
rect 18656 22012 18662 22024
rect 19242 22012 19248 22024
rect 18656 21984 19248 22012
rect 18656 21972 18662 21984
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19392 21984 20361 22012
rect 19392 21972 19398 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 22940 22012 22968 22052
rect 23431 22049 23443 22052
rect 23477 22049 23480 22083
rect 23431 22043 23480 22049
rect 23474 22040 23480 22043
rect 23532 22080 23538 22092
rect 25240 22089 25268 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 25225 22083 25283 22089
rect 23532 22052 24992 22080
rect 23532 22040 23538 22052
rect 22428 21984 22968 22012
rect 23201 22015 23259 22021
rect 22428 21972 22434 21984
rect 23201 21981 23213 22015
rect 23247 22012 23259 22015
rect 24210 22012 24216 22024
rect 23247 21984 24216 22012
rect 23247 21981 23259 21984
rect 23201 21975 23259 21981
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 24964 22021 24992 22052
rect 25225 22049 25237 22083
rect 25271 22080 25283 22083
rect 25271 22052 25305 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 16574 21904 16580 21956
rect 16632 21944 16638 21956
rect 16632 21916 17724 21944
rect 16632 21904 16638 21916
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 14608 21848 16037 21876
rect 14608 21836 14614 21848
rect 16025 21845 16037 21848
rect 16071 21845 16083 21879
rect 16025 21839 16083 21845
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 16942 21836 16948 21888
rect 17000 21836 17006 21888
rect 17696 21885 17724 21916
rect 17770 21904 17776 21956
rect 17828 21944 17834 21956
rect 17828 21916 19334 21944
rect 17828 21904 17834 21916
rect 17681 21879 17739 21885
rect 17681 21845 17693 21879
rect 17727 21845 17739 21879
rect 17681 21839 17739 21845
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 17920 21848 18061 21876
rect 17920 21836 17926 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18506 21876 18512 21888
rect 18196 21848 18512 21876
rect 18196 21836 18202 21848
rect 18506 21836 18512 21848
rect 18564 21836 18570 21888
rect 19306 21876 19334 21916
rect 19518 21904 19524 21956
rect 19576 21904 19582 21956
rect 21082 21904 21088 21956
rect 21140 21904 21146 21956
rect 21910 21904 21916 21956
rect 21968 21944 21974 21956
rect 25130 21944 25136 21956
rect 21968 21916 25136 21944
rect 21968 21904 21974 21916
rect 19981 21879 20039 21885
rect 19981 21876 19993 21879
rect 19306 21848 19993 21876
rect 19981 21845 19993 21848
rect 20027 21845 20039 21879
rect 19981 21839 20039 21845
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 21634 21876 21640 21888
rect 20128 21848 21640 21876
rect 20128 21836 20134 21848
rect 21634 21836 21640 21848
rect 21692 21836 21698 21888
rect 22112 21885 22140 21916
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22143 21848 22177 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 24486 21836 24492 21888
rect 24544 21876 24550 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 24544 21848 24593 21876
rect 24544 21836 24550 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25590 21876 25596 21888
rect 25087 21848 25596 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 6730 21672 6736 21684
rect 2976 21644 6736 21672
rect 1394 21564 1400 21616
rect 1452 21604 1458 21616
rect 1673 21607 1731 21613
rect 1673 21604 1685 21607
rect 1452 21576 1685 21604
rect 1452 21564 1458 21576
rect 1673 21573 1685 21576
rect 1719 21604 1731 21607
rect 2133 21607 2191 21613
rect 2133 21604 2145 21607
rect 1719 21576 2145 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 2133 21573 2145 21576
rect 2179 21573 2191 21607
rect 2133 21567 2191 21573
rect 2976 21545 3004 21644
rect 6730 21632 6736 21644
rect 6788 21632 6794 21684
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 7282 21672 7288 21684
rect 6972 21644 7288 21672
rect 6972 21632 6978 21644
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 11333 21675 11391 21681
rect 11333 21672 11345 21675
rect 11195 21644 11345 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 11333 21641 11345 21644
rect 11379 21672 11391 21675
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 11379 21644 11989 21672
rect 11379 21641 11391 21644
rect 11333 21635 11391 21641
rect 11977 21641 11989 21644
rect 12023 21672 12035 21675
rect 12066 21672 12072 21684
rect 12023 21644 12072 21672
rect 12023 21641 12035 21644
rect 11977 21635 12035 21641
rect 8478 21604 8484 21616
rect 4816 21576 8484 21604
rect 4816 21545 4844 21576
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 10778 21604 10784 21616
rect 10534 21576 10784 21604
rect 10778 21564 10784 21576
rect 10836 21604 10842 21616
rect 11164 21604 11192 21635
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21641 12311 21675
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 12253 21635 12311 21641
rect 12360 21644 12633 21672
rect 10836 21576 11192 21604
rect 10836 21564 10842 21576
rect 11606 21564 11612 21616
rect 11664 21564 11670 21616
rect 12268 21604 12296 21635
rect 12176 21576 12296 21604
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 6733 21539 6791 21545
rect 6733 21536 6745 21539
rect 6144 21508 6745 21536
rect 6144 21496 6150 21508
rect 6733 21505 6745 21508
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 10686 21496 10692 21548
rect 10744 21536 10750 21548
rect 12176 21536 12204 21576
rect 10744 21508 12204 21536
rect 10744 21496 10750 21508
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7340 21440 7665 21468
rect 7340 21428 7346 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 8294 21428 8300 21480
rect 8352 21468 8358 21480
rect 8570 21468 8576 21480
rect 8352 21440 8576 21468
rect 8352 21428 8358 21440
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 10870 21468 10876 21480
rect 9355 21440 10876 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 12360 21468 12388 21644
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 12713 21675 12771 21681
rect 12713 21641 12725 21675
rect 12759 21672 12771 21675
rect 13722 21672 13728 21684
rect 12759 21644 13728 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21641 13875 21675
rect 13817 21635 13875 21641
rect 15013 21675 15071 21681
rect 15013 21641 15025 21675
rect 15059 21672 15071 21675
rect 17310 21672 17316 21684
rect 15059 21644 17316 21672
rect 15059 21641 15071 21644
rect 15013 21635 15071 21641
rect 13832 21604 13860 21635
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 17770 21672 17776 21684
rect 17420 21644 17776 21672
rect 10980 21440 12388 21468
rect 12544 21576 13860 21604
rect 14185 21607 14243 21613
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21400 1915 21403
rect 7926 21400 7932 21412
rect 1903 21372 7932 21400
rect 1903 21369 1915 21372
rect 1857 21363 1915 21369
rect 7926 21360 7932 21372
rect 7984 21360 7990 21412
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 10980 21400 11008 21440
rect 10652 21372 11008 21400
rect 11793 21403 11851 21409
rect 10652 21360 10658 21372
rect 11793 21369 11805 21403
rect 11839 21400 11851 21403
rect 12342 21400 12348 21412
rect 11839 21372 12348 21400
rect 11839 21369 11851 21372
rect 11793 21363 11851 21369
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 12434 21360 12440 21412
rect 12492 21400 12498 21412
rect 12544 21400 12572 21576
rect 14185 21573 14197 21607
rect 14231 21604 14243 21607
rect 14274 21604 14280 21616
rect 14231 21576 14280 21604
rect 14231 21573 14243 21576
rect 14185 21567 14243 21573
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 16482 21604 16488 21616
rect 15304 21576 16488 21604
rect 15304 21536 15332 21576
rect 16482 21564 16488 21576
rect 16540 21564 16546 21616
rect 17420 21604 17448 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 19116 21644 20453 21672
rect 19116 21632 19122 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 20441 21635 20499 21641
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20772 21644 20913 21672
rect 20772 21632 20778 21644
rect 20901 21641 20913 21644
rect 20947 21672 20959 21675
rect 21358 21672 21364 21684
rect 20947 21644 21364 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 21358 21632 21364 21644
rect 21416 21672 21422 21684
rect 22186 21672 22192 21684
rect 21416 21644 22192 21672
rect 21416 21632 21422 21644
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22336 21644 22477 21672
rect 22336 21632 22342 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 17328 21576 17448 21604
rect 14292 21508 15332 21536
rect 12802 21428 12808 21480
rect 12860 21428 12866 21480
rect 13998 21468 14004 21480
rect 13280 21440 14004 21468
rect 12492 21372 12572 21400
rect 12492 21360 12498 21372
rect 6549 21335 6607 21341
rect 6549 21301 6561 21335
rect 6595 21332 6607 21335
rect 6638 21332 6644 21344
rect 6595 21304 6644 21332
rect 6595 21301 6607 21304
rect 6549 21295 6607 21301
rect 6638 21292 6644 21304
rect 6696 21292 6702 21344
rect 8570 21292 8576 21344
rect 8628 21332 8634 21344
rect 10410 21332 10416 21344
rect 8628 21304 10416 21332
rect 8628 21292 8634 21304
rect 10410 21292 10416 21304
rect 10468 21292 10474 21344
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10560 21304 10793 21332
rect 10560 21292 10566 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 10870 21292 10876 21344
rect 10928 21332 10934 21344
rect 11146 21332 11152 21344
rect 10928 21304 11152 21332
rect 10928 21292 10934 21304
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 12066 21292 12072 21344
rect 12124 21332 12130 21344
rect 13280 21332 13308 21440
rect 13998 21428 14004 21440
rect 14056 21428 14062 21480
rect 14292 21477 14320 21508
rect 15378 21496 15384 21548
rect 15436 21496 15442 21548
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 16390 21536 16396 21548
rect 15519 21508 16396 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21437 14335 21471
rect 14277 21431 14335 21437
rect 14461 21471 14519 21477
rect 14461 21437 14473 21471
rect 14507 21468 14519 21471
rect 15102 21468 15108 21480
rect 14507 21440 15108 21468
rect 14507 21437 14519 21440
rect 14461 21431 14519 21437
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15654 21428 15660 21480
rect 15712 21428 15718 21480
rect 15930 21428 15936 21480
rect 15988 21468 15994 21480
rect 16025 21471 16083 21477
rect 16025 21468 16037 21471
rect 15988 21440 16037 21468
rect 15988 21428 15994 21440
rect 16025 21437 16037 21440
rect 16071 21437 16083 21471
rect 16025 21431 16083 21437
rect 16298 21428 16304 21480
rect 16356 21468 16362 21480
rect 17328 21468 17356 21576
rect 17494 21564 17500 21616
rect 17552 21564 17558 21616
rect 18233 21607 18291 21613
rect 18233 21573 18245 21607
rect 18279 21604 18291 21607
rect 18506 21604 18512 21616
rect 18279 21576 18512 21604
rect 18279 21573 18291 21576
rect 18233 21567 18291 21573
rect 18506 21564 18512 21576
rect 18564 21604 18570 21616
rect 21450 21604 21456 21616
rect 18564 21576 21456 21604
rect 18564 21564 18570 21576
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 21634 21564 21640 21616
rect 21692 21604 21698 21616
rect 21692 21576 22600 21604
rect 21692 21564 21698 21576
rect 17402 21496 17408 21548
rect 17460 21496 17466 21548
rect 17512 21536 17540 21564
rect 20438 21536 20444 21548
rect 17512 21508 20444 21536
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 22370 21496 22376 21548
rect 22428 21496 22434 21548
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 16356 21440 17509 21468
rect 16356 21428 16362 21440
rect 17497 21437 17509 21440
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 17678 21428 17684 21480
rect 17736 21428 17742 21480
rect 19426 21468 19432 21480
rect 17926 21440 19432 21468
rect 13357 21403 13415 21409
rect 13357 21369 13369 21403
rect 13403 21400 13415 21403
rect 13538 21400 13544 21412
rect 13403 21372 13544 21400
rect 13403 21369 13415 21372
rect 13357 21363 13415 21369
rect 13538 21360 13544 21372
rect 13596 21360 13602 21412
rect 13814 21360 13820 21412
rect 13872 21400 13878 21412
rect 17770 21400 17776 21412
rect 13872 21372 17776 21400
rect 13872 21360 13878 21372
rect 17770 21360 17776 21372
rect 17828 21360 17834 21412
rect 12124 21304 13308 21332
rect 12124 21292 12130 21304
rect 13446 21292 13452 21344
rect 13504 21332 13510 21344
rect 15562 21332 15568 21344
rect 13504 21304 15568 21332
rect 13504 21292 13510 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16390 21332 16396 21344
rect 16347 21304 16396 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 16632 21304 16681 21332
rect 16632 21292 16638 21304
rect 16669 21301 16681 21304
rect 16715 21332 16727 21335
rect 16758 21332 16764 21344
rect 16715 21304 16764 21332
rect 16715 21301 16727 21304
rect 16669 21295 16727 21301
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 17926 21332 17954 21440
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 22388 21468 22416 21496
rect 22572 21477 22600 21576
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 23934 21564 23940 21616
rect 23992 21604 23998 21616
rect 23992 21576 24150 21604
rect 23992 21564 23998 21576
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 21560 21440 22416 21468
rect 22557 21471 22615 21477
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 21560 21400 21588 21440
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 24670 21468 24676 21480
rect 22557 21431 22615 21437
rect 22664 21440 24676 21468
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 19208 21372 21588 21400
rect 21652 21372 22017 21400
rect 19208 21360 19214 21372
rect 17083 21304 17954 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19521 21295 19579 21301
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 21652 21332 21680 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 22186 21360 22192 21412
rect 22244 21400 22250 21412
rect 22664 21400 22692 21440
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 22244 21372 22692 21400
rect 22244 21360 22250 21372
rect 20036 21304 21680 21332
rect 20036 21292 20042 21304
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 22554 21332 22560 21344
rect 21968 21304 22560 21332
rect 21968 21292 21974 21304
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 23017 21335 23075 21341
rect 23017 21332 23029 21335
rect 22888 21304 23029 21332
rect 22888 21292 22894 21304
rect 23017 21301 23029 21304
rect 23063 21301 23075 21335
rect 23017 21295 23075 21301
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 23808 21304 25145 21332
rect 23808 21292 23814 21304
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 25406 21292 25412 21344
rect 25464 21292 25470 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 5810 21088 5816 21140
rect 5868 21088 5874 21140
rect 8665 21131 8723 21137
rect 8665 21097 8677 21131
rect 8711 21128 8723 21131
rect 9122 21128 9128 21140
rect 8711 21100 9128 21128
rect 8711 21097 8723 21100
rect 8665 21091 8723 21097
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 10520 21100 13584 21128
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 2832 21032 2912 21060
rect 2832 21020 2838 21032
rect 2884 21001 2912 21032
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 6273 21063 6331 21069
rect 6273 21060 6285 21063
rect 5224 21032 6285 21060
rect 5224 21020 5230 21032
rect 6273 21029 6285 21032
rect 6319 21029 6331 21063
rect 6273 21023 6331 21029
rect 6472 21032 8432 21060
rect 2869 20995 2927 21001
rect 2240 20964 2774 20992
rect 2240 20933 2268 20964
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2746 20856 2774 20964
rect 2869 20961 2881 20995
rect 2915 20961 2927 20995
rect 2869 20955 2927 20961
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 5810 20924 5816 20936
rect 4111 20896 5816 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 6472 20933 6500 21032
rect 6546 20952 6552 21004
rect 6604 20992 6610 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6604 20964 7389 20992
rect 6604 20952 6610 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 8404 20992 8432 21032
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 9953 21063 10011 21069
rect 9953 21060 9965 21063
rect 8536 21032 9965 21060
rect 8536 21020 8542 21032
rect 9953 21029 9965 21032
rect 9999 21029 10011 21063
rect 10520 21060 10548 21100
rect 9953 21023 10011 21029
rect 10428 21032 10548 21060
rect 9214 20992 9220 21004
rect 8404 20964 9220 20992
rect 7377 20955 7435 20961
rect 9214 20952 9220 20964
rect 9272 20952 9278 21004
rect 10042 20952 10048 21004
rect 10100 20992 10106 21004
rect 10428 21001 10456 21032
rect 12710 21020 12716 21072
rect 12768 21060 12774 21072
rect 12897 21063 12955 21069
rect 12897 21060 12909 21063
rect 12768 21032 12909 21060
rect 12768 21020 12774 21032
rect 12897 21029 12909 21032
rect 12943 21029 12955 21063
rect 13556 21060 13584 21100
rect 13630 21088 13636 21140
rect 13688 21088 13694 21140
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 13780 21100 16681 21128
rect 13780 21088 13786 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 16850 21088 16856 21140
rect 16908 21128 16914 21140
rect 16908 21100 17724 21128
rect 16908 21088 16914 21100
rect 15473 21063 15531 21069
rect 15473 21060 15485 21063
rect 13556 21032 15485 21060
rect 12897 21023 12955 21029
rect 15473 21029 15485 21032
rect 15519 21029 15531 21063
rect 15473 21023 15531 21029
rect 16758 21020 16764 21072
rect 16816 21060 16822 21072
rect 17034 21060 17040 21072
rect 16816 21032 17040 21060
rect 16816 21020 16822 21032
rect 17034 21020 17040 21032
rect 17092 21020 17098 21072
rect 10413 20995 10471 21001
rect 10100 20964 10364 20992
rect 10100 20952 10106 20964
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7340 20896 7880 20924
rect 7340 20884 7346 20896
rect 7650 20856 7656 20868
rect 2746 20828 7656 20856
rect 7650 20816 7656 20828
rect 7708 20816 7714 20868
rect 7852 20856 7880 20896
rect 7926 20884 7932 20936
rect 7984 20924 7990 20936
rect 9766 20924 9772 20936
rect 7984 20896 9772 20924
rect 7984 20884 7990 20896
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 10336 20933 10364 20964
rect 10413 20961 10425 20995
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10502 20952 10508 21004
rect 10560 20952 10566 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 11112 20964 11161 20992
rect 11112 20952 11118 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20992 11483 20995
rect 12802 20992 12808 21004
rect 11471 20964 12808 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 12802 20952 12808 20964
rect 12860 20992 12866 21004
rect 13630 20992 13636 21004
rect 12860 20964 13636 20992
rect 12860 20952 12866 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 14090 20952 14096 21004
rect 14148 20992 14154 21004
rect 16025 20995 16083 21001
rect 16025 20992 16037 20995
rect 14148 20964 16037 20992
rect 14148 20952 14154 20964
rect 16025 20961 16037 20964
rect 16071 20961 16083 20995
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 16025 20955 16083 20961
rect 16132 20964 17233 20992
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 14369 20927 14427 20933
rect 13228 20896 14136 20924
rect 13228 20884 13234 20896
rect 8941 20859 8999 20865
rect 8941 20856 8953 20859
rect 7852 20828 8953 20856
rect 8941 20825 8953 20828
rect 8987 20825 8999 20859
rect 8941 20819 8999 20825
rect 9309 20859 9367 20865
rect 9309 20825 9321 20859
rect 9355 20856 9367 20859
rect 12894 20856 12900 20868
rect 9355 20828 10916 20856
rect 12650 20828 12900 20856
rect 9355 20825 9367 20828
rect 9309 20819 9367 20825
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 4028 20760 5733 20788
rect 4028 20748 4034 20760
rect 5721 20757 5733 20760
rect 5767 20788 5779 20791
rect 8846 20788 8852 20800
rect 5767 20760 8852 20788
rect 5767 20757 5779 20760
rect 5721 20751 5779 20757
rect 8846 20748 8852 20760
rect 8904 20748 8910 20800
rect 8956 20788 8984 20819
rect 10594 20788 10600 20800
rect 8956 20760 10600 20788
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 10888 20788 10916 20828
rect 12894 20816 12900 20828
rect 12952 20856 12958 20868
rect 13446 20856 13452 20868
rect 12952 20828 13452 20856
rect 12952 20816 12958 20828
rect 13446 20816 13452 20828
rect 13504 20816 13510 20868
rect 13538 20816 13544 20868
rect 13596 20816 13602 20868
rect 14108 20856 14136 20896
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14826 20924 14832 20936
rect 14415 20896 14832 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 15930 20884 15936 20936
rect 15988 20884 15994 20936
rect 14108 20828 14583 20856
rect 12434 20788 12440 20800
rect 10888 20760 12440 20788
rect 12434 20748 12440 20760
rect 12492 20748 12498 20800
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 13722 20788 13728 20800
rect 13412 20760 13728 20788
rect 13412 20748 13418 20760
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 14458 20748 14464 20800
rect 14516 20748 14522 20800
rect 14555 20788 14583 20828
rect 14642 20816 14648 20868
rect 14700 20856 14706 20868
rect 16132 20856 16160 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 17696 20992 17724 21100
rect 17770 21088 17776 21140
rect 17828 21128 17834 21140
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 17828 21100 17877 21128
rect 17828 21088 17834 21100
rect 17865 21097 17877 21100
rect 17911 21097 17923 21131
rect 22370 21128 22376 21140
rect 17865 21091 17923 21097
rect 18340 21100 22376 21128
rect 17770 20992 17776 21004
rect 17696 20964 17776 20992
rect 17221 20955 17279 20961
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 18340 21001 18368 21100
rect 22370 21088 22376 21100
rect 22428 21088 22434 21140
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 22833 21131 22891 21137
rect 22833 21128 22845 21131
rect 22520 21100 22845 21128
rect 22520 21088 22526 21100
rect 22833 21097 22845 21100
rect 22879 21097 22891 21131
rect 22833 21091 22891 21097
rect 18782 21020 18788 21072
rect 18840 21060 18846 21072
rect 18877 21063 18935 21069
rect 18877 21060 18889 21063
rect 18840 21032 18889 21060
rect 18840 21020 18846 21032
rect 18877 21029 18889 21032
rect 18923 21029 18935 21063
rect 18877 21023 18935 21029
rect 21174 21020 21180 21072
rect 21232 21060 21238 21072
rect 21232 21032 23428 21060
rect 21232 21020 21238 21032
rect 18325 20995 18383 21001
rect 18325 20961 18337 20995
rect 18371 20961 18383 20995
rect 18325 20955 18383 20961
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20992 18754 21004
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 18748 20964 19717 20992
rect 18748 20952 18754 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 21634 20952 21640 21004
rect 21692 20992 21698 21004
rect 23400 21001 23428 21032
rect 23934 21020 23940 21072
rect 23992 21060 23998 21072
rect 24029 21063 24087 21069
rect 24029 21060 24041 21063
rect 23992 21032 24041 21060
rect 23992 21020 23998 21032
rect 24029 21029 24041 21032
rect 24075 21060 24087 21063
rect 24118 21060 24124 21072
rect 24075 21032 24124 21060
rect 24075 21029 24087 21032
rect 24029 21023 24087 21029
rect 24118 21020 24124 21032
rect 24176 21060 24182 21072
rect 24394 21060 24400 21072
rect 24176 21032 24400 21060
rect 24176 21020 24182 21032
rect 24394 21020 24400 21032
rect 24452 21020 24458 21072
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 21692 20964 22201 20992
rect 21692 20952 21698 20964
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 23293 20995 23351 21001
rect 23293 20992 23305 20995
rect 22189 20955 22247 20961
rect 22296 20964 23305 20992
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17862 20924 17868 20936
rect 17000 20896 17868 20924
rect 17000 20884 17006 20896
rect 17862 20884 17868 20896
rect 17920 20884 17926 20936
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18414 20924 18420 20936
rect 18279 20896 18420 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 21910 20884 21916 20936
rect 21968 20924 21974 20936
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21968 20896 22017 20924
rect 21968 20884 21974 20896
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22094 20884 22100 20936
rect 22152 20884 22158 20936
rect 14700 20828 16160 20856
rect 17037 20859 17095 20865
rect 14700 20816 14706 20828
rect 17037 20825 17049 20859
rect 17083 20856 17095 20859
rect 17310 20856 17316 20868
rect 17083 20828 17316 20856
rect 17083 20825 17095 20828
rect 17037 20819 17095 20825
rect 17310 20816 17316 20828
rect 17368 20816 17374 20868
rect 21082 20856 21088 20868
rect 20930 20828 21088 20856
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21192 20828 21772 20856
rect 14829 20791 14887 20797
rect 14829 20788 14841 20791
rect 14555 20760 14841 20788
rect 14829 20757 14841 20760
rect 14875 20788 14887 20791
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14875 20760 15025 20788
rect 14875 20757 14887 20760
rect 14829 20751 14887 20757
rect 15013 20757 15025 20760
rect 15059 20788 15071 20791
rect 15378 20788 15384 20800
rect 15059 20760 15384 20788
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16206 20788 16212 20800
rect 15988 20760 16212 20788
rect 15988 20748 15994 20760
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 16390 20748 16396 20800
rect 16448 20788 16454 20800
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16448 20760 17141 20788
rect 16448 20748 16454 20760
rect 17129 20757 17141 20760
rect 17175 20757 17187 20791
rect 17129 20751 17187 20757
rect 19242 20748 19248 20800
rect 19300 20788 19306 20800
rect 19794 20788 19800 20800
rect 19300 20760 19800 20788
rect 19300 20748 19306 20760
rect 19794 20748 19800 20760
rect 19852 20788 19858 20800
rect 21192 20788 21220 20828
rect 19852 20760 21220 20788
rect 19852 20748 19858 20760
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 21637 20791 21695 20797
rect 21637 20788 21649 20791
rect 21416 20760 21649 20788
rect 21416 20748 21422 20760
rect 21637 20757 21649 20760
rect 21683 20757 21695 20791
rect 21744 20788 21772 20828
rect 22296 20788 22324 20964
rect 23293 20961 23305 20964
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 23658 20952 23664 21004
rect 23716 20992 23722 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 23716 20964 25145 20992
rect 23716 20952 23722 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 23106 20924 23112 20936
rect 22428 20896 23112 20924
rect 22428 20884 22434 20896
rect 23106 20884 23112 20896
rect 23164 20884 23170 20936
rect 23198 20884 23204 20936
rect 23256 20884 23262 20936
rect 24670 20884 24676 20936
rect 24728 20924 24734 20936
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24728 20896 25053 20924
rect 24728 20884 24734 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 24397 20859 24455 20865
rect 24397 20856 24409 20859
rect 23440 20828 24409 20856
rect 23440 20816 23446 20828
rect 24397 20825 24409 20828
rect 24443 20856 24455 20859
rect 24949 20859 25007 20865
rect 24949 20856 24961 20859
rect 24443 20828 24961 20856
rect 24443 20825 24455 20828
rect 24397 20819 24455 20825
rect 24949 20825 24961 20828
rect 24995 20825 25007 20859
rect 24949 20819 25007 20825
rect 21744 20760 22324 20788
rect 21637 20751 21695 20757
rect 23106 20748 23112 20800
rect 23164 20788 23170 20800
rect 24581 20791 24639 20797
rect 24581 20788 24593 20791
rect 23164 20760 24593 20788
rect 23164 20748 23170 20760
rect 24581 20757 24593 20760
rect 24627 20757 24639 20791
rect 24581 20751 24639 20757
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 25958 20788 25964 20800
rect 24912 20760 25964 20788
rect 24912 20748 24918 20760
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 26050 20680 26056 20732
rect 26108 20720 26114 20732
rect 26418 20720 26424 20732
rect 26108 20692 26424 20720
rect 26108 20680 26114 20692
rect 26418 20680 26424 20692
rect 26476 20680 26482 20732
rect 1104 20624 25852 20646
rect 6457 20587 6515 20593
rect 6457 20553 6469 20587
rect 6503 20584 6515 20587
rect 6822 20584 6828 20596
rect 6503 20556 6828 20584
rect 6503 20553 6515 20556
rect 6457 20547 6515 20553
rect 6822 20544 6828 20556
rect 6880 20584 6886 20596
rect 7282 20584 7288 20596
rect 6880 20556 7288 20584
rect 6880 20544 6886 20556
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 10042 20584 10048 20596
rect 7791 20556 10048 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 10962 20544 10968 20596
rect 11020 20584 11026 20596
rect 12069 20587 12127 20593
rect 12069 20584 12081 20587
rect 11020 20556 12081 20584
rect 11020 20544 11026 20556
rect 12069 20553 12081 20556
rect 12115 20553 12127 20587
rect 12069 20547 12127 20553
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 13170 20544 13176 20596
rect 13228 20544 13234 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14182 20584 14188 20596
rect 13872 20556 14188 20584
rect 13872 20544 13878 20556
rect 14182 20544 14188 20556
rect 14240 20584 14246 20596
rect 14240 20556 16528 20584
rect 14240 20544 14246 20556
rect 1673 20519 1731 20525
rect 1673 20485 1685 20519
rect 1719 20516 1731 20519
rect 2133 20519 2191 20525
rect 2133 20516 2145 20519
rect 1719 20488 2145 20516
rect 1719 20485 1731 20488
rect 1673 20479 1731 20485
rect 2133 20485 2145 20488
rect 2179 20516 2191 20519
rect 3418 20516 3424 20528
rect 2179 20488 3424 20516
rect 2179 20485 2191 20488
rect 2133 20479 2191 20485
rect 3418 20476 3424 20488
rect 3476 20476 3482 20528
rect 4890 20476 4896 20528
rect 4948 20476 4954 20528
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 5169 20519 5227 20525
rect 5169 20516 5181 20519
rect 5123 20488 5181 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 5169 20485 5181 20488
rect 5215 20516 5227 20519
rect 5350 20516 5356 20528
rect 5215 20488 5356 20516
rect 5215 20485 5227 20488
rect 5169 20479 5227 20485
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 9582 20516 9588 20528
rect 7300 20488 9588 20516
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 5534 20448 5540 20460
rect 3099 20420 5540 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20448 6055 20451
rect 7006 20448 7012 20460
rect 6043 20420 7012 20448
rect 6043 20417 6055 20420
rect 5997 20411 6055 20417
rect 7006 20408 7012 20420
rect 7064 20408 7070 20460
rect 7300 20457 7328 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 10594 20516 10600 20528
rect 10534 20488 10600 20516
rect 10594 20476 10600 20488
rect 10652 20516 10658 20528
rect 11054 20516 11060 20528
rect 10652 20488 11060 20516
rect 10652 20476 10658 20488
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 11793 20519 11851 20525
rect 11793 20485 11805 20519
rect 11839 20516 11851 20519
rect 11974 20516 11980 20528
rect 11839 20488 11980 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 11974 20476 11980 20488
rect 12032 20476 12038 20528
rect 12529 20519 12587 20525
rect 12529 20485 12541 20519
rect 12575 20516 12587 20519
rect 13832 20516 13860 20544
rect 15194 20516 15200 20528
rect 12575 20488 13492 20516
rect 12575 20485 12587 20488
rect 12529 20479 12587 20485
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 8570 20408 8576 20460
rect 8628 20408 8634 20460
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 6641 20383 6699 20389
rect 6641 20349 6653 20383
rect 6687 20380 6699 20383
rect 7926 20380 7932 20392
rect 6687 20352 7932 20380
rect 6687 20349 6699 20352
rect 6641 20343 6699 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 10502 20380 10508 20392
rect 9355 20352 10508 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 1857 20315 1915 20321
rect 1857 20281 1869 20315
rect 1903 20312 1915 20315
rect 1903 20284 2774 20312
rect 1903 20281 1915 20284
rect 1857 20275 1915 20281
rect 2746 20244 2774 20284
rect 4246 20272 4252 20324
rect 4304 20312 4310 20324
rect 5813 20315 5871 20321
rect 5813 20312 5825 20315
rect 4304 20284 5825 20312
rect 4304 20272 4310 20284
rect 5813 20281 5825 20284
rect 5859 20281 5871 20315
rect 5813 20275 5871 20281
rect 6825 20315 6883 20321
rect 6825 20281 6837 20315
rect 6871 20312 6883 20315
rect 13354 20312 13360 20324
rect 6871 20284 8524 20312
rect 6871 20281 6883 20284
rect 6825 20275 6883 20281
rect 6840 20244 6868 20275
rect 2746 20216 6868 20244
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6972 20216 7113 20244
rect 6972 20204 6978 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 8389 20247 8447 20253
rect 8389 20244 8401 20247
rect 7248 20216 8401 20244
rect 7248 20204 7254 20216
rect 8389 20213 8401 20216
rect 8435 20213 8447 20247
rect 8496 20244 8524 20284
rect 10704 20284 13360 20312
rect 10704 20244 10732 20284
rect 13354 20272 13360 20284
rect 13412 20272 13418 20324
rect 8496 20216 10732 20244
rect 8389 20207 8447 20213
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11149 20247 11207 20253
rect 11149 20244 11161 20247
rect 11112 20216 11161 20244
rect 11112 20204 11118 20216
rect 11149 20213 11161 20216
rect 11195 20244 11207 20247
rect 11333 20247 11391 20253
rect 11333 20244 11345 20247
rect 11195 20216 11345 20244
rect 11195 20213 11207 20216
rect 11149 20207 11207 20213
rect 11333 20213 11345 20216
rect 11379 20244 11391 20247
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11379 20216 11621 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 11609 20213 11621 20216
rect 11655 20244 11667 20247
rect 12434 20244 12440 20256
rect 11655 20216 12440 20244
rect 11655 20213 11667 20216
rect 11609 20207 11667 20213
rect 12434 20204 12440 20216
rect 12492 20244 12498 20256
rect 12894 20244 12900 20256
rect 12492 20216 12900 20244
rect 12492 20204 12498 20216
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 13464 20244 13492 20488
rect 13556 20488 13860 20516
rect 15042 20488 15200 20516
rect 13556 20457 13584 20488
rect 15194 20476 15200 20488
rect 15252 20516 15258 20528
rect 15562 20516 15568 20528
rect 15252 20488 15568 20516
rect 15252 20476 15258 20488
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 16500 20460 16528 20556
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 18138 20584 18144 20596
rect 17276 20556 18144 20584
rect 17276 20544 17282 20556
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 20993 20587 21051 20593
rect 18932 20556 20852 20584
rect 18932 20544 18938 20556
rect 18782 20516 18788 20528
rect 18446 20502 18788 20516
rect 18432 20488 18788 20502
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 15470 20408 15476 20460
rect 15528 20448 15534 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15528 20420 15853 20448
rect 15528 20408 15534 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16540 20420 16957 20448
rect 16540 20408 16546 20420
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 14550 20380 14556 20392
rect 13863 20352 14556 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 15010 20340 15016 20392
rect 15068 20380 15074 20392
rect 16758 20380 16764 20392
rect 15068 20352 16764 20380
rect 15068 20340 15074 20352
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 18230 20380 18236 20392
rect 17267 20352 18236 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 18230 20340 18236 20352
rect 18288 20340 18294 20392
rect 15102 20272 15108 20324
rect 15160 20312 15166 20324
rect 15289 20315 15347 20321
rect 15289 20312 15301 20315
rect 15160 20284 15301 20312
rect 15160 20272 15166 20284
rect 15289 20281 15301 20284
rect 15335 20281 15347 20315
rect 15289 20275 15347 20281
rect 15838 20244 15844 20256
rect 13464 20216 15844 20244
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 15930 20204 15936 20256
rect 15988 20204 15994 20256
rect 16393 20247 16451 20253
rect 16393 20213 16405 20247
rect 16439 20244 16451 20247
rect 17034 20244 17040 20256
rect 16439 20216 17040 20244
rect 16439 20213 16451 20216
rect 16393 20207 16451 20213
rect 17034 20204 17040 20216
rect 17092 20244 17098 20256
rect 18432 20244 18460 20488
rect 18782 20476 18788 20488
rect 18840 20516 18846 20528
rect 18840 20488 20010 20516
rect 18840 20476 18846 20488
rect 20824 20448 20852 20556
rect 20993 20553 21005 20587
rect 21039 20584 21051 20587
rect 21266 20584 21272 20596
rect 21039 20556 21272 20584
rect 21039 20553 21051 20556
rect 20993 20547 21051 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 21910 20584 21916 20596
rect 21416 20556 21916 20584
rect 21416 20544 21422 20556
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22462 20584 22468 20596
rect 22143 20556 22468 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 22554 20544 22560 20596
rect 22612 20584 22618 20596
rect 25406 20584 25412 20596
rect 22612 20556 25412 20584
rect 22612 20544 22618 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 20898 20476 20904 20528
rect 20956 20516 20962 20528
rect 23658 20516 23664 20528
rect 20956 20488 23664 20516
rect 20956 20476 20962 20488
rect 23658 20476 23664 20488
rect 23716 20476 23722 20528
rect 23750 20476 23756 20528
rect 23808 20476 23814 20528
rect 24394 20476 24400 20528
rect 24452 20476 24458 20528
rect 22370 20448 22376 20460
rect 20824 20420 22376 20448
rect 22370 20408 22376 20420
rect 22428 20448 22434 20460
rect 22465 20451 22523 20457
rect 22465 20448 22477 20451
rect 22428 20420 22477 20448
rect 22428 20408 22434 20420
rect 22465 20417 22477 20420
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 22554 20380 22560 20392
rect 20220 20352 22560 20380
rect 20220 20340 20226 20352
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 22646 20340 22652 20392
rect 22704 20340 22710 20392
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 21453 20315 21511 20321
rect 21453 20312 21465 20315
rect 20772 20284 21465 20312
rect 20772 20272 20778 20284
rect 21453 20281 21465 20284
rect 21499 20281 21511 20315
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 21453 20275 21511 20281
rect 22066 20284 23121 20312
rect 17092 20216 18460 20244
rect 17092 20204 17098 20216
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 20530 20244 20536 20256
rect 19668 20216 20536 20244
rect 19668 20204 19674 20216
rect 20530 20204 20536 20216
rect 20588 20244 20594 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 20588 20216 21281 20244
rect 20588 20204 20594 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 21818 20244 21824 20256
rect 21416 20216 21824 20244
rect 21416 20204 21422 20216
rect 21818 20204 21824 20216
rect 21876 20244 21882 20256
rect 22066 20244 22094 20284
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 21876 20216 22094 20244
rect 21876 20204 21882 20216
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 23842 20244 23848 20256
rect 22520 20216 23848 20244
rect 22520 20204 22526 20216
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 10413 20043 10471 20049
rect 10413 20040 10425 20043
rect 7064 20012 10425 20040
rect 7064 20000 7070 20012
rect 10413 20009 10425 20012
rect 10459 20009 10471 20043
rect 10413 20003 10471 20009
rect 11422 20000 11428 20052
rect 11480 20040 11486 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 11480 20012 14933 20040
rect 11480 20000 11486 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 15896 20012 17693 20040
rect 15896 20000 15902 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18230 20040 18236 20052
rect 18012 20012 18236 20040
rect 18012 20000 18018 20012
rect 18230 20000 18236 20012
rect 18288 20040 18294 20052
rect 20898 20040 20904 20052
rect 18288 20012 20904 20040
rect 18288 20000 18294 20012
rect 20898 20000 20904 20012
rect 20956 20000 20962 20052
rect 21348 20043 21406 20049
rect 21348 20009 21360 20043
rect 21394 20040 21406 20043
rect 23934 20040 23940 20052
rect 21394 20012 23940 20040
rect 21394 20009 21406 20012
rect 21348 20003 21406 20009
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 4525 19975 4583 19981
rect 4525 19941 4537 19975
rect 4571 19972 4583 19975
rect 7650 19972 7656 19984
rect 4571 19944 7656 19972
rect 4571 19941 4583 19944
rect 4525 19935 4583 19941
rect 7650 19932 7656 19944
rect 7708 19932 7714 19984
rect 7926 19932 7932 19984
rect 7984 19972 7990 19984
rect 11514 19972 11520 19984
rect 7984 19944 11520 19972
rect 7984 19932 7990 19944
rect 11514 19932 11520 19944
rect 11572 19932 11578 19984
rect 13357 19975 13415 19981
rect 13357 19941 13369 19975
rect 13403 19972 13415 19975
rect 13630 19972 13636 19984
rect 13403 19944 13636 19972
rect 13403 19941 13415 19944
rect 13357 19935 13415 19941
rect 13630 19932 13636 19944
rect 13688 19932 13694 19984
rect 14366 19932 14372 19984
rect 14424 19972 14430 19984
rect 14424 19944 15608 19972
rect 14424 19932 14430 19944
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2501 19907 2559 19913
rect 2501 19904 2513 19907
rect 2096 19876 2513 19904
rect 2096 19864 2102 19876
rect 2501 19873 2513 19876
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 5166 19864 5172 19916
rect 5224 19864 5230 19916
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19904 5503 19907
rect 6178 19904 6184 19916
rect 5491 19876 6184 19904
rect 5491 19873 5503 19876
rect 5445 19867 5503 19873
rect 6178 19864 6184 19876
rect 6236 19864 6242 19916
rect 7377 19907 7435 19913
rect 6656 19876 7328 19904
rect 2222 19796 2228 19848
rect 2280 19796 2286 19848
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4890 19836 4896 19848
rect 4755 19808 4896 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 6656 19845 6684 19876
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7300 19836 7328 19876
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 7466 19904 7472 19916
rect 7423 19876 7472 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 10778 19864 10784 19916
rect 10836 19864 10842 19916
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 11072 19876 15485 19904
rect 7834 19836 7840 19848
rect 7300 19808 7840 19836
rect 7101 19799 7159 19805
rect 5350 19660 5356 19712
rect 5408 19700 5414 19712
rect 6457 19703 6515 19709
rect 6457 19700 6469 19703
rect 5408 19672 6469 19700
rect 5408 19660 5414 19672
rect 6457 19669 6469 19672
rect 6503 19669 6515 19703
rect 7116 19700 7144 19799
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 10796 19836 10824 19864
rect 11072 19836 11100 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15580 19904 15608 19944
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 18782 19972 18788 19984
rect 17184 19944 18788 19972
rect 17184 19932 17190 19944
rect 18782 19932 18788 19944
rect 18840 19972 18846 19984
rect 18877 19975 18935 19981
rect 18877 19972 18889 19975
rect 18840 19944 18889 19972
rect 18840 19932 18846 19944
rect 18877 19941 18889 19944
rect 18923 19941 18935 19975
rect 19150 19972 19156 19984
rect 18877 19935 18935 19941
rect 18984 19944 19156 19972
rect 17221 19907 17279 19913
rect 17221 19904 17233 19907
rect 15580 19876 17233 19904
rect 15473 19867 15531 19873
rect 17221 19873 17233 19876
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18138 19864 18144 19916
rect 18196 19864 18202 19916
rect 18230 19864 18236 19916
rect 18288 19864 18294 19916
rect 18690 19864 18696 19916
rect 18748 19864 18754 19916
rect 10796 19808 11100 19836
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 13998 19836 14004 19848
rect 13188 19808 14004 19836
rect 8389 19771 8447 19777
rect 8389 19737 8401 19771
rect 8435 19768 8447 19771
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 8435 19740 10793 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 10781 19731 10839 19737
rect 10873 19771 10931 19777
rect 10873 19737 10885 19771
rect 10919 19768 10931 19771
rect 11422 19768 11428 19780
rect 10919 19740 11428 19768
rect 10919 19737 10931 19740
rect 10873 19731 10931 19737
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 11885 19771 11943 19777
rect 11885 19737 11897 19771
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 7466 19700 7472 19712
rect 7116 19672 7472 19700
rect 6457 19663 6515 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8202 19700 8208 19712
rect 7708 19672 8208 19700
rect 7708 19660 7714 19672
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 9122 19660 9128 19712
rect 9180 19660 9186 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 11146 19700 11152 19712
rect 9815 19672 11152 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11900 19700 11928 19731
rect 12434 19728 12440 19780
rect 12492 19728 12498 19780
rect 13188 19700 13216 19808
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 18049 19839 18107 19845
rect 18049 19836 18061 19839
rect 14608 19808 18061 19836
rect 14608 19796 14614 19808
rect 18049 19805 18061 19808
rect 18095 19805 18107 19839
rect 18156 19836 18184 19864
rect 18984 19836 19012 19944
rect 19150 19932 19156 19944
rect 19208 19972 19214 19984
rect 20622 19972 20628 19984
rect 19208 19944 20628 19972
rect 19208 19932 19214 19944
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 20073 19907 20131 19913
rect 20073 19904 20085 19907
rect 18156 19808 19012 19836
rect 19306 19876 20085 19904
rect 18049 19799 18107 19805
rect 13262 19728 13268 19780
rect 13320 19768 13326 19780
rect 14918 19768 14924 19780
rect 13320 19740 14924 19768
rect 13320 19728 13326 19740
rect 14918 19728 14924 19740
rect 14976 19728 14982 19780
rect 15010 19728 15016 19780
rect 15068 19768 15074 19780
rect 15378 19768 15384 19780
rect 15068 19740 15384 19768
rect 15068 19728 15074 19740
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 15930 19728 15936 19780
rect 15988 19768 15994 19780
rect 16173 19771 16231 19777
rect 16173 19768 16185 19771
rect 15988 19740 16185 19768
rect 15988 19728 15994 19740
rect 16173 19737 16185 19740
rect 16219 19737 16231 19771
rect 16173 19731 16231 19737
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17037 19771 17095 19777
rect 17037 19768 17049 19771
rect 16816 19740 17049 19768
rect 16816 19728 16822 19740
rect 17037 19737 17049 19740
rect 17083 19737 17095 19771
rect 19306 19768 19334 19876
rect 20073 19873 20085 19876
rect 20119 19904 20131 19907
rect 20714 19904 20720 19916
rect 20119 19876 20720 19904
rect 20119 19873 20131 19876
rect 20073 19867 20131 19873
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23290 19904 23296 19916
rect 21131 19876 23296 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19904 23995 19907
rect 24394 19904 24400 19916
rect 23983 19876 24400 19904
rect 23983 19873 23995 19876
rect 23937 19867 23995 19873
rect 24394 19864 24400 19876
rect 24452 19864 24458 19916
rect 25038 19864 25044 19916
rect 25096 19864 25102 19916
rect 25130 19864 25136 19916
rect 25188 19864 25194 19916
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19836 19855 19839
rect 20622 19836 20628 19848
rect 19843 19808 20628 19836
rect 19843 19805 19855 19808
rect 19797 19799 19855 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23658 19836 23664 19848
rect 23532 19808 23664 19836
rect 23532 19796 23538 19808
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 17037 19731 17095 19737
rect 17144 19740 19334 19768
rect 11900 19672 13216 19700
rect 13630 19660 13636 19712
rect 13688 19660 13694 19712
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 14458 19700 14464 19712
rect 13955 19672 14464 19700
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 15286 19660 15292 19712
rect 15344 19660 15350 19712
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 16850 19660 16856 19712
rect 16908 19700 16914 19712
rect 17144 19700 17172 19740
rect 19518 19728 19524 19780
rect 19576 19768 19582 19780
rect 20441 19771 20499 19777
rect 20441 19768 20453 19771
rect 19576 19740 20453 19768
rect 19576 19728 19582 19740
rect 20441 19737 20453 19740
rect 20487 19737 20499 19771
rect 20441 19731 20499 19737
rect 21818 19728 21824 19780
rect 21876 19728 21882 19780
rect 24118 19728 24124 19780
rect 24176 19768 24182 19780
rect 25038 19768 25044 19780
rect 24176 19740 25044 19768
rect 24176 19728 24182 19740
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 16908 19672 17172 19700
rect 16908 19660 16914 19672
rect 17218 19660 17224 19712
rect 17276 19700 17282 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 17276 19672 19441 19700
rect 17276 19660 17282 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 19702 19660 19708 19712
rect 19760 19700 19766 19712
rect 19889 19703 19947 19709
rect 19889 19700 19901 19703
rect 19760 19672 19901 19700
rect 19760 19660 19766 19672
rect 19889 19669 19901 19672
rect 19935 19669 19947 19703
rect 19889 19663 19947 19669
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 21692 19672 22845 19700
rect 21692 19660 21698 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 22833 19663 22891 19669
rect 23293 19703 23351 19709
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23474 19700 23480 19712
rect 23339 19672 23480 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24302 19700 24308 19712
rect 23808 19672 24308 19700
rect 23808 19660 23814 19672
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19700 25007 19703
rect 26050 19700 26056 19712
rect 24995 19672 26056 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 26050 19660 26056 19672
rect 26108 19660 26114 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 4614 19496 4620 19508
rect 3988 19468 4620 19496
rect 3988 19428 4016 19468
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 5813 19499 5871 19505
rect 5813 19465 5825 19499
rect 5859 19496 5871 19499
rect 6270 19496 6276 19508
rect 5859 19468 6276 19496
rect 5859 19465 5871 19468
rect 5813 19459 5871 19465
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7282 19496 7288 19508
rect 7147 19468 7288 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 8386 19456 8392 19508
rect 8444 19456 8450 19508
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10870 19496 10876 19508
rect 9732 19468 10876 19496
rect 9732 19456 9738 19468
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11054 19456 11060 19508
rect 11112 19496 11118 19508
rect 11517 19499 11575 19505
rect 11517 19496 11529 19499
rect 11112 19468 11529 19496
rect 11112 19456 11118 19468
rect 11517 19465 11529 19468
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 13814 19496 13820 19508
rect 11664 19468 13820 19496
rect 11664 19456 11670 19468
rect 5902 19428 5908 19440
rect 1964 19400 4016 19428
rect 4080 19400 5908 19428
rect 1964 19369 1992 19400
rect 4080 19369 4108 19400
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 8294 19428 8300 19440
rect 6012 19400 8300 19428
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5442 19360 5448 19372
rect 4847 19332 5448 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 6012 19369 6040 19400
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 11072 19428 11100 19456
rect 10534 19400 11100 19428
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19329 6055 19363
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 5997 19323 6055 19329
rect 6656 19332 7297 19360
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1912 19264 2237 19292
rect 1912 19252 1918 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 2924 19264 4537 19292
rect 2924 19252 2930 19264
rect 4525 19261 4537 19264
rect 4571 19261 4583 19295
rect 4525 19255 4583 19261
rect 6457 19295 6515 19301
rect 6457 19261 6469 19295
rect 6503 19292 6515 19295
rect 6546 19292 6552 19304
rect 6503 19264 6552 19292
rect 6503 19261 6515 19264
rect 6457 19255 6515 19261
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 6656 19301 6684 19332
rect 7285 19329 7297 19332
rect 7331 19360 7343 19363
rect 7742 19360 7748 19372
rect 7331 19332 7748 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8938 19360 8944 19372
rect 8619 19332 8944 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 12544 19360 12572 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 14056 19468 14473 19496
rect 14056 19456 14062 19468
rect 14461 19465 14473 19468
rect 14507 19496 14519 19499
rect 14642 19496 14648 19508
rect 14507 19468 14648 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 14918 19456 14924 19508
rect 14976 19456 14982 19508
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 15562 19496 15568 19508
rect 15335 19468 15568 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 17034 19456 17040 19508
rect 17092 19456 17098 19508
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 18785 19499 18843 19505
rect 18785 19496 18797 19499
rect 18196 19468 18797 19496
rect 18196 19456 18202 19468
rect 18785 19465 18797 19468
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19659 19468 20453 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 20990 19496 20996 19508
rect 20947 19468 20996 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21232 19468 22017 19496
rect 21232 19456 21238 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22370 19456 22376 19508
rect 22428 19456 22434 19508
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 25130 19496 25136 19508
rect 25087 19468 25136 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 25130 19456 25136 19468
rect 25188 19496 25194 19508
rect 25314 19496 25320 19508
rect 25188 19468 25320 19496
rect 25188 19456 25194 19468
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 13262 19428 13268 19440
rect 12676 19400 13268 19428
rect 12676 19388 12682 19400
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 14274 19388 14280 19440
rect 14332 19428 14338 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14332 19400 15393 19428
rect 14332 19388 14338 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 16574 19428 16580 19440
rect 15381 19391 15439 19397
rect 16316 19400 16580 19428
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12544 19332 12725 19360
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 14458 19360 14464 19372
rect 14122 19332 14464 19360
rect 12713 19323 12771 19329
rect 14458 19320 14464 19332
rect 14516 19360 14522 19372
rect 15194 19360 15200 19372
rect 14516 19332 15200 19360
rect 14516 19320 14522 19332
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 16316 19369 16344 19400
rect 16574 19388 16580 19400
rect 16632 19388 16638 19440
rect 17052 19428 17080 19456
rect 17052 19400 17802 19428
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 19705 19431 19763 19437
rect 19705 19428 19717 19431
rect 19484 19400 19717 19428
rect 19484 19388 19490 19400
rect 19705 19397 19717 19400
rect 19751 19397 19763 19431
rect 19705 19391 19763 19397
rect 20809 19431 20867 19437
rect 20809 19397 20821 19431
rect 20855 19428 20867 19431
rect 23566 19428 23572 19440
rect 20855 19400 23572 19428
rect 20855 19397 20867 19400
rect 20809 19391 20867 19397
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17026 19363 17084 19369
rect 17026 19360 17038 19363
rect 16540 19332 17038 19360
rect 16540 19320 16546 19332
rect 17026 19329 17038 19332
rect 17072 19329 17084 19363
rect 21266 19360 21272 19372
rect 17026 19323 17084 19329
rect 19260 19332 21272 19360
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 6730 19252 6736 19304
rect 6788 19252 6794 19304
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 10778 19292 10784 19304
rect 9355 19264 10784 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 11790 19252 11796 19304
rect 11848 19252 11854 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 15102 19292 15108 19304
rect 13035 19264 15108 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16390 19252 16396 19304
rect 16448 19252 16454 19304
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 17678 19292 17684 19304
rect 17368 19264 17684 19292
rect 17368 19252 17374 19264
rect 17678 19252 17684 19264
rect 17736 19292 17742 19304
rect 17736 19264 18460 19292
rect 17736 19252 17742 19264
rect 6914 19184 6920 19236
rect 6972 19224 6978 19236
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 6972 19196 7757 19224
rect 6972 19184 6978 19196
rect 7745 19193 7757 19196
rect 7791 19193 7803 19227
rect 11808 19224 11836 19252
rect 7745 19187 7803 19193
rect 10336 19196 11836 19224
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 8570 19156 8576 19168
rect 3384 19128 8576 19156
rect 3384 19116 3390 19128
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9398 19116 9404 19168
rect 9456 19156 9462 19168
rect 10336 19156 10364 19196
rect 15654 19184 15660 19236
rect 15712 19224 15718 19236
rect 16408 19224 16436 19252
rect 16669 19227 16727 19233
rect 16669 19224 16681 19227
rect 15712 19196 16681 19224
rect 15712 19184 15718 19196
rect 16669 19193 16681 19196
rect 16715 19193 16727 19227
rect 16669 19187 16727 19193
rect 9456 19128 10364 19156
rect 9456 19116 9462 19128
rect 10778 19116 10784 19168
rect 10836 19116 10842 19168
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19156 11391 19159
rect 11422 19156 11428 19168
rect 11379 19128 11428 19156
rect 11379 19125 11391 19128
rect 11333 19119 11391 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 11790 19116 11796 19168
rect 11848 19116 11854 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13630 19156 13636 19168
rect 12492 19128 13636 19156
rect 12492 19116 12498 19128
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14734 19156 14740 19168
rect 14516 19128 14740 19156
rect 14516 19116 14522 19128
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16390 19156 16396 19168
rect 16163 19128 16396 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 18432 19156 18460 19264
rect 19260 19233 19288 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21358 19320 21364 19372
rect 21416 19320 21422 19372
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20404 19264 21005 19292
rect 20404 19252 20410 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19193 19303 19227
rect 19245 19187 19303 19193
rect 21082 19184 21088 19236
rect 21140 19224 21146 19236
rect 21376 19224 21404 19320
rect 22002 19252 22008 19304
rect 22060 19292 22066 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22060 19264 22477 19292
rect 22060 19252 22066 19264
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 25222 19292 25228 19304
rect 23615 19264 25228 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 21453 19227 21511 19233
rect 21453 19224 21465 19227
rect 21140 19196 21465 19224
rect 21140 19184 21146 19196
rect 21453 19193 21465 19196
rect 21499 19193 21511 19227
rect 21453 19187 21511 19193
rect 21726 19184 21732 19236
rect 21784 19224 21790 19236
rect 22572 19224 22600 19255
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 21784 19196 22600 19224
rect 21784 19184 21790 19196
rect 24670 19184 24676 19236
rect 24728 19224 24734 19236
rect 25038 19224 25044 19236
rect 24728 19196 25044 19224
rect 24728 19184 24734 19196
rect 25038 19184 25044 19196
rect 25096 19224 25102 19236
rect 25317 19227 25375 19233
rect 25317 19224 25329 19227
rect 25096 19196 25329 19224
rect 25096 19184 25102 19196
rect 25317 19193 25329 19196
rect 25363 19193 25375 19227
rect 25317 19187 25375 19193
rect 19702 19156 19708 19168
rect 18432 19128 19708 19156
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20990 19156 20996 19168
rect 20404 19128 20996 19156
rect 20404 19116 20410 19128
rect 20990 19116 20996 19128
rect 21048 19156 21054 19168
rect 22186 19156 22192 19168
rect 21048 19128 22192 19156
rect 21048 19116 21054 19128
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18952 2007 18955
rect 2406 18952 2412 18964
rect 1995 18924 2412 18952
rect 1995 18921 2007 18924
rect 1949 18915 2007 18921
rect 2406 18912 2412 18924
rect 2464 18912 2470 18964
rect 3602 18952 3608 18964
rect 2746 18924 3608 18952
rect 2593 18887 2651 18893
rect 2593 18853 2605 18887
rect 2639 18884 2651 18887
rect 2746 18884 2774 18924
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 3694 18912 3700 18964
rect 3752 18952 3758 18964
rect 3881 18955 3939 18961
rect 3881 18952 3893 18955
rect 3752 18924 3893 18952
rect 3752 18912 3758 18924
rect 3881 18921 3893 18924
rect 3927 18952 3939 18955
rect 5534 18952 5540 18964
rect 3927 18924 5540 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 5902 18912 5908 18964
rect 5960 18952 5966 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 5960 18924 8401 18952
rect 5960 18912 5966 18924
rect 8389 18921 8401 18924
rect 8435 18921 8447 18955
rect 8389 18915 8447 18921
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 10686 18952 10692 18964
rect 8628 18924 10692 18952
rect 8628 18912 8634 18924
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 14182 18952 14188 18964
rect 12575 18924 14188 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 14182 18912 14188 18924
rect 14240 18912 14246 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 23198 18952 23204 18964
rect 14384 18924 23204 18952
rect 9217 18887 9275 18893
rect 9217 18884 9229 18887
rect 2639 18856 2774 18884
rect 3436 18856 9229 18884
rect 2639 18853 2651 18856
rect 2593 18847 2651 18853
rect 2130 18708 2136 18760
rect 2188 18708 2194 18760
rect 3436 18757 3464 18856
rect 9217 18853 9229 18856
rect 9263 18853 9275 18887
rect 12989 18887 13047 18893
rect 12989 18884 13001 18887
rect 9217 18847 9275 18853
rect 9416 18856 13001 18884
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 5813 18819 5871 18825
rect 4111 18788 5120 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 5092 18760 5120 18788
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 6546 18816 6552 18828
rect 5859 18788 6552 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7190 18816 7196 18828
rect 7147 18788 7196 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 7377 18819 7435 18825
rect 7377 18785 7389 18819
rect 7423 18816 7435 18819
rect 7558 18816 7564 18828
rect 7423 18788 7564 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 7834 18776 7840 18828
rect 7892 18816 7898 18828
rect 9416 18816 9444 18856
rect 12989 18853 13001 18856
rect 13035 18853 13047 18887
rect 14384 18884 14412 18924
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 25038 18912 25044 18964
rect 25096 18912 25102 18964
rect 14918 18884 14924 18896
rect 12989 18847 13047 18853
rect 13464 18856 14412 18884
rect 14844 18856 14924 18884
rect 7892 18788 9444 18816
rect 7892 18776 7898 18788
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9548 18788 9781 18816
rect 9548 18776 9554 18788
rect 9769 18785 9781 18788
rect 9815 18785 9827 18819
rect 9769 18779 9827 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 13464 18816 13492 18856
rect 11020 18788 13492 18816
rect 11020 18776 11026 18788
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 14734 18816 14740 18828
rect 13740 18788 14740 18816
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 4706 18748 4712 18760
rect 4203 18720 4712 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 2792 18680 2820 18711
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5132 18720 5365 18748
rect 5132 18708 5138 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18748 6147 18751
rect 6178 18748 6184 18760
rect 6135 18720 6184 18748
rect 6135 18717 6147 18720
rect 6089 18711 6147 18717
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 4246 18680 4252 18692
rect 2792 18652 4252 18680
rect 4246 18640 4252 18652
rect 4304 18640 4310 18692
rect 5718 18680 5724 18692
rect 4540 18652 5724 18680
rect 3234 18572 3240 18624
rect 3292 18572 3298 18624
rect 4540 18621 4568 18652
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 8588 18680 8616 18711
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9180 18720 9597 18748
rect 9180 18708 9186 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11790 18748 11796 18760
rect 10459 18720 11796 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 13740 18748 13768 18788
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 14844 18825 14872 18856
rect 14918 18844 14924 18856
rect 14976 18844 14982 18896
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17862 18884 17868 18896
rect 17267 18856 17868 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 18049 18887 18107 18893
rect 18049 18853 18061 18887
rect 18095 18884 18107 18887
rect 19058 18884 19064 18896
rect 18095 18856 19064 18884
rect 18095 18853 18107 18856
rect 18049 18847 18107 18853
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 21634 18844 21640 18896
rect 21692 18844 21698 18896
rect 22557 18887 22615 18893
rect 22557 18853 22569 18887
rect 22603 18884 22615 18887
rect 25056 18884 25084 18912
rect 22603 18856 25084 18884
rect 22603 18853 22615 18856
rect 22557 18847 22615 18853
rect 14829 18819 14887 18825
rect 14829 18785 14841 18819
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 17678 18816 17684 18828
rect 15068 18788 17684 18816
rect 15068 18776 15074 18788
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 18380 18788 18613 18816
rect 18380 18776 18386 18788
rect 18601 18785 18613 18788
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 21652 18816 21680 18844
rect 20671 18788 21680 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22520 18788 23121 18816
rect 22520 18776 22526 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 25041 18819 25099 18825
rect 25041 18816 25053 18819
rect 23109 18779 23167 18785
rect 23216 18788 25053 18816
rect 12406 18720 13768 18748
rect 9306 18680 9312 18692
rect 8588 18652 9312 18680
rect 9306 18640 9312 18652
rect 9364 18640 9370 18692
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 12406 18680 12434 18720
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14918 18748 14924 18760
rect 13872 18720 14924 18748
rect 13872 18708 13878 18720
rect 14918 18708 14924 18720
rect 14976 18748 14982 18760
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 14976 18720 15485 18748
rect 14976 18708 14982 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18874 18748 18880 18760
rect 18463 18720 18880 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 22094 18748 22100 18760
rect 20349 18711 20407 18717
rect 21836 18720 22100 18748
rect 9723 18652 12434 18680
rect 13357 18683 13415 18689
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13722 18680 13728 18692
rect 13403 18652 13728 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 14645 18683 14703 18689
rect 14645 18649 14657 18683
rect 14691 18680 14703 18683
rect 15010 18680 15016 18692
rect 14691 18652 15016 18680
rect 14691 18649 14703 18652
rect 14645 18643 14703 18649
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16298 18640 16304 18692
rect 16356 18640 16362 18692
rect 18322 18640 18328 18692
rect 18380 18680 18386 18692
rect 19242 18680 19248 18692
rect 18380 18652 19248 18680
rect 18380 18640 18386 18652
rect 19242 18640 19248 18652
rect 19300 18680 19306 18692
rect 20364 18680 20392 18711
rect 21082 18680 21088 18692
rect 19300 18652 20392 18680
rect 21008 18652 21088 18680
rect 19300 18640 19306 18652
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18581 4583 18615
rect 4525 18575 4583 18581
rect 5169 18615 5227 18621
rect 5169 18581 5181 18615
rect 5215 18612 5227 18615
rect 8202 18612 8208 18624
rect 5215 18584 8208 18612
rect 5215 18581 5227 18584
rect 5169 18575 5227 18581
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 10502 18612 10508 18624
rect 8628 18584 10508 18612
rect 8628 18572 8634 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 13446 18572 13452 18624
rect 13504 18572 13510 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 14737 18615 14795 18621
rect 14737 18612 14749 18615
rect 13596 18584 14749 18612
rect 13596 18572 13602 18584
rect 14737 18581 14749 18584
rect 14783 18612 14795 18615
rect 15654 18612 15660 18624
rect 14783 18584 15660 18612
rect 14783 18581 14795 18584
rect 14737 18575 14795 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17184 18584 17509 18612
rect 17184 18572 17190 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 17678 18572 17684 18624
rect 17736 18572 17742 18624
rect 18509 18615 18567 18621
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 19429 18615 19487 18621
rect 19429 18612 19441 18615
rect 18555 18584 19441 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19429 18581 19441 18584
rect 19475 18581 19487 18615
rect 19429 18575 19487 18581
rect 19702 18572 19708 18624
rect 19760 18612 19766 18624
rect 19889 18615 19947 18621
rect 19889 18612 19901 18615
rect 19760 18584 19901 18612
rect 19760 18572 19766 18584
rect 19889 18581 19901 18584
rect 19935 18581 19947 18615
rect 21008 18612 21036 18652
rect 21082 18640 21088 18652
rect 21140 18640 21146 18692
rect 21836 18680 21864 18720
rect 22094 18708 22100 18720
rect 22152 18708 22158 18760
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 22244 18720 22324 18748
rect 22244 18708 22250 18720
rect 21836 18666 21956 18680
rect 21850 18652 21956 18666
rect 21928 18612 21956 18652
rect 21008 18584 21956 18612
rect 22097 18615 22155 18621
rect 19889 18575 19947 18581
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22186 18612 22192 18624
rect 22143 18584 22192 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 22296 18612 22324 18720
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22888 18720 23029 18748
rect 22888 18708 22894 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23216 18748 23244 18788
rect 25041 18785 25053 18788
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 23017 18711 23075 18717
rect 23124 18720 23244 18748
rect 23845 18751 23903 18757
rect 22554 18640 22560 18692
rect 22612 18680 22618 18692
rect 23124 18680 23152 18720
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 24118 18748 24124 18760
rect 23891 18720 24124 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 22612 18652 23152 18680
rect 22612 18640 22618 18652
rect 22830 18612 22836 18624
rect 22296 18584 22836 18612
rect 22830 18572 22836 18584
rect 22888 18612 22894 18624
rect 22925 18615 22983 18621
rect 22925 18612 22937 18615
rect 22888 18584 22937 18612
rect 22888 18572 22894 18584
rect 22925 18581 22937 18584
rect 22971 18581 22983 18615
rect 22925 18575 22983 18581
rect 23014 18572 23020 18624
rect 23072 18612 23078 18624
rect 23860 18612 23888 18711
rect 24118 18708 24124 18720
rect 24176 18708 24182 18760
rect 24029 18683 24087 18689
rect 24029 18649 24041 18683
rect 24075 18680 24087 18683
rect 25682 18680 25688 18692
rect 24075 18652 25688 18680
rect 24075 18649 24087 18652
rect 24029 18643 24087 18649
rect 25682 18640 25688 18652
rect 25740 18640 25746 18692
rect 23072 18584 23888 18612
rect 23072 18572 23078 18584
rect 24578 18572 24584 18624
rect 24636 18572 24642 18624
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 2130 18368 2136 18420
rect 2188 18408 2194 18420
rect 2225 18411 2283 18417
rect 2225 18408 2237 18411
rect 2188 18380 2237 18408
rect 2188 18368 2194 18380
rect 2225 18377 2237 18380
rect 2271 18377 2283 18411
rect 2225 18371 2283 18377
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 2866 18408 2872 18420
rect 2639 18380 2872 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3237 18411 3295 18417
rect 3237 18377 3249 18411
rect 3283 18408 3295 18411
rect 4062 18408 4068 18420
rect 3283 18380 4068 18408
rect 3283 18377 3295 18380
rect 3237 18371 3295 18377
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4522 18368 4528 18420
rect 4580 18368 4586 18420
rect 5810 18368 5816 18420
rect 5868 18368 5874 18420
rect 7006 18408 7012 18420
rect 5920 18380 7012 18408
rect 5920 18340 5948 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 7650 18368 7656 18420
rect 7708 18368 7714 18420
rect 8294 18368 8300 18420
rect 8352 18368 8358 18420
rect 10778 18408 10784 18420
rect 9232 18380 10784 18408
rect 4724 18312 5948 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 1811 18244 2145 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2133 18241 2145 18244
rect 2179 18272 2191 18275
rect 2498 18272 2504 18284
rect 2179 18244 2504 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18272 2835 18275
rect 3326 18272 3332 18284
rect 2823 18244 3332 18272
rect 2823 18241 2835 18244
rect 2777 18235 2835 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18272 3479 18275
rect 3694 18272 3700 18284
rect 3467 18244 3700 18272
rect 3467 18241 3479 18244
rect 3421 18235 3479 18241
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 4724 18281 4752 18312
rect 6730 18300 6736 18352
rect 6788 18340 6794 18352
rect 9122 18340 9128 18352
rect 6788 18312 7236 18340
rect 6788 18300 6794 18312
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 5350 18232 5356 18284
rect 5408 18232 5414 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6914 18272 6920 18284
rect 6043 18244 6920 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7208 18281 7236 18312
rect 7852 18312 9128 18340
rect 7852 18284 7880 18312
rect 9122 18300 9128 18312
rect 9180 18300 9186 18352
rect 9232 18349 9260 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12124 18380 12173 18408
rect 12124 18368 12130 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13872 18380 14289 18408
rect 13872 18368 13878 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14792 18380 15209 18408
rect 14792 18368 14798 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15654 18368 15660 18420
rect 15712 18368 15718 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 18506 18408 18512 18420
rect 16347 18380 18512 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 9217 18343 9275 18349
rect 9217 18309 9229 18343
rect 9263 18309 9275 18343
rect 10870 18340 10876 18352
rect 10442 18312 10876 18340
rect 9217 18303 9275 18309
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 10962 18300 10968 18352
rect 11020 18340 11026 18352
rect 11241 18343 11299 18349
rect 11241 18340 11253 18343
rect 11020 18312 11253 18340
rect 11020 18300 11026 18312
rect 11241 18309 11253 18312
rect 11287 18309 11299 18343
rect 11241 18303 11299 18309
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 11848 18312 13001 18340
rect 11848 18300 11854 18312
rect 12989 18309 13001 18312
rect 13035 18340 13047 18343
rect 16316 18340 16344 18371
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 20346 18408 20352 18420
rect 19659 18380 20352 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 23106 18408 23112 18420
rect 21192 18380 23112 18408
rect 13035 18312 16344 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 17402 18300 17408 18352
rect 17460 18300 17466 18352
rect 17954 18300 17960 18352
rect 18012 18340 18018 18352
rect 20530 18340 20536 18352
rect 18012 18312 20536 18340
rect 18012 18300 18018 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 20627 18312 20852 18340
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3835 18176 3893 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3881 18173 3893 18176
rect 3927 18204 3939 18207
rect 5534 18204 5540 18216
rect 3927 18176 5540 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 6549 18207 6607 18213
rect 6549 18173 6561 18207
rect 6595 18204 6607 18207
rect 8754 18204 8760 18216
rect 6595 18176 8760 18204
rect 6595 18173 6607 18176
rect 6549 18167 6607 18173
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 8956 18204 8984 18235
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 10560 18244 15577 18272
rect 10560 18232 10566 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16393 18275 16451 18281
rect 16393 18272 16405 18275
rect 16356 18244 16405 18272
rect 16356 18232 16362 18244
rect 16393 18241 16405 18244
rect 16439 18272 16451 18275
rect 17126 18272 17132 18284
rect 16439 18244 17132 18272
rect 16439 18241 16451 18244
rect 16393 18235 16451 18241
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 17420 18272 17448 18300
rect 18230 18272 18236 18284
rect 17420 18244 18236 18272
rect 18230 18232 18236 18244
rect 18288 18272 18294 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18288 18244 18429 18272
rect 18288 18232 18294 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 20438 18272 20444 18284
rect 18417 18235 18475 18241
rect 18616 18244 20444 18272
rect 8956 18176 9076 18204
rect 1581 18139 1639 18145
rect 1581 18105 1593 18139
rect 1627 18136 1639 18139
rect 2774 18136 2780 18148
rect 1627 18108 2780 18136
rect 1627 18105 1639 18108
rect 1581 18099 1639 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 3160 18108 5181 18136
rect 2682 18028 2688 18080
rect 2740 18068 2746 18080
rect 3160 18068 3188 18108
rect 5169 18105 5181 18108
rect 5215 18105 5227 18139
rect 5169 18099 5227 18105
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 8386 18136 8392 18148
rect 7055 18108 8392 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 9048 18080 9076 18176
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 12253 18207 12311 18213
rect 9364 18176 11836 18204
rect 9364 18164 9370 18176
rect 11808 18145 11836 18176
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11793 18139 11851 18145
rect 10735 18108 11744 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 2740 18040 3188 18068
rect 2740 18028 2746 18040
rect 3234 18028 3240 18080
rect 3292 18068 3298 18080
rect 6546 18068 6552 18080
rect 3292 18040 6552 18068
rect 3292 18028 3298 18040
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 6733 18071 6791 18077
rect 6733 18037 6745 18071
rect 6779 18068 6791 18071
rect 7834 18068 7840 18080
rect 6779 18040 7840 18068
rect 6779 18037 6791 18040
rect 6733 18031 6791 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 9030 18028 9036 18080
rect 9088 18028 9094 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10704 18068 10732 18099
rect 9824 18040 10732 18068
rect 9824 18028 9830 18040
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 10928 18040 11161 18068
rect 10928 18028 10934 18040
rect 11149 18037 11161 18040
rect 11195 18068 11207 18071
rect 11606 18068 11612 18080
rect 11195 18040 11612 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 11716 18068 11744 18108
rect 11793 18105 11805 18139
rect 11839 18105 11851 18139
rect 12268 18136 12296 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 12492 18176 15761 18204
rect 12492 18164 12498 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 17313 18207 17371 18213
rect 17313 18204 17325 18207
rect 16264 18176 17325 18204
rect 16264 18164 16270 18176
rect 17313 18173 17325 18176
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 17494 18164 17500 18216
rect 17552 18204 17558 18216
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 17552 18176 18521 18204
rect 17552 18164 17558 18176
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 12268 18108 13860 18136
rect 11793 18099 11851 18105
rect 12434 18068 12440 18080
rect 11716 18040 12440 18068
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 13832 18068 13860 18108
rect 14660 18108 16865 18136
rect 14660 18068 14688 18108
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 18616 18136 18644 18244
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 18690 18164 18696 18216
rect 18748 18164 18754 18216
rect 19518 18164 19524 18216
rect 19576 18204 19582 18216
rect 19705 18207 19763 18213
rect 19705 18204 19717 18207
rect 19576 18176 19717 18204
rect 19576 18164 19582 18176
rect 19705 18173 19717 18176
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 19794 18164 19800 18216
rect 19852 18164 19858 18216
rect 20627 18204 20655 18312
rect 20824 18281 20852 18312
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 21192 18340 21220 18380
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 24118 18368 24124 18420
rect 24176 18408 24182 18420
rect 24213 18411 24271 18417
rect 24213 18408 24225 18411
rect 24176 18380 24225 18408
rect 24176 18368 24182 18380
rect 24213 18377 24225 18380
rect 24259 18408 24271 18411
rect 24670 18408 24676 18420
rect 24259 18380 24676 18408
rect 24259 18377 24271 18380
rect 24213 18371 24271 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 21048 18312 21220 18340
rect 21048 18300 21054 18312
rect 21450 18300 21456 18352
rect 21508 18340 21514 18352
rect 22005 18343 22063 18349
rect 22005 18340 22017 18343
rect 21508 18312 22017 18340
rect 21508 18300 21514 18312
rect 22005 18309 22017 18312
rect 22051 18340 22063 18343
rect 24029 18343 24087 18349
rect 24029 18340 24041 18343
rect 22051 18312 24041 18340
rect 22051 18309 22063 18312
rect 22005 18303 22063 18309
rect 24029 18309 24041 18312
rect 24075 18309 24087 18343
rect 24029 18303 24087 18309
rect 24302 18300 24308 18352
rect 24360 18340 24366 18352
rect 24489 18343 24547 18349
rect 24489 18340 24501 18343
rect 24360 18312 24501 18340
rect 24360 18300 24366 18312
rect 24489 18309 24501 18312
rect 24535 18340 24547 18343
rect 24949 18343 25007 18349
rect 24949 18340 24961 18343
rect 24535 18312 24961 18340
rect 24535 18309 24547 18312
rect 24489 18303 24547 18309
rect 24949 18309 24961 18312
rect 24995 18340 25007 18343
rect 25866 18340 25872 18352
rect 24995 18312 25872 18340
rect 24995 18309 25007 18312
rect 24949 18303 25007 18309
rect 25866 18300 25872 18312
rect 25924 18300 25930 18352
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18272 20867 18275
rect 21818 18272 21824 18284
rect 20855 18244 21824 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 20364 18176 20655 18204
rect 20364 18136 20392 18176
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 20901 18207 20959 18213
rect 20901 18204 20913 18207
rect 20772 18176 20913 18204
rect 20772 18164 20778 18176
rect 20901 18173 20913 18176
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 20990 18164 20996 18216
rect 21048 18164 21054 18216
rect 21266 18164 21272 18216
rect 21324 18204 21330 18216
rect 24670 18204 24676 18216
rect 21324 18176 24676 18204
rect 21324 18164 21330 18176
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24780 18176 25053 18204
rect 16853 18099 16911 18105
rect 16960 18108 18644 18136
rect 19168 18108 20392 18136
rect 20441 18139 20499 18145
rect 13832 18040 14688 18068
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 16960 18068 16988 18108
rect 14792 18040 16988 18068
rect 14792 18028 14798 18040
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17552 18040 18061 18068
rect 17552 18028 17558 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 18230 18028 18236 18080
rect 18288 18068 18294 18080
rect 19168 18068 19196 18108
rect 20441 18105 20453 18139
rect 20487 18136 20499 18139
rect 20530 18136 20536 18148
rect 20487 18108 20536 18136
rect 20487 18105 20499 18108
rect 20441 18099 20499 18105
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 21453 18139 21511 18145
rect 21453 18136 21465 18139
rect 20995 18108 21465 18136
rect 18288 18040 19196 18068
rect 18288 18028 18294 18040
rect 19242 18028 19248 18080
rect 19300 18028 19306 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20995 18068 21023 18108
rect 21453 18105 21465 18108
rect 21499 18105 21511 18139
rect 21453 18099 21511 18105
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 22094 18136 22100 18148
rect 21876 18108 22100 18136
rect 21876 18096 21882 18108
rect 22094 18096 22100 18108
rect 22152 18096 22158 18148
rect 23382 18096 23388 18148
rect 23440 18136 23446 18148
rect 24581 18139 24639 18145
rect 24581 18136 24593 18139
rect 23440 18108 24593 18136
rect 23440 18096 23446 18108
rect 24581 18105 24593 18108
rect 24627 18105 24639 18139
rect 24581 18099 24639 18105
rect 20772 18040 21023 18068
rect 20772 18028 20778 18040
rect 22554 18028 22560 18080
rect 22612 18068 22618 18080
rect 24780 18068 24808 18176
rect 25041 18173 25053 18176
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25498 18204 25504 18216
rect 25271 18176 25504 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 22612 18040 24808 18068
rect 22612 18028 22618 18040
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 2777 17867 2835 17873
rect 2777 17864 2789 17867
rect 1504 17836 2789 17864
rect 1504 17660 1532 17836
rect 2777 17833 2789 17836
rect 2823 17864 2835 17867
rect 4982 17864 4988 17876
rect 2823 17836 4988 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 4982 17824 4988 17836
rect 5040 17824 5046 17876
rect 6454 17824 6460 17876
rect 6512 17824 6518 17876
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 7064 17836 7113 17864
rect 7064 17824 7070 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7101 17827 7159 17833
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7248 17836 7757 17864
rect 7248 17824 7254 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 7745 17827 7803 17833
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 8754 17864 8760 17876
rect 7892 17836 8760 17864
rect 7892 17824 7898 17836
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 11238 17864 11244 17876
rect 9364 17836 11244 17864
rect 9364 17824 9370 17836
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 13354 17864 13360 17876
rect 11348 17836 13360 17864
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 8294 17796 8300 17808
rect 1627 17768 8300 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 11054 17756 11060 17808
rect 11112 17796 11118 17808
rect 11348 17796 11376 17836
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 13504 17836 17141 17864
rect 13504 17824 13510 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 17129 17827 17187 17833
rect 18233 17867 18291 17873
rect 18233 17833 18245 17867
rect 18279 17864 18291 17867
rect 18874 17864 18880 17876
rect 18279 17836 18880 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18874 17824 18880 17836
rect 18932 17864 18938 17876
rect 19150 17864 19156 17876
rect 18932 17836 19156 17864
rect 18932 17824 18938 17836
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19886 17824 19892 17876
rect 19944 17864 19950 17876
rect 20714 17864 20720 17876
rect 19944 17836 20720 17864
rect 19944 17824 19950 17836
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 20980 17867 21038 17873
rect 20980 17833 20992 17867
rect 21026 17864 21038 17867
rect 22186 17864 22192 17876
rect 21026 17836 22192 17864
rect 21026 17833 21038 17836
rect 20980 17827 21038 17833
rect 22186 17824 22192 17836
rect 22244 17824 22250 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22646 17864 22652 17876
rect 22511 17836 22652 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 24581 17867 24639 17873
rect 22888 17836 23428 17864
rect 22888 17824 22894 17836
rect 11112 17768 11376 17796
rect 16669 17799 16727 17805
rect 11112 17756 11118 17768
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 17310 17796 17316 17808
rect 16715 17768 17316 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 23293 17799 23351 17805
rect 23293 17765 23305 17799
rect 23339 17765 23351 17799
rect 23400 17796 23428 17836
rect 24581 17833 24593 17867
rect 24627 17864 24639 17867
rect 24854 17864 24860 17876
rect 24627 17836 24860 17864
rect 24627 17833 24639 17836
rect 24581 17827 24639 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 23400 17768 25084 17796
rect 23293 17759 23351 17765
rect 2222 17688 2228 17740
rect 2280 17688 2286 17740
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17728 5227 17731
rect 5258 17728 5264 17740
rect 5215 17700 5264 17728
rect 5215 17697 5227 17700
rect 5169 17691 5227 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17728 5503 17731
rect 5994 17728 6000 17740
rect 5491 17700 6000 17728
rect 5491 17697 5503 17700
rect 5445 17691 5503 17697
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 6362 17688 6368 17740
rect 6420 17728 6426 17740
rect 6420 17700 7972 17728
rect 6420 17688 6426 17700
rect 1765 17663 1823 17669
rect 1765 17660 1777 17663
rect 1504 17632 1777 17660
rect 1765 17629 1777 17632
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 4249 17663 4307 17669
rect 3467 17632 3924 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3896 17536 3924 17632
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4706 17660 4712 17672
rect 4295 17632 4712 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17660 7343 17663
rect 7834 17660 7840 17672
rect 7331 17632 7840 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 7944 17669 7972 17700
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9088 17700 9720 17728
rect 9088 17688 9094 17700
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8619 17632 9260 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8478 17592 8484 17604
rect 4540 17564 8484 17592
rect 3237 17527 3295 17533
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 3326 17524 3332 17536
rect 3283 17496 3332 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 3326 17484 3332 17496
rect 3384 17484 3390 17536
rect 3878 17484 3884 17536
rect 3936 17484 3942 17536
rect 4540 17533 4568 17564
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17493 4583 17527
rect 4525 17487 4583 17493
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 7558 17524 7564 17536
rect 4672 17496 7564 17524
rect 4672 17484 4678 17496
rect 7558 17484 7564 17496
rect 7616 17484 7622 17536
rect 8386 17484 8392 17536
rect 8444 17484 8450 17536
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 9232 17524 9260 17632
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 9692 17660 9720 17700
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11756 17700 11989 17728
rect 11756 17688 11762 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12618 17728 12624 17740
rect 12299 17700 12624 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13780 17700 14289 17728
rect 13780 17688 13786 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15654 17688 15660 17740
rect 15712 17728 15718 17740
rect 15838 17728 15844 17740
rect 15712 17700 15844 17728
rect 15712 17688 15718 17700
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 16390 17688 16396 17740
rect 16448 17688 16454 17740
rect 16758 17688 16764 17740
rect 16816 17728 16822 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16816 17700 17693 17728
rect 16816 17688 16822 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 18524 17700 19748 17728
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9692 17632 9781 17660
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16408 17660 16436 17688
rect 18524 17660 18552 17700
rect 16408 17632 18552 17660
rect 18598 17620 18604 17672
rect 18656 17620 18662 17672
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 10042 17592 10048 17604
rect 9548 17564 10048 17592
rect 9548 17552 9554 17564
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 11606 17592 11612 17604
rect 11270 17564 11612 17592
rect 11606 17552 11612 17564
rect 11664 17592 11670 17604
rect 12710 17592 12716 17604
rect 11664 17564 12716 17592
rect 11664 17552 11670 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 15194 17592 15200 17604
rect 13688 17564 15200 17592
rect 13688 17552 13694 17564
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 17402 17592 17408 17604
rect 16500 17564 17408 17592
rect 11422 17524 11428 17536
rect 9232 17496 11428 17524
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 11974 17524 11980 17536
rect 11563 17496 11980 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 12584 17496 13737 17524
rect 12584 17484 12590 17496
rect 13725 17493 13737 17496
rect 13771 17524 13783 17527
rect 16500 17524 16528 17564
rect 17402 17552 17408 17564
rect 17460 17552 17466 17604
rect 17497 17595 17555 17601
rect 17497 17561 17509 17595
rect 17543 17592 17555 17595
rect 18616 17592 18644 17620
rect 17543 17564 18828 17592
rect 17543 17561 17555 17564
rect 17497 17555 17555 17561
rect 18800 17536 18828 17564
rect 13771 17496 16528 17524
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 16632 17496 17601 17524
rect 16632 17484 16638 17496
rect 17589 17493 17601 17496
rect 17635 17524 17647 17527
rect 17678 17524 17684 17536
rect 17635 17496 17684 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19610 17524 19616 17536
rect 19475 17496 19616 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 19720 17524 19748 17700
rect 19886 17688 19892 17740
rect 19944 17688 19950 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20346 17728 20352 17740
rect 20119 17700 20352 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 22554 17728 22560 17740
rect 20763 17700 22560 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 22554 17688 22560 17700
rect 22612 17728 22618 17740
rect 23198 17728 23204 17740
rect 22612 17700 23204 17728
rect 22612 17688 22618 17700
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 23308 17660 23336 17759
rect 23934 17688 23940 17740
rect 23992 17728 23998 17740
rect 24302 17728 24308 17740
rect 23992 17700 24308 17728
rect 23992 17688 23998 17700
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 25056 17737 25084 17768
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17728 25283 17731
rect 25774 17728 25780 17740
rect 25271 17700 25780 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 23382 17660 23388 17672
rect 23308 17632 23388 17660
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 23658 17620 23664 17672
rect 23716 17620 23722 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24486 17660 24492 17672
rect 23799 17632 24492 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24486 17620 24492 17632
rect 24544 17620 24550 17672
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 19843 17564 20944 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 20714 17524 20720 17536
rect 19720 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 20916 17524 20944 17564
rect 21266 17552 21272 17604
rect 21324 17592 21330 17604
rect 23566 17592 23572 17604
rect 21324 17564 21482 17592
rect 22664 17564 23572 17592
rect 21324 17552 21330 17564
rect 22664 17524 22692 17564
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 20916 17496 22692 17524
rect 22833 17527 22891 17533
rect 22833 17493 22845 17527
rect 22879 17524 22891 17527
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22879 17496 23029 17524
rect 22879 17493 22891 17496
rect 22833 17487 22891 17493
rect 23017 17493 23029 17496
rect 23063 17524 23075 17527
rect 24118 17524 24124 17536
rect 23063 17496 24124 17524
rect 23063 17493 23075 17496
rect 23017 17487 23075 17493
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24486 17524 24492 17536
rect 24268 17496 24492 17524
rect 24268 17484 24274 17496
rect 24486 17484 24492 17496
rect 24544 17484 24550 17536
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24636 17496 24961 17524
rect 24636 17484 24642 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6914 17320 6920 17332
rect 5859 17292 6920 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7024 17292 7512 17320
rect 7024 17252 7052 17292
rect 6012 17224 7052 17252
rect 7484 17252 7512 17292
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 8444 17292 15853 17320
rect 8444 17280 8450 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16574 17320 16580 17332
rect 15979 17292 16580 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 23106 17320 23112 17332
rect 16908 17292 23112 17320
rect 16908 17280 16914 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23658 17320 23664 17332
rect 23216 17292 23664 17320
rect 9122 17252 9128 17264
rect 7484 17224 9128 17252
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4614 17184 4620 17196
rect 4111 17156 4620 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 4798 17144 4804 17196
rect 4856 17144 4862 17196
rect 6012 17193 6040 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 9493 17255 9551 17261
rect 9493 17221 9505 17255
rect 9539 17252 9551 17255
rect 9766 17252 9772 17264
rect 9539 17224 9772 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 11333 17255 11391 17261
rect 11333 17252 11345 17255
rect 10718 17224 11345 17252
rect 11333 17221 11345 17224
rect 11379 17252 11391 17255
rect 11606 17252 11612 17264
rect 11379 17224 11612 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 11974 17212 11980 17264
rect 12032 17212 12038 17264
rect 12710 17212 12716 17264
rect 12768 17212 12774 17264
rect 13446 17212 13452 17264
rect 13504 17252 13510 17264
rect 17862 17252 17868 17264
rect 13504 17224 16068 17252
rect 13504 17212 13510 17224
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 6733 17188 6791 17193
rect 6733 17187 6868 17188
rect 6733 17153 6745 17187
rect 6779 17184 6868 17187
rect 6914 17184 6920 17196
rect 6779 17160 6920 17184
rect 6779 17153 6791 17160
rect 6840 17156 6920 17160
rect 6733 17147 6791 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17188 7435 17193
rect 7377 17187 7512 17188
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17184 7512 17187
rect 7558 17184 7564 17196
rect 7423 17160 7564 17184
rect 7423 17153 7435 17160
rect 7484 17156 7564 17160
rect 7377 17147 7435 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 8021 17188 8079 17193
rect 7944 17187 8079 17188
rect 7944 17184 8033 17187
rect 7668 17160 8033 17184
rect 7668 17156 7972 17160
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4706 17116 4712 17128
rect 4571 17088 4712 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 7668 17116 7696 17156
rect 8021 17153 8033 17160
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8754 17184 8760 17196
rect 8352 17156 8760 17184
rect 8352 17144 8358 17156
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 9088 17156 9229 17184
rect 9088 17144 9094 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 11698 17184 11704 17196
rect 9217 17147 9275 17153
rect 11072 17156 11704 17184
rect 6604 17088 7696 17116
rect 6604 17076 6610 17088
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 9858 17116 9864 17128
rect 7984 17088 9864 17116
rect 7984 17076 7990 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10100 17088 10977 17116
rect 10100 17076 10106 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 3881 17051 3939 17057
rect 3881 17017 3893 17051
rect 3927 17048 3939 17051
rect 7466 17048 7472 17060
rect 3927 17020 6684 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 6546 16940 6552 16992
rect 6604 16940 6610 16992
rect 6656 16980 6684 17020
rect 6840 17020 7472 17048
rect 6840 16980 6868 17020
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 7616 17020 7849 17048
rect 7616 17008 7622 17020
rect 7837 17017 7849 17020
rect 7883 17017 7895 17051
rect 7837 17011 7895 17017
rect 8570 17008 8576 17060
rect 8628 17008 8634 17060
rect 6656 16952 6868 16980
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 8846 16980 8852 16992
rect 7239 16952 8852 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 11072 16980 11100 17156
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 14366 17144 14372 17196
rect 14424 17144 14430 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 12676 17088 13461 17116
rect 12676 17076 12682 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 16040 17125 16068 17224
rect 16132 17224 17868 17252
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 16025 17119 16083 17125
rect 13909 17079 13967 17085
rect 14292 17088 15240 17116
rect 9088 16952 11100 16980
rect 9088 16940 9094 16952
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 14292 16980 14320 17088
rect 14829 17051 14887 17057
rect 14829 17017 14841 17051
rect 14875 17048 14887 17051
rect 15102 17048 15108 17060
rect 14875 17020 15108 17048
rect 14875 17017 14887 17020
rect 14829 17011 14887 17017
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 15212 17048 15240 17088
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16132 17048 16160 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 18874 17252 18880 17264
rect 18248 17224 18880 17252
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 18248 17184 18276 17224
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 21453 17255 21511 17261
rect 21453 17221 21465 17255
rect 21499 17252 21511 17255
rect 21542 17252 21548 17264
rect 21499 17224 21548 17252
rect 21499 17221 21511 17224
rect 21453 17215 21511 17221
rect 21542 17212 21548 17224
rect 21600 17212 21606 17264
rect 22094 17212 22100 17264
rect 22152 17252 22158 17264
rect 23216 17252 23244 17292
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 24302 17280 24308 17332
rect 24360 17280 24366 17332
rect 24118 17252 24124 17264
rect 22152 17224 23244 17252
rect 24058 17224 24124 17252
rect 22152 17212 22158 17224
rect 24118 17212 24124 17224
rect 24176 17212 24182 17264
rect 25130 17252 25136 17264
rect 24780 17224 25136 17252
rect 17359 17156 18276 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 20809 17187 20867 17193
rect 19734 17156 20484 17184
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17736 17088 17877 17116
rect 17736 17076 17742 17088
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 19150 17116 19156 17128
rect 18647 17088 19156 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 20070 17116 20076 17128
rect 19392 17088 20076 17116
rect 19392 17076 19398 17088
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20456 17125 20484 17156
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 22278 17184 22284 17196
rect 20855 17156 22284 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 24780 17184 24808 17224
rect 25130 17212 25136 17224
rect 25188 17212 25194 17264
rect 24044 17156 24808 17184
rect 24857 17187 24915 17193
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 21266 17116 21272 17128
rect 20487 17088 21272 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 21266 17076 21272 17088
rect 21324 17116 21330 17128
rect 21818 17116 21824 17128
rect 21324 17088 21824 17116
rect 21324 17076 21330 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22833 17119 22891 17125
rect 22833 17085 22845 17119
rect 22879 17116 22891 17119
rect 24044 17116 24072 17156
rect 24857 17153 24869 17187
rect 24903 17153 24915 17187
rect 24857 17147 24915 17153
rect 22879 17088 24072 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 15212 17020 16160 17048
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 16540 17020 18000 17048
rect 16540 17008 16546 17020
rect 12032 16952 14320 16980
rect 12032 16940 12038 16952
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 15068 16952 15485 16980
rect 15068 16940 15074 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16632 16952 16865 16980
rect 16632 16940 16638 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 17972 16980 18000 17020
rect 19628 17020 22692 17048
rect 19628 16980 19656 17020
rect 17972 16952 19656 16980
rect 16853 16943 16911 16949
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 21266 16980 21272 16992
rect 20680 16952 21272 16980
rect 20680 16940 20686 16952
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21876 16952 22017 16980
rect 21876 16940 21882 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 22005 16943 22063 16949
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22370 16980 22376 16992
rect 22327 16952 22376 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 22664 16980 22692 17020
rect 24872 16980 24900 17147
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 25498 17048 25504 17060
rect 25087 17020 25504 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 25498 17008 25504 17020
rect 25556 17008 25562 17060
rect 25317 16983 25375 16989
rect 25317 16980 25329 16983
rect 22664 16952 25329 16980
rect 25317 16949 25329 16952
rect 25363 16949 25375 16983
rect 25317 16943 25375 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 4249 16779 4307 16785
rect 4249 16745 4261 16779
rect 4295 16776 4307 16779
rect 4614 16776 4620 16788
rect 4295 16748 4620 16776
rect 4295 16745 4307 16748
rect 4249 16739 4307 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 7926 16776 7932 16788
rect 4764 16748 7932 16776
rect 4764 16736 4770 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8386 16736 8392 16788
rect 8444 16736 8450 16788
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9398 16776 9404 16788
rect 9079 16748 9404 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 15010 16776 15016 16788
rect 11256 16748 15016 16776
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 11054 16708 11060 16720
rect 6972 16680 11060 16708
rect 6972 16668 6978 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 7282 16600 7288 16652
rect 7340 16600 7346 16652
rect 7469 16643 7527 16649
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 8662 16640 8668 16652
rect 7515 16612 8668 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 7944 16581 7972 16612
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 10042 16640 10048 16652
rect 9263 16612 10048 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 11256 16649 11284 16748
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 19692 16779 19750 16785
rect 19692 16745 19704 16779
rect 19738 16776 19750 16779
rect 21726 16776 21732 16788
rect 19738 16748 21732 16776
rect 19738 16745 19750 16748
rect 19692 16739 19750 16745
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 25225 16779 25283 16785
rect 25225 16776 25237 16779
rect 22336 16748 25237 16776
rect 22336 16736 22342 16748
rect 25225 16745 25237 16748
rect 25271 16745 25283 16779
rect 25225 16739 25283 16745
rect 19334 16668 19340 16720
rect 19392 16668 19398 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21542 16708 21548 16720
rect 20772 16680 21548 16708
rect 20772 16668 20778 16680
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11425 16643 11483 16649
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 12250 16640 12256 16652
rect 11471 16612 12256 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14918 16640 14924 16652
rect 14323 16612 14924 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 19352 16640 19380 16668
rect 17451 16612 19380 16640
rect 19429 16643 19487 16649
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 22278 16640 22284 16652
rect 19475 16612 22284 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 22646 16640 22652 16652
rect 22603 16612 22652 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 8754 16572 8760 16584
rect 8619 16544 8760 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10962 16572 10968 16584
rect 9723 16544 10968 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11146 16532 11152 16584
rect 11204 16532 11210 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 21266 16532 21272 16584
rect 21324 16572 21330 16584
rect 21637 16575 21695 16581
rect 21637 16572 21649 16575
rect 21324 16544 21649 16572
rect 21324 16532 21330 16544
rect 21637 16541 21649 16544
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16572 24639 16575
rect 25222 16572 25228 16584
rect 24627 16544 25228 16572
rect 24627 16541 24639 16544
rect 24581 16535 24639 16541
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 5353 16507 5411 16513
rect 5353 16473 5365 16507
rect 5399 16504 5411 16507
rect 11790 16504 11796 16516
rect 5399 16476 11796 16504
rect 5399 16473 5411 16476
rect 5353 16467 5411 16473
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 12253 16507 12311 16513
rect 12253 16473 12265 16507
rect 12299 16504 12311 16507
rect 12526 16504 12532 16516
rect 12299 16476 12532 16504
rect 12299 16473 12311 16476
rect 12253 16467 12311 16473
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 14384 16476 14565 16504
rect 14384 16448 14412 16476
rect 14553 16473 14565 16476
rect 14599 16504 14611 16507
rect 14599 16476 14964 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 14936 16448 14964 16476
rect 15010 16464 15016 16516
rect 15068 16464 15074 16516
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 21818 16504 21824 16516
rect 16356 16476 17894 16504
rect 20930 16476 21824 16504
rect 16356 16464 16362 16476
rect 21468 16448 21496 16476
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 24118 16504 24124 16516
rect 23782 16476 24124 16504
rect 24118 16464 24124 16476
rect 24176 16464 24182 16516
rect 4706 16396 4712 16448
rect 4764 16396 4770 16448
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 8846 16436 8852 16448
rect 7791 16408 8852 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 9490 16396 9496 16448
rect 9548 16396 9554 16448
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 10778 16396 10784 16448
rect 10836 16396 10842 16448
rect 12342 16396 12348 16448
rect 12400 16436 12406 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12400 16408 13737 16436
rect 12400 16396 12406 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 14366 16396 14372 16448
rect 14424 16396 14430 16448
rect 14918 16396 14924 16448
rect 14976 16396 14982 16448
rect 16485 16439 16543 16445
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 18322 16436 18328 16448
rect 16531 16408 18328 16436
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 19150 16396 19156 16448
rect 19208 16436 19214 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 19208 16408 21189 16436
rect 19208 16396 19214 16408
rect 21177 16405 21189 16408
rect 21223 16436 21235 16439
rect 21266 16436 21272 16448
rect 21223 16408 21272 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21450 16396 21456 16448
rect 21508 16396 21514 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23992 16408 24041 16436
rect 23992 16396 23998 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 8021 16235 8079 16241
rect 8021 16201 8033 16235
rect 8067 16232 8079 16235
rect 8294 16232 8300 16244
rect 8067 16204 8300 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 9674 16232 9680 16244
rect 8404 16204 9680 16232
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 8404 16164 8432 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 9766 16192 9772 16244
rect 9824 16192 9830 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10192 16204 10793 16232
rect 10192 16192 10198 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 10980 16204 13400 16232
rect 4764 16136 8432 16164
rect 4764 16124 4770 16136
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 10980 16164 11008 16204
rect 9548 16136 11008 16164
rect 9548 16124 9554 16136
rect 12618 16124 12624 16176
rect 12676 16124 12682 16176
rect 13372 16164 13400 16204
rect 13446 16192 13452 16244
rect 13504 16192 13510 16244
rect 14550 16232 14556 16244
rect 13556 16204 14556 16232
rect 13556 16164 13584 16204
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 15010 16192 15016 16244
rect 15068 16232 15074 16244
rect 16298 16232 16304 16244
rect 15068 16204 16304 16232
rect 15068 16192 15074 16204
rect 16298 16192 16304 16204
rect 16356 16232 16362 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 16356 16204 16681 16232
rect 16356 16192 16362 16204
rect 16669 16201 16681 16204
rect 16715 16201 16727 16235
rect 16669 16195 16727 16201
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 18506 16232 18512 16244
rect 18463 16204 18512 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 19337 16235 19395 16241
rect 19337 16201 19349 16235
rect 19383 16201 19395 16235
rect 19337 16195 19395 16201
rect 13372 16136 13584 16164
rect 14369 16167 14427 16173
rect 14369 16133 14381 16167
rect 14415 16164 14427 16167
rect 19352 16164 19380 16195
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20533 16235 20591 16241
rect 19760 16204 19840 16232
rect 19760 16192 19766 16204
rect 14415 16136 19380 16164
rect 14415 16133 14427 16136
rect 14369 16127 14427 16133
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8662 16096 8668 16108
rect 8251 16068 8668 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16096 9367 16099
rect 9398 16096 9404 16108
rect 9355 16068 9404 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 10042 16096 10048 16108
rect 9999 16068 10048 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 11514 16096 11520 16108
rect 10152 16068 11520 16096
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 10152 16028 10180 16068
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13964 16068 14289 16096
rect 13964 16056 13970 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15562 16096 15568 16108
rect 15243 16068 15568 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15804 16068 15853 16096
rect 15804 16056 15810 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 18966 16096 18972 16108
rect 17175 16068 18972 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 19702 16056 19708 16108
rect 19760 16056 19766 16108
rect 8444 16000 10180 16028
rect 10873 16031 10931 16037
rect 8444 15988 8450 16000
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 6086 15920 6092 15972
rect 6144 15960 6150 15972
rect 6144 15932 9536 15960
rect 6144 15920 6150 15932
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 9122 15852 9128 15904
rect 9180 15852 9186 15904
rect 9508 15892 9536 15932
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 9640 15932 10425 15960
rect 9640 15920 9646 15932
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 10778 15892 10784 15904
rect 9508 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 10888 15892 10916 15991
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12342 16028 12348 16040
rect 12023 16000 12348 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13354 16028 13360 16040
rect 12492 16000 13360 16028
rect 12492 15988 12498 16000
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15580 16028 15608 16056
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15580 16000 15945 16028
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 16022 15988 16028 16040
rect 16080 15988 16086 16040
rect 19812 16037 19840 16204
rect 20533 16201 20545 16235
rect 20579 16201 20591 16235
rect 20533 16195 20591 16201
rect 20901 16235 20959 16241
rect 20901 16201 20913 16235
rect 20947 16232 20959 16235
rect 21082 16232 21088 16244
rect 20947 16204 21088 16232
rect 20947 16201 20959 16204
rect 20901 16195 20959 16201
rect 20548 16164 20576 16195
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 21910 16192 21916 16244
rect 21968 16232 21974 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 21968 16204 22477 16232
rect 21968 16192 21974 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 23842 16192 23848 16244
rect 23900 16192 23906 16244
rect 25222 16192 25228 16244
rect 25280 16192 25286 16244
rect 25774 16164 25780 16176
rect 20548 16136 25780 16164
rect 25774 16124 25780 16136
rect 25832 16124 25838 16176
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 20993 16099 21051 16105
rect 20993 16096 21005 16099
rect 20956 16068 21005 16096
rect 20956 16056 20962 16068
rect 20993 16065 21005 16068
rect 21039 16096 21051 16099
rect 21039 16068 21772 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 13372 15932 15485 15960
rect 13372 15892 13400 15932
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 17586 15960 17592 15972
rect 15473 15923 15531 15929
rect 15580 15932 17592 15960
rect 10888 15864 13400 15892
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13909 15895 13967 15901
rect 13909 15892 13921 15895
rect 13596 15864 13921 15892
rect 13596 15852 13602 15864
rect 13909 15861 13921 15864
rect 13955 15861 13967 15895
rect 13909 15855 13967 15861
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 15580 15892 15608 15932
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 19812 15960 19840 15991
rect 19886 15988 19892 16040
rect 19944 15988 19950 16040
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 19812 15932 20944 15960
rect 15068 15864 15608 15892
rect 15068 15852 15074 15864
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 20806 15892 20812 15904
rect 17460 15864 20812 15892
rect 17460 15852 17466 15864
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 20916 15892 20944 15932
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 21192 15960 21220 15991
rect 21140 15932 21220 15960
rect 21744 15960 21772 16068
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 23750 16056 23756 16108
rect 23808 16056 23814 16108
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 24578 16096 24584 16108
rect 24084 16068 24584 16096
rect 24084 16056 24090 16068
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22244 16000 22569 16028
rect 22244 15988 22250 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 23934 15988 23940 16040
rect 23992 15988 23998 16040
rect 23017 15963 23075 15969
rect 23017 15960 23029 15963
rect 21744 15932 23029 15960
rect 21140 15920 21146 15932
rect 23017 15929 23029 15932
rect 23063 15929 23075 15963
rect 23017 15923 23075 15929
rect 21545 15895 21603 15901
rect 21545 15892 21557 15895
rect 20916 15864 21557 15892
rect 21545 15861 21557 15864
rect 21591 15861 21603 15895
rect 21545 15855 21603 15861
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22186 15892 22192 15904
rect 22051 15864 22192 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22646 15852 22652 15904
rect 22704 15892 22710 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 22704 15864 23397 15892
rect 22704 15852 22710 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 9950 15688 9956 15700
rect 9907 15660 9956 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 12158 15688 12164 15700
rect 10612 15660 12164 15688
rect 9217 15623 9275 15629
rect 9217 15589 9229 15623
rect 9263 15620 9275 15623
rect 10612 15620 10640 15660
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 12526 15688 12532 15700
rect 12268 15660 12532 15688
rect 9263 15592 10640 15620
rect 9263 15589 9275 15592
rect 9217 15583 9275 15589
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 12268 15620 12296 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 14090 15688 14096 15700
rect 13863 15660 14096 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 15252 15660 16037 15688
rect 15252 15648 15258 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 16025 15651 16083 15657
rect 16666 15648 16672 15700
rect 16724 15648 16730 15700
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18012 15660 18705 15688
rect 18012 15648 18018 15660
rect 18693 15657 18705 15660
rect 18739 15688 18751 15691
rect 19794 15688 19800 15700
rect 18739 15660 19800 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19794 15648 19800 15660
rect 19852 15648 19858 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22738 15688 22744 15700
rect 22244 15660 22744 15688
rect 22244 15648 22250 15660
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 22833 15691 22891 15697
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 22922 15688 22928 15700
rect 22879 15660 22928 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 22922 15648 22928 15660
rect 22980 15648 22986 15700
rect 24118 15648 24124 15700
rect 24176 15648 24182 15700
rect 24578 15648 24584 15700
rect 24636 15688 24642 15700
rect 25317 15691 25375 15697
rect 25317 15688 25329 15691
rect 24636 15660 25329 15688
rect 24636 15648 24642 15660
rect 25317 15657 25329 15660
rect 25363 15657 25375 15691
rect 25317 15651 25375 15657
rect 11848 15592 12296 15620
rect 11848 15580 11854 15592
rect 12342 15580 12348 15632
rect 12400 15620 12406 15632
rect 13538 15620 13544 15632
rect 12400 15592 13544 15620
rect 12400 15580 12406 15592
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 21634 15620 21640 15632
rect 18380 15592 21640 15620
rect 18380 15580 18386 15592
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 24026 15620 24032 15632
rect 22066 15592 24032 15620
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 10410 15552 10416 15564
rect 8996 15524 10416 15552
rect 8996 15512 9002 15524
rect 10410 15512 10416 15524
rect 10468 15512 10474 15564
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 13262 15552 13268 15564
rect 10827 15524 13268 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14182 15552 14188 15564
rect 13403 15524 14188 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 16850 15552 16856 15564
rect 14332 15524 16856 15552
rect 14332 15512 14338 15524
rect 16850 15512 16856 15524
rect 16908 15552 16914 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16908 15524 16957 15552
rect 16908 15512 16914 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 18874 15552 18880 15564
rect 17267 15524 18880 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 18874 15512 18880 15524
rect 18932 15552 18938 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 18932 15524 20085 15552
rect 18932 15512 18938 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 21174 15512 21180 15564
rect 21232 15512 21238 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 22066 15552 22094 15592
rect 24026 15580 24032 15592
rect 24084 15580 24090 15632
rect 21560 15524 22094 15552
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10226 15484 10232 15496
rect 10091 15456 10232 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13814 15484 13820 15496
rect 13127 15456 13820 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 10520 15416 10548 15447
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 16298 15484 16304 15496
rect 15686 15456 16304 15484
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 18322 15444 18328 15496
rect 18380 15444 18386 15496
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 20898 15484 20904 15496
rect 18656 15456 20904 15484
rect 18656 15444 18662 15456
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21560 15484 21588 15524
rect 22830 15512 22836 15564
rect 22888 15552 22894 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 22888 15524 25145 15552
rect 22888 15512 22894 15524
rect 24688 15493 24716 15524
rect 25133 15521 25145 15524
rect 25179 15521 25191 15555
rect 25133 15515 25191 15521
rect 25590 15512 25596 15564
rect 25648 15552 25654 15564
rect 26234 15552 26240 15564
rect 25648 15524 26240 15552
rect 25648 15512 25654 15524
rect 26234 15512 26240 15524
rect 26292 15512 26298 15564
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 21131 15456 21588 15484
rect 21652 15456 23397 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 10686 15416 10692 15428
rect 10520 15388 10692 15416
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 12618 15416 12624 15428
rect 12006 15388 12624 15416
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 10962 15348 10968 15360
rect 7800 15320 10968 15348
rect 7800 15308 7806 15320
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 12084 15348 12112 15388
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13173 15419 13231 15425
rect 13173 15385 13185 15419
rect 13219 15416 13231 15419
rect 14553 15419 14611 15425
rect 13219 15388 14504 15416
rect 13219 15385 13231 15388
rect 13173 15379 13231 15385
rect 11204 15320 12112 15348
rect 11204 15308 11210 15320
rect 12250 15308 12256 15360
rect 12308 15308 12314 15360
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 12400 15320 12725 15348
rect 12400 15308 12406 15320
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 14476 15348 14504 15388
rect 14553 15385 14565 15419
rect 14599 15416 14611 15419
rect 14642 15416 14648 15428
rect 14599 15388 14648 15416
rect 14599 15385 14611 15388
rect 14553 15379 14611 15385
rect 14642 15376 14648 15388
rect 14700 15376 14706 15428
rect 16574 15416 16580 15428
rect 15856 15388 16580 15416
rect 15856 15348 15884 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 14476 15320 15884 15348
rect 12713 15311 12771 15317
rect 16298 15308 16304 15360
rect 16356 15308 16362 15360
rect 18340 15348 18368 15444
rect 19889 15419 19947 15425
rect 19889 15385 19901 15419
rect 19935 15416 19947 15419
rect 21652 15416 21680 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15453 24731 15487
rect 24673 15447 24731 15453
rect 19935 15388 21680 15416
rect 22005 15419 22063 15425
rect 19935 15385 19947 15388
rect 19889 15379 19947 15385
rect 22005 15385 22017 15419
rect 22051 15385 22063 15419
rect 22005 15379 22063 15385
rect 19061 15351 19119 15357
rect 19061 15348 19073 15351
rect 18340 15320 19073 15348
rect 19061 15317 19073 15320
rect 19107 15348 19119 15351
rect 19242 15348 19248 15360
rect 19107 15320 19248 15348
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 19978 15308 19984 15360
rect 20036 15308 20042 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 22020 15348 22048 15379
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 22741 15419 22799 15425
rect 22741 15416 22753 15419
rect 22428 15388 22753 15416
rect 22428 15376 22434 15388
rect 22741 15385 22753 15388
rect 22787 15416 22799 15419
rect 23845 15419 23903 15425
rect 23845 15416 23857 15419
rect 22787 15388 23857 15416
rect 22787 15385 22799 15388
rect 22741 15379 22799 15385
rect 23845 15385 23857 15388
rect 23891 15385 23903 15419
rect 23845 15379 23903 15385
rect 24857 15419 24915 15425
rect 24857 15385 24869 15419
rect 24903 15416 24915 15419
rect 24946 15416 24952 15428
rect 24903 15388 24952 15416
rect 24903 15385 24915 15388
rect 24857 15379 24915 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 20956 15320 22048 15348
rect 22097 15351 22155 15357
rect 20956 15308 20962 15320
rect 22097 15317 22109 15351
rect 22143 15348 22155 15351
rect 26602 15348 26608 15360
rect 22143 15320 26608 15348
rect 22143 15317 22155 15320
rect 22097 15311 22155 15317
rect 26602 15308 26608 15320
rect 26660 15308 26666 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 9398 15104 9404 15156
rect 9456 15104 9462 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 10226 15144 10232 15156
rect 9723 15116 10232 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 13814 15144 13820 15156
rect 11256 15116 13820 15144
rect 9861 15079 9919 15085
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 11256 15076 11284 15116
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 13906 15104 13912 15156
rect 13964 15104 13970 15156
rect 16117 15147 16175 15153
rect 16117 15113 16129 15147
rect 16163 15144 16175 15147
rect 16163 15116 18920 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 9907 15048 11284 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11256 15008 11284 15048
rect 12618 15036 12624 15088
rect 12676 15036 12682 15088
rect 14642 15036 14648 15088
rect 14700 15076 14706 15088
rect 16758 15076 16764 15088
rect 14700 15048 16764 15076
rect 14700 15036 14706 15048
rect 16758 15036 16764 15048
rect 16816 15036 16822 15088
rect 17402 15076 17408 15088
rect 16868 15048 17408 15076
rect 11195 14980 11284 15008
rect 14553 15011 14611 15017
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 15010 15008 15016 15020
rect 14599 14980 15016 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 16022 15008 16028 15020
rect 15120 14980 16028 15008
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10091 14912 10640 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10318 14832 10324 14884
rect 10376 14832 10382 14884
rect 10612 14872 10640 14912
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12526 14940 12532 14952
rect 12023 14912 12532 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12526 14900 12532 14912
rect 12584 14940 12590 14952
rect 15120 14940 15148 14980
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16868 15008 16896 15048
rect 17402 15036 17408 15048
rect 17460 15036 17466 15088
rect 18892 15076 18920 15116
rect 18966 15104 18972 15156
rect 19024 15104 19030 15156
rect 21266 15144 21272 15156
rect 19996 15116 21272 15144
rect 19996 15076 20024 15116
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 21358 15104 21364 15156
rect 21416 15104 21422 15156
rect 23934 15144 23940 15156
rect 23124 15116 23940 15144
rect 21450 15076 21456 15088
rect 18892 15048 20024 15076
rect 20838 15048 21456 15076
rect 21450 15036 21456 15048
rect 21508 15036 21514 15088
rect 21542 15036 21548 15088
rect 21600 15076 21606 15088
rect 22097 15079 22155 15085
rect 22097 15076 22109 15079
rect 21600 15048 22109 15076
rect 21600 15036 21606 15048
rect 22097 15045 22109 15048
rect 22143 15045 22155 15079
rect 22097 15039 22155 15045
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 23014 15076 23020 15088
rect 22244 15048 23020 15076
rect 22244 15036 22250 15048
rect 23014 15036 23020 15048
rect 23072 15036 23078 15088
rect 23124 15085 23152 15116
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24394 15104 24400 15156
rect 24452 15144 24458 15156
rect 24581 15147 24639 15153
rect 24581 15144 24593 15147
rect 24452 15116 24593 15144
rect 24452 15104 24458 15116
rect 24581 15113 24593 15116
rect 24627 15113 24639 15147
rect 24581 15107 24639 15113
rect 23109 15079 23167 15085
rect 23109 15045 23121 15079
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 16132 14980 16896 15008
rect 12584 14912 15148 14940
rect 12584 14900 12590 14912
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 15436 14912 15485 14940
rect 15436 14900 15442 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 11146 14872 11152 14884
rect 10612 14844 11152 14872
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 16132 14872 16160 14980
rect 18230 14968 18236 15020
rect 18288 14968 18294 15020
rect 21008 14980 22094 15008
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17129 14943 17187 14949
rect 16899 14912 16988 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 13596 14844 16160 14872
rect 13596 14832 13602 14844
rect 10962 14764 10968 14816
rect 11020 14764 11026 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 12066 14804 12072 14816
rect 11112 14776 12072 14804
rect 11112 14764 11118 14776
rect 12066 14764 12072 14776
rect 12124 14804 12130 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 12124 14776 13461 14804
rect 12124 14764 12130 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 13449 14767 13507 14773
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14804 14887 14807
rect 16390 14804 16396 14816
rect 14875 14776 16396 14804
rect 14875 14773 14887 14776
rect 14829 14767 14887 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16960 14804 16988 14912
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17862 14940 17868 14952
rect 17175 14912 17868 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 19334 14940 19340 14952
rect 18156 14912 19340 14940
rect 17126 14804 17132 14816
rect 16540 14776 17132 14804
rect 16540 14764 16546 14776
rect 17126 14764 17132 14776
rect 17184 14804 17190 14816
rect 18156 14804 18184 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 19659 14912 20760 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20732 14884 20760 14912
rect 20714 14832 20720 14884
rect 20772 14832 20778 14884
rect 17184 14776 18184 14804
rect 17184 14764 17190 14776
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19794 14764 19800 14816
rect 19852 14804 19858 14816
rect 21008 14804 21036 14980
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21726 14940 21732 14952
rect 21131 14912 21732 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 21726 14900 21732 14912
rect 21784 14900 21790 14952
rect 22066 14940 22094 14980
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22336 14980 22845 15008
rect 22336 14968 22342 14980
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 24210 14968 24216 15020
rect 24268 14968 24274 15020
rect 25130 14968 25136 15020
rect 25188 14968 25194 15020
rect 23198 14940 23204 14952
rect 22066 14912 23204 14940
rect 23198 14900 23204 14912
rect 23256 14900 23262 14952
rect 21266 14832 21272 14884
rect 21324 14872 21330 14884
rect 22094 14872 22100 14884
rect 21324 14844 22100 14872
rect 21324 14832 21330 14844
rect 22094 14832 22100 14844
rect 22152 14832 22158 14884
rect 25314 14832 25320 14884
rect 25372 14832 25378 14884
rect 19852 14776 21036 14804
rect 19852 14764 19858 14776
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 21508 14776 21557 14804
rect 21508 14764 21514 14776
rect 21545 14773 21557 14776
rect 21591 14773 21603 14807
rect 21545 14767 21603 14773
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 23290 14804 23296 14816
rect 22235 14776 23296 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10502 14600 10508 14612
rect 10459 14572 10508 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12526 14600 12532 14612
rect 12483 14572 12532 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 24762 14600 24768 14612
rect 13872 14572 24768 14600
rect 13872 14560 13878 14572
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 25188 14572 25329 14600
rect 25188 14560 25194 14572
rect 25317 14569 25329 14572
rect 25363 14569 25375 14603
rect 25317 14563 25375 14569
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 16206 14532 16212 14544
rect 15988 14504 16212 14532
rect 15988 14492 15994 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18690 14532 18696 14544
rect 18279 14504 18696 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14532 19487 14535
rect 20070 14532 20076 14544
rect 19475 14504 20076 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 20070 14492 20076 14504
rect 20128 14492 20134 14544
rect 20530 14492 20536 14544
rect 20588 14532 20594 14544
rect 21450 14532 21456 14544
rect 20588 14504 21456 14532
rect 20588 14492 20594 14504
rect 21450 14492 21456 14504
rect 21508 14492 21514 14544
rect 21542 14492 21548 14544
rect 21600 14532 21606 14544
rect 23293 14535 23351 14541
rect 23293 14532 23305 14535
rect 21600 14504 23305 14532
rect 21600 14492 21606 14504
rect 23293 14501 23305 14504
rect 23339 14501 23351 14535
rect 23842 14532 23848 14544
rect 23293 14495 23351 14501
rect 23400 14504 23848 14532
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 12250 14464 12256 14476
rect 11011 14436 12256 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 18598 14464 18604 14476
rect 16807 14436 18604 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18598 14424 18604 14436
rect 18656 14464 18662 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 18656 14436 19993 14464
rect 18656 14424 18662 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 21910 14424 21916 14476
rect 21968 14464 21974 14476
rect 22278 14464 22284 14476
rect 21968 14436 22284 14464
rect 21968 14424 21974 14436
rect 22278 14424 22284 14436
rect 22336 14464 22342 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 22336 14436 22385 14464
rect 22336 14424 22342 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 22925 14467 22983 14473
rect 22925 14433 22937 14467
rect 22971 14464 22983 14467
rect 23400 14464 23428 14504
rect 23842 14492 23848 14504
rect 23900 14532 23906 14544
rect 24210 14532 24216 14544
rect 23900 14504 24216 14532
rect 23900 14492 23906 14504
rect 24210 14492 24216 14504
rect 24268 14532 24274 14544
rect 25225 14535 25283 14541
rect 25225 14532 25237 14535
rect 24268 14504 25237 14532
rect 24268 14492 24274 14504
rect 25225 14501 25237 14504
rect 25271 14501 25283 14535
rect 25225 14495 25283 14501
rect 22971 14436 23428 14464
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23532 14436 23765 14464
rect 23532 14424 23538 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24578 14464 24584 14476
rect 23983 14436 24584 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 14090 14396 14096 14408
rect 13127 14368 14096 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 15930 14396 15936 14408
rect 15686 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14396 15994 14408
rect 16298 14396 16304 14408
rect 15988 14368 16304 14396
rect 15988 14356 15994 14368
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16482 14356 16488 14408
rect 16540 14356 16546 14408
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19889 14399 19947 14405
rect 19889 14396 19901 14399
rect 19484 14368 19901 14396
rect 19484 14356 19490 14368
rect 19889 14365 19901 14368
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14396 20867 14399
rect 21358 14396 21364 14408
rect 20855 14368 21364 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 24118 14356 24124 14408
rect 24176 14396 24182 14408
rect 24673 14399 24731 14405
rect 24673 14396 24685 14399
rect 24176 14368 24685 14396
rect 24176 14356 24182 14368
rect 24673 14365 24685 14368
rect 24719 14365 24731 14399
rect 24673 14359 24731 14365
rect 12618 14328 12624 14340
rect 12190 14300 12624 14328
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 18230 14328 18236 14340
rect 12912 14300 14964 14328
rect 12912 14269 12940 14300
rect 12897 14263 12955 14269
rect 12897 14229 12909 14263
rect 12943 14229 12955 14263
rect 12897 14223 12955 14229
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14090 14260 14096 14272
rect 13872 14232 14096 14260
rect 13872 14220 13878 14232
rect 14090 14220 14096 14232
rect 14148 14260 14154 14272
rect 14366 14260 14372 14272
rect 14148 14232 14372 14260
rect 14148 14220 14154 14232
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 14936 14260 14964 14300
rect 15856 14300 17172 14328
rect 17986 14300 18236 14328
rect 15856 14260 15884 14300
rect 17144 14272 17172 14300
rect 18230 14288 18236 14300
rect 18288 14288 18294 14340
rect 18693 14331 18751 14337
rect 18693 14297 18705 14331
rect 18739 14328 18751 14331
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 18739 14300 19809 14328
rect 18739 14297 18751 14300
rect 18693 14291 18751 14297
rect 19797 14297 19809 14300
rect 19843 14297 19855 14331
rect 23382 14328 23388 14340
rect 19797 14291 19855 14297
rect 19996 14300 23388 14328
rect 14936 14232 15884 14260
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16758 14260 16764 14272
rect 16071 14232 16764 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 17126 14220 17132 14272
rect 17184 14220 17190 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19996 14260 20024 14300
rect 23382 14288 23388 14300
rect 23440 14288 23446 14340
rect 24857 14331 24915 14337
rect 24857 14297 24869 14331
rect 24903 14328 24915 14331
rect 25406 14328 25412 14340
rect 24903 14300 25412 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 25406 14288 25412 14300
rect 25464 14288 25470 14340
rect 18656 14232 20024 14260
rect 18656 14220 18662 14232
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 22002 14260 22008 14272
rect 20956 14232 22008 14260
rect 20956 14220 20962 14232
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 23658 14220 23664 14272
rect 23716 14220 23722 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11330 14056 11336 14068
rect 11195 14028 11336 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11793 14059 11851 14065
rect 11793 14025 11805 14059
rect 11839 14056 11851 14059
rect 11882 14056 11888 14068
rect 11839 14028 11888 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12802 14056 12808 14068
rect 12483 14028 12808 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 13998 14056 14004 14068
rect 13127 14028 14004 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14700 14028 15485 14056
rect 14700 14016 14706 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 15896 14028 16129 14056
rect 15896 14016 15902 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17126 14056 17132 14068
rect 17083 14028 17132 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17604 14028 18644 14056
rect 11348 13920 11376 14016
rect 14274 13988 14280 14000
rect 13740 13960 14280 13988
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11348 13892 11989 13920
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13265 13923 13323 13929
rect 12667 13892 12701 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13630 13920 13636 13932
rect 13311 13892 13636 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 12636 13852 12664 13883
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13740 13929 13768 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 15930 13988 15936 14000
rect 15226 13960 15936 13988
rect 15930 13948 15936 13960
rect 15988 13948 15994 14000
rect 17604 13988 17632 14028
rect 16316 13960 17632 13988
rect 18233 13991 18291 13997
rect 16316 13929 16344 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18506 13988 18512 14000
rect 18279 13960 18512 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 18616 13988 18644 14028
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 20530 14056 20536 14068
rect 19300 14028 20536 14056
rect 19300 14016 19306 14028
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 20680 14028 21189 14056
rect 20680 14016 20686 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 22646 14056 22652 14068
rect 22060 14028 22652 14056
rect 22060 14016 22066 14028
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 19794 13988 19800 14000
rect 18616 13960 19800 13988
rect 19794 13948 19800 13960
rect 19852 13948 19858 14000
rect 20898 13988 20904 14000
rect 19904 13960 20904 13988
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 16448 13892 17356 13920
rect 16448 13880 16454 13892
rect 14458 13852 14464 13864
rect 11379 13824 14464 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 17328 13852 17356 13892
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 19904 13920 19932 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21085 13991 21143 13997
rect 21085 13957 21097 13991
rect 21131 13988 21143 13991
rect 21726 13988 21732 14000
rect 21131 13960 21732 13988
rect 21131 13957 21143 13960
rect 21085 13951 21143 13957
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 23382 13988 23388 14000
rect 22204 13960 23388 13988
rect 17512 13892 19932 13920
rect 17512 13852 17540 13892
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20772 13892 21312 13920
rect 20772 13880 20778 13892
rect 17328 13824 17540 13852
rect 17586 13812 17592 13864
rect 17644 13812 17650 13864
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 21284 13861 21312 13892
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22204 13920 22232 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 23842 13948 23848 14000
rect 23900 13948 23906 14000
rect 22152 13892 22232 13920
rect 22152 13880 22158 13892
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22336 13892 22845 13920
rect 22336 13880 22342 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 25866 13920 25872 13932
rect 25188 13892 25872 13920
rect 25188 13880 25194 13892
rect 25866 13880 25872 13892
rect 25924 13880 25930 13932
rect 21269 13855 21327 13861
rect 20036 13824 21220 13852
rect 20036 13812 20042 13824
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 18506 13784 18512 13796
rect 15620 13756 18512 13784
rect 15620 13744 15626 13756
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 19518 13744 19524 13796
rect 19576 13784 19582 13796
rect 21192 13784 21220 13824
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21450 13852 21456 13864
rect 21315 13824 21456 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21450 13812 21456 13824
rect 21508 13812 21514 13864
rect 23109 13855 23167 13861
rect 21560 13824 22324 13852
rect 21560 13784 21588 13824
rect 22296 13793 22324 13824
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 24394 13852 24400 13864
rect 23155 13824 24400 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24578 13812 24584 13864
rect 24636 13812 24642 13864
rect 25222 13812 25228 13864
rect 25280 13852 25286 13864
rect 25317 13855 25375 13861
rect 25317 13852 25329 13855
rect 25280 13824 25329 13852
rect 25280 13812 25286 13824
rect 25317 13821 25329 13824
rect 25363 13821 25375 13855
rect 25317 13815 25375 13821
rect 19576 13756 20852 13784
rect 21192 13756 21588 13784
rect 22281 13787 22339 13793
rect 19576 13744 19582 13756
rect 13998 13725 14004 13728
rect 13988 13719 14004 13725
rect 13988 13685 14000 13719
rect 13988 13679 14004 13685
rect 13998 13676 14004 13679
rect 14056 13676 14062 13728
rect 15841 13719 15899 13725
rect 15841 13685 15853 13719
rect 15887 13716 15899 13719
rect 15930 13716 15936 13728
rect 15887 13688 15936 13716
rect 15887 13685 15899 13688
rect 15841 13679 15899 13685
rect 15930 13676 15936 13688
rect 15988 13716 15994 13728
rect 16574 13716 16580 13728
rect 15988 13688 16580 13716
rect 15988 13676 15994 13688
rect 16574 13676 16580 13688
rect 16632 13716 16638 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16632 13688 16681 13716
rect 16632 13676 16638 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17310 13716 17316 13728
rect 16816 13688 17316 13716
rect 16816 13676 16822 13688
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 19426 13676 19432 13728
rect 19484 13716 19490 13728
rect 19705 13719 19763 13725
rect 19705 13716 19717 13719
rect 19484 13688 19717 13716
rect 19484 13676 19490 13688
rect 19705 13685 19717 13688
rect 19751 13685 19763 13719
rect 19705 13679 19763 13685
rect 20349 13719 20407 13725
rect 20349 13685 20361 13719
rect 20395 13716 20407 13719
rect 20530 13716 20536 13728
rect 20395 13688 20536 13716
rect 20395 13685 20407 13688
rect 20349 13679 20407 13685
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 20824 13716 20852 13756
rect 22281 13753 22293 13787
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 22738 13716 22744 13728
rect 20824 13688 22744 13716
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 14056 13484 16037 13512
rect 14056 13472 14062 13484
rect 16025 13481 16037 13484
rect 16071 13512 16083 13515
rect 18693 13515 18751 13521
rect 16071 13484 17816 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 13541 13447 13599 13453
rect 13541 13444 13553 13447
rect 13412 13416 13553 13444
rect 13412 13404 13418 13416
rect 13541 13413 13553 13416
rect 13587 13444 13599 13447
rect 17788 13444 17816 13484
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19702 13512 19708 13524
rect 18739 13484 19708 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 19794 13472 19800 13524
rect 19852 13472 19858 13524
rect 19968 13515 20026 13521
rect 19968 13481 19980 13515
rect 20014 13512 20026 13515
rect 20990 13512 20996 13524
rect 20014 13484 20996 13512
rect 20014 13481 20026 13484
rect 19968 13475 20026 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21450 13472 21456 13524
rect 21508 13472 21514 13524
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 23937 13515 23995 13521
rect 23937 13512 23949 13515
rect 23532 13484 23949 13512
rect 23532 13472 23538 13484
rect 23937 13481 23949 13484
rect 23983 13481 23995 13515
rect 23937 13475 23995 13481
rect 19337 13447 19395 13453
rect 13587 13416 14412 13444
rect 17788 13416 18828 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 12066 13336 12072 13388
rect 12124 13336 12130 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14384 13376 14412 13416
rect 14384 13348 15884 13376
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 11514 13240 11520 13252
rect 9631 13212 11520 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10686 13172 10692 13184
rect 10100 13144 10692 13172
rect 10100 13132 10106 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13172 10931 13175
rect 11808 13172 11836 13271
rect 13446 13240 13452 13252
rect 13294 13212 13452 13240
rect 13446 13200 13452 13212
rect 13504 13240 13510 13252
rect 13504 13212 13952 13240
rect 13504 13200 13510 13212
rect 13924 13181 13952 13212
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14550 13240 14556 13252
rect 14240 13212 14556 13240
rect 14240 13200 14246 13212
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 10919 13144 11836 13172
rect 13909 13175 13967 13181
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 15672 13172 15700 13294
rect 15856 13240 15884 13348
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18690 13376 18696 13388
rect 16807 13348 18696 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 18800 13376 18828 13416
rect 19337 13413 19349 13447
rect 19383 13444 19395 13447
rect 19812 13444 19840 13472
rect 19383 13416 19840 13444
rect 21008 13444 21036 13472
rect 21008 13416 22048 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 21910 13376 21916 13388
rect 18800 13348 19656 13376
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19518 13308 19524 13320
rect 18923 13280 19524 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 16758 13240 16764 13252
rect 15856 13212 16764 13240
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 19628 13240 19656 13348
rect 19720 13348 21916 13376
rect 19720 13320 19748 13348
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22020 13376 22048 13416
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23900 13416 24133 13444
rect 23900 13404 23906 13416
rect 24121 13413 24133 13416
rect 24167 13444 24179 13447
rect 24762 13444 24768 13456
rect 24167 13416 24768 13444
rect 24167 13413 24179 13416
rect 24121 13407 24179 13413
rect 24762 13404 24768 13416
rect 24820 13404 24826 13456
rect 23661 13379 23719 13385
rect 23661 13376 23673 13379
rect 22020 13348 23673 13376
rect 23661 13345 23673 13348
rect 23707 13345 23719 13379
rect 23661 13339 23719 13345
rect 19702 13268 19708 13320
rect 19760 13268 19766 13320
rect 23860 13308 23888 13404
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 25041 13379 25099 13385
rect 25041 13376 25053 13379
rect 24912 13348 25053 13376
rect 24912 13336 24918 13348
rect 25041 13345 25053 13348
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 23322 13280 23888 13308
rect 19886 13240 19892 13252
rect 18892 13212 19380 13240
rect 19628 13212 19892 13240
rect 18892 13184 18920 13212
rect 15930 13172 15936 13184
rect 13955 13144 15936 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17586 13172 17592 13184
rect 16356 13144 17592 13172
rect 16356 13132 16362 13144
rect 17586 13132 17592 13144
rect 17644 13172 17650 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 17644 13144 18245 13172
rect 17644 13132 17650 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 18233 13135 18291 13141
rect 18874 13132 18880 13184
rect 18932 13132 18938 13184
rect 19352 13172 19380 13212
rect 19886 13200 19892 13212
rect 19944 13200 19950 13252
rect 20990 13200 20996 13252
rect 21048 13200 21054 13252
rect 22186 13200 22192 13252
rect 22244 13200 22250 13252
rect 24949 13243 25007 13249
rect 23492 13212 24624 13240
rect 23492 13172 23520 13212
rect 24596 13181 24624 13212
rect 24949 13209 24961 13243
rect 24995 13240 25007 13243
rect 25590 13240 25596 13252
rect 24995 13212 25596 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 25590 13200 25596 13212
rect 25648 13200 25654 13252
rect 19352 13144 23520 13172
rect 24581 13175 24639 13181
rect 24581 13141 24593 13175
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11572 12940 12434 12968
rect 11572 12928 11578 12940
rect 12406 12900 12434 12940
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 13446 12968 13452 12980
rect 12676 12940 13452 12968
rect 12676 12928 12682 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14274 12968 14280 12980
rect 13872 12940 14280 12968
rect 13872 12928 13878 12940
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 17368 12940 18460 12968
rect 17368 12928 17374 12940
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12406 12872 13001 12900
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 15562 12900 15568 12912
rect 13035 12872 15568 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 18432 12900 18460 12940
rect 19058 12928 19064 12980
rect 19116 12968 19122 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 19116 12940 19533 12968
rect 19116 12928 19122 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 19610 12928 19616 12980
rect 19668 12968 19674 12980
rect 20717 12971 20775 12977
rect 20717 12968 20729 12971
rect 19668 12940 20729 12968
rect 19668 12928 19674 12940
rect 20717 12937 20729 12940
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 21358 12928 21364 12980
rect 21416 12928 21422 12980
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 23753 12971 23811 12977
rect 23753 12968 23765 12971
rect 22244 12940 23765 12968
rect 22244 12928 22250 12940
rect 23753 12937 23765 12940
rect 23799 12968 23811 12971
rect 25130 12968 25136 12980
rect 23799 12940 25136 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 22554 12900 22560 12912
rect 18432 12872 22560 12900
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 23842 12900 23848 12912
rect 23506 12872 23848 12900
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24213 12903 24271 12909
rect 24213 12900 24225 12903
rect 24084 12872 24225 12900
rect 24084 12860 24090 12872
rect 24213 12869 24225 12872
rect 24259 12869 24271 12903
rect 24213 12863 24271 12869
rect 24762 12860 24768 12912
rect 24820 12900 24826 12912
rect 25317 12903 25375 12909
rect 25317 12900 25329 12903
rect 24820 12872 25329 12900
rect 24820 12860 24826 12872
rect 25317 12869 25329 12872
rect 25363 12869 25375 12903
rect 25317 12863 25375 12869
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 18230 12792 18236 12844
rect 18288 12792 18294 12844
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 18472 12804 19441 12832
rect 18472 12792 18478 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12832 20683 12835
rect 21634 12832 21640 12844
rect 20671 12804 21640 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 24670 12792 24676 12844
rect 24728 12832 24734 12844
rect 25041 12835 25099 12841
rect 25041 12832 25053 12835
rect 24728 12804 25053 12832
rect 24728 12792 24734 12804
rect 25041 12801 25053 12804
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 15194 12724 15200 12776
rect 15252 12724 15258 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 16666 12764 16672 12776
rect 15519 12736 16672 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17494 12764 17500 12776
rect 17175 12736 17500 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17494 12724 17500 12736
rect 17552 12764 17558 12776
rect 18322 12764 18328 12776
rect 17552 12736 18328 12764
rect 17552 12724 17558 12736
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 19058 12764 19064 12776
rect 18840 12736 19064 12764
rect 18840 12724 18846 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19628 12696 19656 12727
rect 18656 12668 19656 12696
rect 18656 12656 18662 12668
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20824 12696 20852 12727
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 20496 12668 20852 12696
rect 20496 12656 20502 12668
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 15988 12600 16405 12628
rect 15988 12588 15994 12600
rect 16393 12597 16405 12600
rect 16439 12628 16451 12631
rect 16574 12628 16580 12640
rect 16439 12600 16580 12628
rect 16439 12597 16451 12600
rect 16393 12591 16451 12597
rect 16574 12588 16580 12600
rect 16632 12628 16638 12640
rect 17862 12628 17868 12640
rect 16632 12600 17868 12628
rect 16632 12588 16638 12600
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18506 12628 18512 12640
rect 18380 12600 18512 12628
rect 18380 12588 18386 12600
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19242 12628 19248 12640
rect 19107 12600 19248 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 20898 12628 20904 12640
rect 20588 12600 20904 12628
rect 20588 12588 20594 12600
rect 20898 12588 20904 12600
rect 20956 12628 20962 12640
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 20956 12600 21465 12628
rect 20956 12588 20962 12600
rect 21453 12597 21465 12600
rect 21499 12597 21511 12631
rect 21453 12591 21511 12597
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22646 12628 22652 12640
rect 22152 12600 22652 12628
rect 22152 12588 22158 12600
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 24026 12588 24032 12640
rect 24084 12628 24090 12640
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 24084 12600 24869 12628
rect 24084 12588 24090 12600
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 14090 12424 14096 12436
rect 13955 12396 14096 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15562 12424 15568 12436
rect 15519 12396 15568 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 15856 12396 17448 12424
rect 15856 12356 15884 12396
rect 14568 12328 15884 12356
rect 17420 12356 17448 12396
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18782 12424 18788 12436
rect 18288 12396 18788 12424
rect 18288 12384 18294 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 20824 12396 21312 12424
rect 17420 12328 19564 12356
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 14568 12297 14596 12328
rect 14553 12291 14611 12297
rect 4120 12260 14504 12288
rect 4120 12248 4126 12260
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13464 12192 14289 12220
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 13464 12093 13492 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 5776 12056 13461 12084
rect 5776 12044 5782 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 13725 12087 13783 12093
rect 13725 12053 13737 12087
rect 13771 12084 13783 12087
rect 14366 12084 14372 12096
rect 13771 12056 14372 12084
rect 13771 12053 13783 12056
rect 13725 12047 13783 12053
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14476 12084 14504 12260
rect 14553 12257 14565 12291
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16758 12288 16764 12300
rect 15795 12260 16764 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17460 12260 17969 12288
rect 17460 12248 17466 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 19536 12288 19564 12328
rect 20824 12288 20852 12396
rect 19536 12260 20852 12288
rect 18230 12220 18236 12232
rect 17158 12192 18236 12220
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16298 12152 16304 12164
rect 16071 12124 16304 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 18690 12161 18696 12164
rect 18657 12155 18696 12161
rect 18657 12152 18669 12155
rect 17328 12124 18669 12152
rect 17328 12084 17356 12124
rect 18657 12121 18669 12124
rect 18657 12115 18696 12121
rect 18690 12112 18696 12115
rect 18748 12112 18754 12164
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 19242 12152 19248 12164
rect 18923 12124 19248 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12121 19763 12155
rect 21284 12152 21312 12396
rect 22370 12384 22376 12436
rect 22428 12424 22434 12436
rect 24029 12427 24087 12433
rect 24029 12424 24041 12427
rect 22428 12396 24041 12424
rect 22428 12384 22434 12396
rect 24029 12393 24041 12396
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 24489 12427 24547 12433
rect 24489 12393 24501 12427
rect 24535 12424 24547 12427
rect 24670 12424 24676 12436
rect 24535 12396 24676 12424
rect 24535 12393 24547 12396
rect 24489 12387 24547 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21910 12288 21916 12300
rect 21416 12260 21916 12288
rect 21416 12248 21422 12260
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 24578 12288 24584 12300
rect 22603 12260 24584 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12220 21879 12223
rect 22094 12220 22100 12232
rect 21867 12192 22100 12220
rect 21867 12189 21879 12192
rect 21821 12183 21879 12189
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 24210 12220 24216 12232
rect 23690 12192 24216 12220
rect 24210 12180 24216 12192
rect 24268 12220 24274 12232
rect 24688 12220 24716 12384
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 24268 12192 24716 12220
rect 24268 12180 24274 12192
rect 21284 12124 22094 12152
rect 19705 12115 19763 12121
rect 14476 12056 17356 12084
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19720 12084 19748 12115
rect 20346 12084 20352 12096
rect 19392 12056 20352 12084
rect 19392 12044 19398 12056
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20496 12056 21189 12084
rect 20496 12044 20502 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 21177 12047 21235 12053
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 21637 12087 21695 12093
rect 21637 12084 21649 12087
rect 21324 12056 21649 12084
rect 21324 12044 21330 12056
rect 21637 12053 21649 12056
rect 21683 12053 21695 12087
rect 22066 12084 22094 12124
rect 23934 12084 23940 12096
rect 22066 12056 23940 12084
rect 21637 12047 21695 12053
rect 23934 12044 23940 12056
rect 23992 12044 23998 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13814 11880 13820 11892
rect 12820 11852 13820 11880
rect 12820 11753 12848 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 14884 11852 16129 11880
rect 14884 11840 14890 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 17310 11880 17316 11892
rect 16807 11852 17316 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13354 11812 13360 11824
rect 13127 11784 13360 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 14366 11812 14372 11824
rect 14306 11784 14372 11812
rect 14366 11772 14372 11784
rect 14424 11812 14430 11824
rect 14734 11812 14740 11824
rect 14424 11784 14740 11812
rect 14424 11772 14430 11784
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 16776 11812 16804 11843
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18877 11883 18935 11889
rect 18877 11849 18889 11883
rect 18923 11880 18935 11883
rect 19334 11880 19340 11892
rect 18923 11852 19340 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19610 11840 19616 11892
rect 19668 11880 19674 11892
rect 19668 11852 21036 11880
rect 19668 11840 19674 11852
rect 18782 11812 18788 11824
rect 16316 11784 16804 11812
rect 18630 11784 18788 11812
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15841 11747 15899 11753
rect 15335 11716 15700 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15672 11688 15700 11716
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 15930 11744 15936 11756
rect 15887 11716 15936 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16316 11753 16344 11784
rect 18782 11772 18788 11784
rect 18840 11772 18846 11824
rect 19702 11812 19708 11824
rect 19444 11784 19708 11812
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 19444 11753 19472 11784
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16632 11716 17141 11744
rect 16632 11704 16638 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 20806 11704 20812 11756
rect 20864 11704 20870 11756
rect 15654 11636 15660 11688
rect 15712 11636 15718 11688
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 18598 11676 18604 11688
rect 17451 11648 18604 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 20438 11676 20444 11688
rect 19751 11648 20444 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 21008 11676 21036 11852
rect 21174 11840 21180 11892
rect 21232 11840 21238 11892
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 22094 11880 22100 11892
rect 21784 11852 22100 11880
rect 21784 11840 21790 11852
rect 22094 11840 22100 11852
rect 22152 11880 22158 11892
rect 23382 11880 23388 11892
rect 22152 11852 23388 11880
rect 22152 11840 22158 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22112 11676 22140 11707
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23624 11716 23949 11744
rect 23624 11704 23630 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 21008 11648 22140 11676
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 23842 11676 23848 11688
rect 22520 11648 23848 11676
rect 22520 11636 22526 11648
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 26326 11676 26332 11688
rect 25188 11648 26332 11676
rect 25188 11636 25194 11648
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 21266 11608 21272 11620
rect 21100 11580 21272 11608
rect 15102 11500 15108 11552
rect 15160 11500 15166 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 21100 11540 21128 11580
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 15620 11512 21128 11540
rect 15620 11500 15626 11512
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16022 11336 16028 11348
rect 15519 11308 16028 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17092 11308 17417 11336
rect 17092 11296 17098 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 20993 11339 21051 11345
rect 18656 11308 20576 11336
rect 18656 11296 18662 11308
rect 14734 11228 14740 11280
rect 14792 11268 14798 11280
rect 15930 11268 15936 11280
rect 14792 11240 15936 11268
rect 14792 11228 14798 11240
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 18690 11228 18696 11280
rect 18748 11268 18754 11280
rect 20441 11271 20499 11277
rect 20441 11268 20453 11271
rect 18748 11240 20453 11268
rect 18748 11228 18754 11240
rect 20441 11237 20453 11240
rect 20487 11237 20499 11271
rect 20548 11268 20576 11308
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 24486 11336 24492 11348
rect 21039 11308 24492 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 24486 11296 24492 11308
rect 24544 11296 24550 11348
rect 25317 11339 25375 11345
rect 25317 11305 25329 11339
rect 25363 11336 25375 11339
rect 26050 11336 26056 11348
rect 25363 11308 26056 11336
rect 25363 11305 25375 11308
rect 25317 11299 25375 11305
rect 26050 11296 26056 11308
rect 26108 11296 26114 11348
rect 20548 11240 22692 11268
rect 20441 11231 20499 11237
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18414 11200 18420 11212
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 21450 11200 21456 11212
rect 18800 11172 21456 11200
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16390 11132 16396 11144
rect 16347 11104 16396 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 18800 11132 18828 11172
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 21634 11160 21640 11212
rect 21692 11160 21698 11212
rect 22186 11160 22192 11212
rect 22244 11160 22250 11212
rect 17635 11104 18828 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 16960 11064 16988 11095
rect 18874 11092 18880 11144
rect 18932 11092 18938 11144
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11101 19395 11135
rect 19337 11095 19395 11101
rect 17126 11064 17132 11076
rect 16960 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11064 17190 11076
rect 18322 11064 18328 11076
rect 17184 11036 18328 11064
rect 17184 11024 17190 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18782 11024 18788 11076
rect 18840 11064 18846 11076
rect 19352 11064 19380 11095
rect 19518 11092 19524 11144
rect 19576 11092 19582 11144
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 19944 11104 19993 11132
rect 19944 11092 19950 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 22664 11141 22692 11240
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24581 11271 24639 11277
rect 24581 11268 24593 11271
rect 23532 11240 24593 11268
rect 23532 11228 23538 11240
rect 24581 11237 24593 11240
rect 24627 11237 24639 11271
rect 24581 11231 24639 11237
rect 25133 11271 25191 11277
rect 25133 11237 25145 11271
rect 25179 11268 25191 11271
rect 25866 11268 25872 11280
rect 25179 11240 25872 11268
rect 25179 11237 25191 11240
rect 25133 11231 25191 11237
rect 25866 11228 25872 11240
rect 25924 11228 25930 11280
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24854 11200 24860 11212
rect 23891 11172 24860 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 20128 11104 21189 11132
rect 20128 11092 20134 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 22796 11104 24777 11132
rect 22796 11092 22802 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 18840 11036 19380 11064
rect 18840 11024 18846 11036
rect 18690 10956 18696 11008
rect 18748 10956 18754 11008
rect 19352 10996 19380 11036
rect 20165 11067 20223 11073
rect 20165 11033 20177 11067
rect 20211 11064 20223 11067
rect 20530 11064 20536 11076
rect 20211 11036 20536 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 24302 11024 24308 11076
rect 24360 11064 24366 11076
rect 25409 11067 25467 11073
rect 25409 11064 25421 11067
rect 24360 11036 25421 11064
rect 24360 11024 24366 11036
rect 25409 11033 25421 11036
rect 25455 11033 25467 11067
rect 25409 11027 25467 11033
rect 20717 10999 20775 11005
rect 20717 10996 20729 10999
rect 19352 10968 20729 10996
rect 20717 10965 20729 10968
rect 20763 10996 20775 10999
rect 20806 10996 20812 11008
rect 20763 10968 20812 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20806 10956 20812 10968
rect 20864 10996 20870 11008
rect 21450 10996 21456 11008
rect 20864 10968 21456 10996
rect 20864 10956 20870 10968
rect 21450 10956 21456 10968
rect 21508 10996 21514 11008
rect 22281 10999 22339 11005
rect 22281 10996 22293 10999
rect 21508 10968 22293 10996
rect 21508 10956 21514 10968
rect 22281 10965 22293 10968
rect 22327 10965 22339 10999
rect 22281 10959 22339 10965
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15712 10764 15761 10792
rect 15712 10752 15718 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 16390 10752 16396 10804
rect 16448 10752 16454 10804
rect 17126 10752 17132 10804
rect 17184 10752 17190 10804
rect 18046 10752 18052 10804
rect 18104 10752 18110 10804
rect 19702 10792 19708 10804
rect 18892 10764 19708 10792
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10656 17003 10659
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 16991 10628 18245 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 18233 10625 18245 10628
rect 18279 10656 18291 10659
rect 18506 10656 18512 10668
rect 18279 10628 18512 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 18892 10665 18920 10764
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 21542 10792 21548 10804
rect 20128 10764 21548 10792
rect 20128 10752 20134 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 22554 10792 22560 10804
rect 22066 10764 22560 10792
rect 20165 10683 20223 10689
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 22066 10724 22094 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 21048 10696 22094 10724
rect 23293 10727 23351 10733
rect 21048 10684 21054 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10656 19579 10659
rect 20070 10656 20076 10668
rect 19567 10628 20076 10656
rect 19567 10625 19579 10628
rect 19521 10619 19579 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20165 10649 20177 10683
rect 20211 10680 20223 10683
rect 20211 10656 20300 10680
rect 20346 10656 20352 10668
rect 20211 10652 20352 10656
rect 20211 10649 20223 10652
rect 20165 10643 20223 10649
rect 20272 10628 20352 10652
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20809 10659 20867 10665
rect 20809 10656 20821 10659
rect 20772 10628 20821 10656
rect 20772 10616 20778 10628
rect 20809 10625 20821 10628
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 22002 10656 22008 10668
rect 21499 10628 22008 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 17405 10591 17463 10597
rect 17405 10557 17417 10591
rect 17451 10588 17463 10591
rect 20162 10588 20168 10600
rect 17451 10560 20168 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 22112 10588 22140 10619
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 21692 10560 22140 10588
rect 21692 10548 21698 10560
rect 24670 10548 24676 10600
rect 24728 10548 24734 10600
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 17828 10492 18705 10520
rect 17828 10480 17834 10492
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 19981 10523 20039 10529
rect 19981 10489 19993 10523
rect 20027 10520 20039 10523
rect 23934 10520 23940 10532
rect 20027 10492 23940 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 19334 10412 19340 10464
rect 19392 10412 19398 10464
rect 19702 10412 19708 10464
rect 19760 10452 19766 10464
rect 20346 10452 20352 10464
rect 19760 10424 20352 10452
rect 19760 10412 19766 10424
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 20806 10452 20812 10464
rect 20671 10424 20812 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 19702 10248 19708 10260
rect 17451 10220 19708 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 21634 10248 21640 10260
rect 20272 10220 21640 10248
rect 16666 10140 16672 10192
rect 16724 10180 16730 10192
rect 20272 10180 20300 10220
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 21876 10220 24593 10248
rect 21876 10208 21882 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 24581 10211 24639 10217
rect 16724 10152 20300 10180
rect 16724 10140 16730 10152
rect 20714 10140 20720 10192
rect 20772 10140 20778 10192
rect 22738 10140 22744 10192
rect 22796 10180 22802 10192
rect 23109 10183 23167 10189
rect 23109 10180 23121 10183
rect 22796 10152 23121 10180
rect 22796 10140 22802 10152
rect 23109 10149 23121 10152
rect 23155 10180 23167 10183
rect 23155 10152 25176 10180
rect 23155 10149 23167 10152
rect 23109 10143 23167 10149
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 21266 10112 21272 10124
rect 18095 10084 21272 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 23569 10115 23627 10121
rect 23569 10112 23581 10115
rect 22756 10084 23581 10112
rect 17586 10004 17592 10056
rect 17644 10004 17650 10056
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10044 18383 10047
rect 19426 10044 19432 10056
rect 18371 10016 19432 10044
rect 18371 10013 18383 10016
rect 18325 10007 18383 10013
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 19702 10044 19708 10056
rect 19659 10016 19708 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10044 20959 10047
rect 20990 10044 20996 10056
rect 20947 10016 20996 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 22756 10030 22784 10084
rect 23569 10081 23581 10084
rect 23615 10112 23627 10115
rect 24210 10112 24216 10124
rect 23615 10084 24216 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 25148 10121 25176 10152
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10044 24087 10047
rect 24118 10044 24124 10056
rect 24075 10016 24124 10044
rect 24075 10013 24087 10016
rect 24029 10007 24087 10013
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25774 10044 25780 10056
rect 25087 10016 25780 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25774 10004 25780 10016
rect 25832 10004 25838 10056
rect 20073 9979 20131 9985
rect 20073 9945 20085 9979
rect 20119 9976 20131 9979
rect 20119 9948 21128 9976
rect 20119 9945 20131 9948
rect 20073 9939 20131 9945
rect 19429 9911 19487 9917
rect 19429 9877 19441 9911
rect 19475 9908 19487 9911
rect 19518 9908 19524 9920
rect 19475 9880 19524 9908
rect 19475 9877 19487 9880
rect 19429 9871 19487 9877
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 21100 9908 21128 9948
rect 21174 9936 21180 9988
rect 21232 9976 21238 9988
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21232 9948 21649 9976
rect 21232 9936 21238 9948
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 21637 9939 21695 9945
rect 22940 9948 24961 9976
rect 22940 9908 22968 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 21100 9880 22968 9908
rect 23842 9868 23848 9920
rect 23900 9868 23906 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 19702 9664 19708 9716
rect 19760 9704 19766 9716
rect 21269 9707 21327 9713
rect 21269 9704 21281 9707
rect 19760 9676 21281 9704
rect 19760 9664 19766 9676
rect 21269 9673 21281 9676
rect 21315 9704 21327 9707
rect 22094 9704 22100 9716
rect 21315 9676 22100 9704
rect 21315 9673 21327 9676
rect 21269 9667 21327 9673
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19484 9608 22140 9636
rect 19484 9596 19490 9608
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 8536 9540 18245 9568
rect 8536 9528 8542 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18874 9528 18880 9580
rect 18932 9528 18938 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 20162 9528 20168 9580
rect 20220 9528 20226 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20272 9540 20913 9568
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 20272 9500 20300 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21450 9528 21456 9580
rect 21508 9528 21514 9580
rect 21637 9571 21695 9577
rect 21637 9537 21649 9571
rect 21683 9568 21695 9571
rect 21726 9568 21732 9580
rect 21683 9540 21732 9568
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 22112 9577 22140 9608
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 17276 9472 20300 9500
rect 17276 9460 17282 9472
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9432 18107 9435
rect 18598 9432 18604 9444
rect 18095 9404 18604 9432
rect 18095 9401 18107 9404
rect 18049 9395 18107 9401
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 19337 9435 19395 9441
rect 19337 9401 19349 9435
rect 19383 9432 19395 9435
rect 19426 9432 19432 9444
rect 19383 9404 19432 9432
rect 19383 9401 19395 9404
rect 19337 9395 19395 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 20717 9435 20775 9441
rect 20717 9401 20729 9435
rect 20763 9432 20775 9435
rect 22830 9432 22836 9444
rect 20763 9404 22836 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 15988 9336 18705 9364
rect 15988 9324 15994 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 18693 9327 18751 9333
rect 19981 9367 20039 9373
rect 19981 9333 19993 9367
rect 20027 9364 20039 9367
rect 20990 9364 20996 9376
rect 20027 9336 20996 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 14918 9160 14924 9172
rect 11839 9132 14924 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 19576 9132 20913 9160
rect 19576 9120 19582 9132
rect 20901 9129 20913 9132
rect 20947 9160 20959 9163
rect 20947 9132 22692 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19444 9064 21281 9092
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 19444 9033 19472 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 22554 9092 22560 9104
rect 21269 9055 21327 9061
rect 21376 9064 22560 9092
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 8993 19487 9027
rect 21376 9024 21404 9064
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 22664 9092 22692 9132
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 25133 9163 25191 9169
rect 25133 9160 25145 9163
rect 24176 9132 25145 9160
rect 24176 9120 24182 9132
rect 25133 9129 25145 9132
rect 25179 9129 25191 9163
rect 25133 9123 25191 9129
rect 25409 9163 25467 9169
rect 25409 9129 25421 9163
rect 25455 9160 25467 9163
rect 26234 9160 26240 9172
rect 25455 9132 26240 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 26418 9092 26424 9104
rect 22664 9064 26424 9092
rect 26418 9052 26424 9064
rect 26476 9052 26482 9104
rect 19429 8987 19487 8993
rect 19628 8996 21404 9024
rect 22005 9027 22063 9033
rect 18874 8916 18880 8968
rect 18932 8956 18938 8968
rect 19061 8959 19119 8965
rect 19061 8956 19073 8959
rect 18932 8928 19073 8956
rect 18932 8916 18938 8928
rect 19061 8925 19073 8928
rect 19107 8956 19119 8959
rect 19628 8956 19656 8996
rect 22005 8993 22017 9027
rect 22051 9024 22063 9027
rect 23658 9024 23664 9036
rect 22051 8996 23664 9024
rect 22051 8993 22063 8996
rect 22005 8987 22063 8993
rect 23658 8984 23664 8996
rect 23716 8984 23722 9036
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24854 9024 24860 9036
rect 23891 8996 24860 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 19107 8928 19656 8956
rect 19705 8959 19763 8965
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9364 8860 10333 8888
rect 9364 8848 9370 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12069 8891 12127 8897
rect 12069 8888 12081 8891
rect 11546 8860 12081 8888
rect 10321 8851 10379 8857
rect 12069 8857 12081 8860
rect 12115 8888 12127 8891
rect 12526 8888 12532 8900
rect 12115 8860 12532 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 19720 8888 19748 8919
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 20533 8959 20591 8965
rect 20533 8956 20545 8959
rect 19944 8928 20545 8956
rect 19944 8916 19950 8928
rect 20533 8925 20545 8928
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 21082 8916 21088 8968
rect 21140 8956 21146 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21140 8928 21465 8956
rect 21140 8916 21146 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 21692 8928 22661 8956
rect 21692 8916 21698 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 19720 8860 21036 8888
rect 21008 8820 21036 8860
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 24673 8891 24731 8897
rect 24673 8888 24685 8891
rect 22152 8860 24685 8888
rect 22152 8848 22158 8860
rect 24673 8857 24685 8860
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 24857 8891 24915 8897
rect 24857 8857 24869 8891
rect 24903 8888 24915 8891
rect 25038 8888 25044 8900
rect 24903 8860 25044 8888
rect 24903 8857 24915 8860
rect 24857 8851 24915 8857
rect 25038 8848 25044 8860
rect 25096 8848 25102 8900
rect 23842 8820 23848 8832
rect 21008 8792 23848 8820
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 19610 8616 19616 8628
rect 19475 8588 19616 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 20898 8576 20904 8628
rect 20956 8616 20962 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 20956 8588 21373 8616
rect 20956 8576 20962 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 19208 8520 20944 8548
rect 19208 8508 19214 8520
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 20916 8489 20944 8520
rect 20990 8508 20996 8560
rect 21048 8548 21054 8560
rect 23293 8551 23351 8557
rect 21048 8520 22232 8548
rect 21048 8508 21054 8520
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 15344 8452 19625 8480
rect 15344 8440 15350 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 20901 8483 20959 8489
rect 20901 8449 20913 8483
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21910 8480 21916 8492
rect 21315 8452 21916 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 20272 8412 20300 8443
rect 21284 8412 21312 8443
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22204 8480 22232 8520
rect 23293 8517 23305 8551
rect 23339 8548 23351 8551
rect 24854 8548 24860 8560
rect 23339 8520 24860 8548
rect 23339 8517 23351 8520
rect 23293 8511 23351 8517
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22204 8452 23949 8480
rect 22097 8443 22155 8449
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 24946 8480 24952 8492
rect 23937 8443 23995 8449
rect 24044 8452 24952 8480
rect 20272 8384 21312 8412
rect 22112 8412 22140 8443
rect 24044 8412 24072 8452
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 22112 8384 24072 8412
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 16264 8316 20085 8344
rect 16264 8304 16270 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 21726 8344 21732 8356
rect 20763 8316 21732 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 24026 8276 24032 8288
rect 21600 8248 24032 8276
rect 21600 8236 21606 8248
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 22005 8075 22063 8081
rect 22005 8041 22017 8075
rect 22051 8072 22063 8075
rect 22094 8072 22100 8084
rect 22051 8044 22100 8072
rect 22051 8041 22063 8044
rect 22005 8035 22063 8041
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 21361 8007 21419 8013
rect 21361 7973 21373 8007
rect 21407 8004 21419 8007
rect 23566 8004 23572 8016
rect 21407 7976 23572 8004
rect 21407 7973 21419 7976
rect 21361 7967 21419 7973
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 25590 8004 25596 8016
rect 23676 7976 25596 8004
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 23676 7936 23704 7976
rect 25590 7964 25596 7976
rect 25648 7964 25654 8016
rect 19852 7908 22232 7936
rect 19852 7896 19858 7908
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 18748 7840 20913 7868
rect 18748 7828 18754 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21542 7828 21548 7880
rect 21600 7828 21606 7880
rect 22204 7877 22232 7908
rect 22480 7908 23704 7936
rect 23845 7939 23903 7945
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 20073 7803 20131 7809
rect 20073 7769 20085 7803
rect 20119 7800 20131 7803
rect 22480 7800 22508 7908
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24946 7936 24952 7948
rect 23891 7908 24952 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 22879 7840 24164 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 20119 7772 22508 7800
rect 24136 7800 24164 7840
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24544 7840 24869 7868
rect 24544 7828 24550 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 25682 7800 25688 7812
rect 24136 7772 25688 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 25682 7760 25688 7772
rect 25740 7760 25746 7812
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 23532 7704 24685 7732
rect 23532 7692 23538 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 23293 7463 23351 7469
rect 20772 7432 22416 7460
rect 20772 7420 20778 7432
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20312 7364 20821 7392
rect 20312 7352 20318 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22388 7392 22416 7432
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 22388 7364 23949 7392
rect 22281 7355 22339 7361
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 25314 7392 25320 7404
rect 23937 7355 23995 7361
rect 24044 7364 25320 7392
rect 22296 7324 22324 7355
rect 24044 7324 24072 7364
rect 25314 7352 25320 7364
rect 25372 7352 25378 7404
rect 22296 7296 24072 7324
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 20671 7228 22094 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 22066 7188 22094 7228
rect 23290 7188 23296 7200
rect 22066 7160 23296 7188
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 22005 6851 22063 6857
rect 19392 6820 21496 6848
rect 19392 6808 19398 6820
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 21468 6789 21496 6820
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 23750 6848 23756 6860
rect 22051 6820 23756 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 23845 6851 23903 6857
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24854 6848 24860 6860
rect 23891 6820 24860 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 22664 6712 22692 6743
rect 22830 6740 22836 6792
rect 22888 6780 22894 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 22888 6752 24685 6780
rect 22888 6740 22894 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 20640 6684 22692 6712
rect 24857 6715 24915 6721
rect 20640 6653 20668 6684
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25038 6712 25044 6724
rect 24903 6684 25044 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6644 21327 6647
rect 21634 6644 21640 6656
rect 21315 6616 21640 6644
rect 21315 6613 21327 6616
rect 21269 6607 21327 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 21545 6443 21603 6449
rect 21545 6440 21557 6443
rect 21508 6412 21557 6440
rect 21508 6400 21514 6412
rect 21545 6409 21557 6412
rect 21591 6409 21603 6443
rect 24946 6440 24952 6452
rect 21545 6403 21603 6409
rect 22296 6412 24952 6440
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 22296 6313 22324 6412
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 25498 6304 25504 6316
rect 24167 6276 25504 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 25498 6264 25504 6276
rect 25556 6264 25562 6316
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 22005 5899 22063 5905
rect 22005 5896 22017 5899
rect 15252 5868 22017 5896
rect 15252 5856 15258 5868
rect 22005 5865 22017 5868
rect 22051 5865 22063 5899
rect 22005 5859 22063 5865
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 24578 5828 24584 5840
rect 21407 5800 24584 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 21726 5720 21732 5772
rect 21784 5760 21790 5772
rect 21784 5732 24900 5760
rect 21784 5720 21790 5732
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21818 5692 21824 5704
rect 21591 5664 21824 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5692 22891 5695
rect 23474 5692 23480 5704
rect 22879 5664 23480 5692
rect 22879 5661 22891 5664
rect 22833 5655 22891 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 24872 5701 24900 5732
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 23532 5528 24685 5556
rect 23532 5516 23538 5528
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 23293 5287 23351 5293
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 23382 5216 23388 5228
rect 22327 5188 23388 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23900 5188 23949 5216
rect 23900 5176 23906 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 19058 4768 19064 4820
rect 19116 4808 19122 4820
rect 22005 4811 22063 4817
rect 22005 4808 22017 4811
rect 19116 4780 22017 4808
rect 19116 4768 19122 4780
rect 22005 4777 22017 4780
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22189 4607 22247 4613
rect 22189 4604 22201 4607
rect 21775 4576 22201 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22189 4573 22201 4576
rect 22235 4604 22247 4607
rect 22278 4604 22284 4616
rect 22235 4576 22284 4604
rect 22235 4573 22247 4576
rect 22189 4567 22247 4573
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 23290 4564 23296 4616
rect 23348 4604 23354 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 23348 4576 24869 4604
rect 23348 4564 23354 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 22336 4440 24685 4468
rect 22336 4428 22342 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 23952 4168 25176 4196
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 23952 4137 23980 4168
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 20036 4100 20085 4128
rect 20036 4088 20042 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23937 4131 23995 4137
rect 22327 4100 23428 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20162 4060 20168 4072
rect 19024 4032 20168 4060
rect 19024 4020 19030 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22094 4060 22100 4072
rect 21315 4032 22100 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23400 4060 23428 4100
rect 23937 4097 23949 4131
rect 23983 4097 23995 4131
rect 25038 4128 25044 4140
rect 23937 4091 23995 4097
rect 24044 4100 25044 4128
rect 24044 4060 24072 4100
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25148 4128 25176 4168
rect 26602 4128 26608 4140
rect 25148 4100 26608 4128
rect 26602 4088 26608 4100
rect 26660 4088 26666 4140
rect 23400 4032 24072 4060
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7466 3516 7472 3528
rect 6871 3488 7472 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20588 3488 20821 3516
rect 20588 3476 20594 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23474 3516 23480 3528
rect 22879 3488 23480 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 24636 3488 24777 3516
rect 24636 3476 24642 3488
rect 24765 3485 24777 3488
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24946 3448 24952 3460
rect 23891 3420 24952 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 7248 3352 7481 3380
rect 7248 3340 7254 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 24578 3340 24584 3392
rect 24636 3340 24642 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 7466 3136 7472 3188
rect 7524 3136 7530 3188
rect 19242 3068 19248 3120
rect 19300 3108 19306 3120
rect 23293 3111 23351 3117
rect 19300 3080 20116 3108
rect 19300 3068 19306 3080
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19794 3040 19800 3052
rect 18463 3012 19800 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 20088 3049 20116 3080
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25130 3068 25136 3120
rect 25188 3068 25194 3120
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3040 24179 3043
rect 25406 3040 25412 3052
rect 24167 3012 25412 3040
rect 24167 3009 24179 3012
rect 24121 3003 24179 3009
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19518 2972 19524 2984
rect 19475 2944 19524 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 6549 2839 6607 2845
rect 6549 2805 6561 2839
rect 6595 2836 6607 2839
rect 6730 2836 6736 2848
rect 6595 2808 6736 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 25222 2836 25228 2848
rect 19852 2808 25228 2836
rect 19852 2796 19858 2808
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 8662 2632 8668 2644
rect 6595 2604 8668 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 19794 2592 19800 2644
rect 19852 2592 19858 2644
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 6886 2468 7849 2496
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 6886 2428 6914 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 19518 2456 19524 2508
rect 19576 2496 19582 2508
rect 22738 2496 22744 2508
rect 19576 2468 22744 2496
rect 19576 2456 19582 2468
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 6779 2400 6914 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 22646 2428 22652 2440
rect 20303 2400 22652 2428
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2428 22891 2431
rect 24578 2428 24584 2440
rect 22879 2400 24584 2428
rect 22879 2397 22891 2400
rect 22833 2391 22891 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23382 2360 23388 2372
rect 21315 2332 23388 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 23382 2320 23388 2332
rect 23440 2320 23446 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 3056 26392 3108 26444
rect 3332 26392 3384 26444
rect 2504 26188 2556 26240
rect 12624 26188 12676 26240
rect 9128 25032 9180 25084
rect 20904 25032 20956 25084
rect 4804 24964 4856 25016
rect 18696 24964 18748 25016
rect 10232 24896 10284 24948
rect 22376 24896 22428 24948
rect 7748 24828 7800 24880
rect 18420 24828 18472 24880
rect 20536 24828 20588 24880
rect 23388 24828 23440 24880
rect 2412 24760 2464 24812
rect 15200 24760 15252 24812
rect 17408 24760 17460 24812
rect 17776 24760 17828 24812
rect 24124 24760 24176 24812
rect 5816 24692 5868 24744
rect 7288 24692 7340 24744
rect 10416 24692 10468 24744
rect 19248 24692 19300 24744
rect 2320 24624 2372 24676
rect 7104 24624 7156 24676
rect 14832 24624 14884 24676
rect 22836 24624 22888 24676
rect 5908 24556 5960 24608
rect 10324 24556 10376 24608
rect 11704 24556 11756 24608
rect 14556 24556 14608 24608
rect 22652 24556 22704 24608
rect 23112 24556 23164 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 3976 24395 4028 24404
rect 3976 24361 3985 24395
rect 3985 24361 4019 24395
rect 4019 24361 4028 24395
rect 3976 24352 4028 24361
rect 6736 24352 6788 24404
rect 9128 24395 9180 24404
rect 9128 24361 9137 24395
rect 9137 24361 9171 24395
rect 9171 24361 9180 24395
rect 9128 24352 9180 24361
rect 11060 24284 11112 24336
rect 6460 24216 6512 24268
rect 9680 24216 9732 24268
rect 11244 24216 11296 24268
rect 3884 24148 3936 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 6736 24191 6788 24200
rect 6736 24157 6745 24191
rect 6745 24157 6779 24191
rect 6779 24157 6788 24191
rect 6736 24148 6788 24157
rect 7288 24191 7340 24200
rect 7288 24157 7297 24191
rect 7297 24157 7331 24191
rect 7331 24157 7340 24191
rect 7288 24148 7340 24157
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 1584 24123 1636 24132
rect 1584 24089 1593 24123
rect 1593 24089 1627 24123
rect 1627 24089 1636 24123
rect 1584 24080 1636 24089
rect 8668 24080 8720 24132
rect 2320 24012 2372 24064
rect 6368 24012 6420 24064
rect 7472 24012 7524 24064
rect 9956 24148 10008 24200
rect 17316 24352 17368 24404
rect 12348 24284 12400 24336
rect 22100 24352 22152 24404
rect 12440 24216 12492 24268
rect 17408 24216 17460 24268
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18512 24259 18564 24268
rect 18512 24225 18521 24259
rect 18521 24225 18555 24259
rect 18555 24225 18564 24259
rect 18512 24216 18564 24225
rect 20720 24216 20772 24268
rect 22560 24216 22612 24268
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 14004 24148 14056 24200
rect 9588 24080 9640 24132
rect 15844 24148 15896 24200
rect 9864 24012 9916 24064
rect 17592 24080 17644 24132
rect 18236 24080 18288 24132
rect 19156 24080 19208 24132
rect 16212 24055 16264 24064
rect 16212 24021 16221 24055
rect 16221 24021 16255 24055
rect 16255 24021 16264 24055
rect 16212 24012 16264 24021
rect 16396 24055 16448 24064
rect 16396 24021 16405 24055
rect 16405 24021 16439 24055
rect 16439 24021 16448 24055
rect 16396 24012 16448 24021
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 17224 24055 17276 24064
rect 17224 24021 17233 24055
rect 17233 24021 17267 24055
rect 17267 24021 17276 24055
rect 17224 24012 17276 24021
rect 18972 24012 19024 24064
rect 19340 24055 19392 24064
rect 19340 24021 19349 24055
rect 19349 24021 19383 24055
rect 19383 24021 19392 24055
rect 19340 24012 19392 24021
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 23848 24216 23900 24268
rect 25044 24191 25096 24200
rect 25044 24157 25053 24191
rect 25053 24157 25087 24191
rect 25087 24157 25096 24191
rect 25044 24148 25096 24157
rect 22468 24080 22520 24132
rect 23940 24080 23992 24132
rect 19524 24012 19576 24064
rect 20628 24055 20680 24064
rect 20628 24021 20637 24055
rect 20637 24021 20671 24055
rect 20671 24021 20680 24055
rect 20628 24012 20680 24021
rect 22008 24012 22060 24064
rect 22928 24012 22980 24064
rect 24124 24012 24176 24064
rect 24860 24012 24912 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 2320 23851 2372 23860
rect 2320 23817 2329 23851
rect 2329 23817 2363 23851
rect 2363 23817 2372 23851
rect 2320 23808 2372 23817
rect 6828 23808 6880 23860
rect 5356 23740 5408 23792
rect 5816 23783 5868 23792
rect 5816 23749 5825 23783
rect 5825 23749 5859 23783
rect 5859 23749 5868 23783
rect 5816 23740 5868 23749
rect 8024 23808 8076 23860
rect 9312 23808 9364 23860
rect 11704 23808 11756 23860
rect 14004 23808 14056 23860
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 3608 23672 3660 23724
rect 6736 23672 6788 23724
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 6000 23604 6052 23656
rect 10140 23740 10192 23792
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 10968 23740 11020 23792
rect 20628 23808 20680 23860
rect 22928 23808 22980 23860
rect 25504 23808 25556 23860
rect 15200 23783 15252 23792
rect 15200 23749 15209 23783
rect 15209 23749 15243 23783
rect 15243 23749 15252 23783
rect 15200 23740 15252 23749
rect 15384 23783 15436 23792
rect 15384 23749 15393 23783
rect 15393 23749 15427 23783
rect 15427 23749 15436 23783
rect 15384 23740 15436 23749
rect 16120 23740 16172 23792
rect 17408 23740 17460 23792
rect 5908 23536 5960 23588
rect 5448 23468 5500 23520
rect 9772 23672 9824 23724
rect 8024 23604 8076 23656
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 15844 23672 15896 23724
rect 10048 23604 10100 23656
rect 11980 23604 12032 23656
rect 12716 23536 12768 23588
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 16304 23604 16356 23656
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 17316 23672 17368 23681
rect 18420 23740 18472 23792
rect 18880 23740 18932 23792
rect 23940 23740 23992 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 17776 23604 17828 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 20720 23672 20772 23724
rect 19984 23604 20036 23656
rect 20628 23647 20680 23656
rect 20628 23613 20637 23647
rect 20637 23613 20671 23647
rect 20671 23613 20680 23647
rect 20628 23604 20680 23613
rect 17960 23536 18012 23588
rect 22100 23604 22152 23656
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 23296 23604 23348 23656
rect 24308 23604 24360 23656
rect 9220 23468 9272 23520
rect 10968 23468 11020 23520
rect 12624 23468 12676 23520
rect 13360 23468 13412 23520
rect 16672 23468 16724 23520
rect 16856 23511 16908 23520
rect 16856 23477 16865 23511
rect 16865 23477 16899 23511
rect 16899 23477 16908 23511
rect 16856 23468 16908 23477
rect 17224 23468 17276 23520
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 21364 23468 21416 23520
rect 25872 23536 25924 23588
rect 22376 23468 22428 23520
rect 22560 23468 22612 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 3608 23264 3660 23316
rect 3976 23264 4028 23316
rect 6736 23264 6788 23316
rect 9128 23264 9180 23316
rect 13268 23264 13320 23316
rect 1952 23196 2004 23248
rect 7012 23196 7064 23248
rect 4620 23128 4672 23180
rect 7656 23128 7708 23180
rect 9404 23196 9456 23248
rect 15660 23264 15712 23316
rect 16856 23264 16908 23316
rect 8668 23128 8720 23180
rect 16304 23196 16356 23248
rect 17040 23196 17092 23248
rect 19432 23196 19484 23248
rect 23388 23239 23440 23248
rect 23388 23205 23397 23239
rect 23397 23205 23431 23239
rect 23431 23205 23440 23239
rect 23388 23196 23440 23205
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11612 23128 11664 23180
rect 12256 23128 12308 23180
rect 14924 23128 14976 23180
rect 18512 23128 18564 23180
rect 18696 23171 18748 23180
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 21180 23128 21232 23180
rect 22284 23128 22336 23180
rect 23296 23128 23348 23180
rect 4344 23103 4396 23112
rect 4344 23069 4353 23103
rect 4353 23069 4387 23103
rect 4387 23069 4396 23103
rect 4344 23060 4396 23069
rect 5540 23060 5592 23112
rect 6276 23060 6328 23112
rect 9588 23060 9640 23112
rect 5816 22992 5868 23044
rect 7564 22992 7616 23044
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14188 23060 14240 23112
rect 16396 23060 16448 23112
rect 16672 23060 16724 23112
rect 10048 22992 10100 23044
rect 13912 22992 13964 23044
rect 14004 22992 14056 23044
rect 14556 22992 14608 23044
rect 15384 22992 15436 23044
rect 17868 23060 17920 23112
rect 18052 23060 18104 23112
rect 19340 23060 19392 23112
rect 24768 23060 24820 23112
rect 12532 22924 12584 22976
rect 12808 22924 12860 22976
rect 13544 22967 13596 22976
rect 13544 22933 13553 22967
rect 13553 22933 13587 22967
rect 13587 22933 13596 22967
rect 13544 22924 13596 22933
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 15660 22924 15712 22976
rect 16304 22924 16356 22976
rect 16580 22924 16632 22976
rect 17224 22967 17276 22976
rect 17224 22933 17233 22967
rect 17233 22933 17267 22967
rect 17267 22933 17276 22967
rect 17224 22924 17276 22933
rect 18788 22992 18840 23044
rect 19984 22992 20036 23044
rect 20168 22992 20220 23044
rect 21916 23035 21968 23044
rect 21916 23001 21925 23035
rect 21925 23001 21959 23035
rect 21959 23001 21968 23035
rect 21916 22992 21968 23001
rect 17776 22924 17828 22976
rect 18696 22924 18748 22976
rect 20720 22924 20772 22976
rect 21824 22924 21876 22976
rect 23756 22992 23808 23044
rect 25320 22992 25372 23044
rect 23572 22924 23624 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1492 22720 1544 22772
rect 6920 22720 6972 22772
rect 7104 22720 7156 22772
rect 4252 22652 4304 22704
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 8392 22652 8444 22704
rect 4528 22584 4580 22636
rect 5632 22584 5684 22636
rect 6736 22584 6788 22636
rect 3608 22516 3660 22568
rect 4160 22448 4212 22500
rect 12256 22720 12308 22772
rect 12716 22720 12768 22772
rect 13268 22720 13320 22772
rect 14556 22720 14608 22772
rect 14740 22720 14792 22772
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 11152 22652 11204 22704
rect 10784 22584 10836 22636
rect 9036 22516 9088 22568
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 12440 22516 12492 22568
rect 10876 22448 10928 22500
rect 13360 22448 13412 22500
rect 2228 22423 2280 22432
rect 2228 22389 2237 22423
rect 2237 22389 2271 22423
rect 2271 22389 2280 22423
rect 2228 22380 2280 22389
rect 5816 22380 5868 22432
rect 10048 22380 10100 22432
rect 11244 22380 11296 22432
rect 12256 22380 12308 22432
rect 12992 22380 13044 22432
rect 14188 22652 14240 22704
rect 15292 22652 15344 22704
rect 16488 22720 16540 22772
rect 16028 22652 16080 22704
rect 16212 22652 16264 22704
rect 17868 22720 17920 22772
rect 18512 22720 18564 22772
rect 19248 22763 19300 22772
rect 19248 22729 19257 22763
rect 19257 22729 19291 22763
rect 19291 22729 19300 22763
rect 19248 22720 19300 22729
rect 15568 22584 15620 22636
rect 16580 22584 16632 22636
rect 17040 22652 17092 22704
rect 18420 22652 18472 22704
rect 18880 22584 18932 22636
rect 15752 22516 15804 22568
rect 20628 22584 20680 22636
rect 23756 22720 23808 22772
rect 23940 22720 23992 22772
rect 20168 22516 20220 22568
rect 21088 22516 21140 22568
rect 21824 22516 21876 22568
rect 15200 22448 15252 22500
rect 16396 22448 16448 22500
rect 16856 22448 16908 22500
rect 16304 22380 16356 22432
rect 16672 22380 16724 22432
rect 17684 22380 17736 22432
rect 17776 22380 17828 22432
rect 20996 22448 21048 22500
rect 22100 22448 22152 22500
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 24124 22516 24176 22568
rect 25780 22516 25832 22568
rect 18880 22380 18932 22432
rect 20076 22380 20128 22432
rect 20260 22380 20312 22432
rect 22652 22380 22704 22432
rect 23664 22380 23716 22432
rect 24768 22380 24820 22432
rect 25688 22380 25740 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 2228 22176 2280 22228
rect 1676 22083 1728 22092
rect 1676 22049 1685 22083
rect 1685 22049 1719 22083
rect 1719 22049 1728 22083
rect 1676 22040 1728 22049
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22108 8352 22160
rect 9496 22176 9548 22228
rect 13452 22176 13504 22228
rect 14740 22176 14792 22228
rect 10600 22108 10652 22160
rect 12716 22108 12768 22160
rect 9036 22040 9088 22092
rect 11060 22040 11112 22092
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12440 22040 12492 22049
rect 16304 22108 16356 22160
rect 18880 22176 18932 22228
rect 19432 22176 19484 22228
rect 21272 22176 21324 22228
rect 23848 22176 23900 22228
rect 17684 22108 17736 22160
rect 22376 22108 22428 22160
rect 22652 22108 22704 22160
rect 2688 21972 2740 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4436 21972 4488 22024
rect 6460 21972 6512 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 9496 22015 9548 22024
rect 9496 21981 9505 22015
rect 9505 21981 9539 22015
rect 9539 21981 9548 22015
rect 9496 21972 9548 21981
rect 12072 21972 12124 22024
rect 13452 21972 13504 22024
rect 14188 21972 14240 22024
rect 15568 21972 15620 22024
rect 16396 22040 16448 22092
rect 17224 22040 17276 22092
rect 18144 22083 18196 22092
rect 18144 22049 18153 22083
rect 18153 22049 18187 22083
rect 18187 22049 18196 22083
rect 18144 22040 18196 22049
rect 18420 22040 18472 22092
rect 9404 21904 9456 21956
rect 10416 21904 10468 21956
rect 13544 21947 13596 21956
rect 2136 21836 2188 21888
rect 8208 21836 8260 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 10508 21836 10560 21888
rect 13544 21913 13553 21947
rect 13553 21913 13587 21947
rect 13587 21913 13596 21947
rect 13544 21904 13596 21913
rect 12716 21836 12768 21888
rect 13360 21836 13412 21888
rect 14556 21836 14608 21888
rect 18604 21972 18656 22024
rect 19248 21972 19300 22024
rect 19340 21972 19392 22024
rect 22376 21972 22428 22024
rect 23480 22040 23532 22092
rect 25412 22108 25464 22160
rect 24216 21972 24268 22024
rect 16580 21904 16632 21956
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 16948 21879 17000 21888
rect 16948 21845 16957 21879
rect 16957 21845 16991 21879
rect 16991 21845 17000 21879
rect 16948 21836 17000 21845
rect 17776 21904 17828 21956
rect 17868 21836 17920 21888
rect 18144 21836 18196 21888
rect 18512 21836 18564 21888
rect 19524 21947 19576 21956
rect 19524 21913 19533 21947
rect 19533 21913 19567 21947
rect 19567 21913 19576 21947
rect 19524 21904 19576 21913
rect 21088 21904 21140 21956
rect 21916 21904 21968 21956
rect 20076 21836 20128 21888
rect 21640 21836 21692 21888
rect 25136 21904 25188 21956
rect 24492 21836 24544 21888
rect 25596 21836 25648 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 1400 21564 1452 21616
rect 6736 21632 6788 21684
rect 6920 21632 6972 21684
rect 7288 21632 7340 21684
rect 8484 21564 8536 21616
rect 10784 21564 10836 21616
rect 12072 21632 12124 21684
rect 11612 21607 11664 21616
rect 11612 21573 11621 21607
rect 11621 21573 11655 21607
rect 11655 21573 11664 21607
rect 11612 21564 11664 21573
rect 6092 21496 6144 21548
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 10692 21496 10744 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 7288 21428 7340 21480
rect 8300 21428 8352 21480
rect 8576 21428 8628 21480
rect 10876 21428 10928 21480
rect 13728 21632 13780 21684
rect 17316 21632 17368 21684
rect 7932 21360 7984 21412
rect 10600 21360 10652 21412
rect 12348 21360 12400 21412
rect 12440 21360 12492 21412
rect 14280 21564 14332 21616
rect 16488 21564 16540 21616
rect 17776 21632 17828 21684
rect 19064 21632 19116 21684
rect 20720 21632 20772 21684
rect 21364 21632 21416 21684
rect 22192 21632 22244 21684
rect 22284 21632 22336 21684
rect 12808 21471 12860 21480
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 6644 21292 6696 21344
rect 8576 21292 8628 21344
rect 10416 21292 10468 21344
rect 10508 21292 10560 21344
rect 10876 21292 10928 21344
rect 11152 21292 11204 21344
rect 12072 21292 12124 21344
rect 14004 21428 14056 21480
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 16396 21496 16448 21548
rect 15108 21428 15160 21480
rect 15660 21471 15712 21480
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 15936 21428 15988 21480
rect 16304 21428 16356 21480
rect 17500 21564 17552 21616
rect 18512 21564 18564 21616
rect 21456 21607 21508 21616
rect 21456 21573 21465 21607
rect 21465 21573 21499 21607
rect 21499 21573 21508 21607
rect 21456 21564 21508 21573
rect 21640 21564 21692 21616
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 20444 21496 20496 21548
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 22376 21539 22428 21548
rect 22376 21505 22385 21539
rect 22385 21505 22419 21539
rect 22419 21505 22428 21539
rect 22376 21496 22428 21505
rect 17684 21471 17736 21480
rect 17684 21437 17693 21471
rect 17693 21437 17727 21471
rect 17727 21437 17736 21471
rect 17684 21428 17736 21437
rect 13544 21360 13596 21412
rect 13820 21360 13872 21412
rect 17776 21360 17828 21412
rect 13452 21335 13504 21344
rect 13452 21301 13461 21335
rect 13461 21301 13495 21335
rect 13495 21301 13504 21335
rect 13452 21292 13504 21301
rect 15568 21292 15620 21344
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 16580 21292 16632 21344
rect 16764 21292 16816 21344
rect 19432 21428 19484 21480
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 23940 21564 23992 21616
rect 23296 21496 23348 21548
rect 19156 21360 19208 21412
rect 19340 21292 19392 21344
rect 19984 21292 20036 21344
rect 22192 21360 22244 21412
rect 24676 21428 24728 21480
rect 21916 21292 21968 21344
rect 22560 21292 22612 21344
rect 22836 21292 22888 21344
rect 23756 21292 23808 21344
rect 25412 21335 25464 21344
rect 25412 21301 25421 21335
rect 25421 21301 25455 21335
rect 25455 21301 25464 21335
rect 25412 21292 25464 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 5816 21131 5868 21140
rect 5816 21097 5825 21131
rect 5825 21097 5859 21131
rect 5859 21097 5868 21131
rect 5816 21088 5868 21097
rect 9128 21088 9180 21140
rect 2780 21020 2832 21072
rect 5172 21020 5224 21072
rect 4160 20952 4212 21004
rect 5816 20884 5868 20936
rect 6552 20952 6604 21004
rect 8484 21020 8536 21072
rect 9220 20952 9272 21004
rect 10048 20952 10100 21004
rect 12716 21020 12768 21072
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 13728 21088 13780 21140
rect 16856 21088 16908 21140
rect 16764 21020 16816 21072
rect 17040 21020 17092 21072
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 7288 20884 7340 20936
rect 7656 20816 7708 20868
rect 7932 20884 7984 20936
rect 9772 20884 9824 20936
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 11060 20952 11112 21004
rect 12808 20952 12860 21004
rect 13636 20952 13688 21004
rect 14096 20952 14148 21004
rect 13176 20884 13228 20936
rect 3976 20748 4028 20800
rect 8852 20748 8904 20800
rect 10600 20748 10652 20800
rect 12900 20816 12952 20868
rect 13452 20816 13504 20868
rect 13544 20859 13596 20868
rect 13544 20825 13553 20859
rect 13553 20825 13587 20859
rect 13587 20825 13596 20859
rect 13544 20816 13596 20825
rect 14832 20884 14884 20936
rect 15936 20927 15988 20936
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 12440 20748 12492 20800
rect 13360 20748 13412 20800
rect 13728 20748 13780 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 14648 20816 14700 20868
rect 17776 21088 17828 21140
rect 17776 20952 17828 21004
rect 22376 21088 22428 21140
rect 22468 21088 22520 21140
rect 18788 21020 18840 21072
rect 21180 21063 21232 21072
rect 21180 21029 21189 21063
rect 21189 21029 21223 21063
rect 21223 21029 21232 21063
rect 21180 21020 21232 21029
rect 18696 20952 18748 21004
rect 21640 20952 21692 21004
rect 23940 21063 23992 21072
rect 23940 21029 23949 21063
rect 23949 21029 23983 21063
rect 23983 21029 23992 21063
rect 23940 21020 23992 21029
rect 24124 21020 24176 21072
rect 24400 21020 24452 21072
rect 16948 20884 17000 20936
rect 17868 20884 17920 20936
rect 18420 20884 18472 20936
rect 19340 20884 19392 20936
rect 21916 20884 21968 20936
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22100 20884 22152 20893
rect 17316 20816 17368 20868
rect 21088 20816 21140 20868
rect 15384 20748 15436 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 15936 20748 15988 20800
rect 16212 20748 16264 20800
rect 16396 20748 16448 20800
rect 19248 20748 19300 20800
rect 19800 20748 19852 20800
rect 21364 20748 21416 20800
rect 23664 20952 23716 21004
rect 22376 20884 22428 20936
rect 23112 20884 23164 20936
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 24676 20884 24728 20936
rect 23388 20816 23440 20868
rect 23112 20748 23164 20800
rect 24860 20748 24912 20800
rect 25964 20748 26016 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 26056 20680 26108 20732
rect 26424 20680 26476 20732
rect 6828 20544 6880 20596
rect 7288 20544 7340 20596
rect 10048 20544 10100 20596
rect 10968 20544 11020 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 13176 20587 13228 20596
rect 13176 20553 13185 20587
rect 13185 20553 13219 20587
rect 13219 20553 13228 20587
rect 13176 20544 13228 20553
rect 13820 20544 13872 20596
rect 14188 20544 14240 20596
rect 3424 20476 3476 20528
rect 4896 20519 4948 20528
rect 4896 20485 4905 20519
rect 4905 20485 4939 20519
rect 4939 20485 4948 20519
rect 4896 20476 4948 20485
rect 5356 20476 5408 20528
rect 5540 20408 5592 20460
rect 7012 20408 7064 20460
rect 9588 20476 9640 20528
rect 10600 20476 10652 20528
rect 11060 20476 11112 20528
rect 11980 20476 12032 20528
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 7932 20340 7984 20392
rect 10508 20340 10560 20392
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 4252 20272 4304 20324
rect 6920 20204 6972 20256
rect 7196 20204 7248 20256
rect 13360 20272 13412 20324
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 11060 20204 11112 20256
rect 12440 20204 12492 20256
rect 12900 20204 12952 20256
rect 15200 20476 15252 20528
rect 15568 20476 15620 20528
rect 17224 20544 17276 20596
rect 18144 20544 18196 20596
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 18880 20544 18932 20596
rect 15476 20408 15528 20460
rect 16488 20408 16540 20460
rect 14556 20340 14608 20392
rect 15016 20340 15068 20392
rect 16764 20340 16816 20392
rect 18236 20340 18288 20392
rect 15108 20272 15160 20324
rect 15844 20204 15896 20256
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 17040 20204 17092 20256
rect 18788 20476 18840 20528
rect 21272 20544 21324 20596
rect 21364 20544 21416 20596
rect 21916 20544 21968 20596
rect 22468 20544 22520 20596
rect 22560 20587 22612 20596
rect 22560 20553 22569 20587
rect 22569 20553 22603 20587
rect 22603 20553 22612 20587
rect 22560 20544 22612 20553
rect 25412 20544 25464 20596
rect 20904 20476 20956 20528
rect 23664 20476 23716 20528
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 24400 20476 24452 20528
rect 22376 20408 22428 20460
rect 23296 20408 23348 20460
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19892 20340 19944 20392
rect 20168 20340 20220 20392
rect 22560 20340 22612 20392
rect 22652 20383 22704 20392
rect 22652 20349 22661 20383
rect 22661 20349 22695 20383
rect 22695 20349 22704 20383
rect 22652 20340 22704 20349
rect 20720 20272 20772 20324
rect 19616 20204 19668 20256
rect 20536 20204 20588 20256
rect 21364 20204 21416 20256
rect 21824 20204 21876 20256
rect 22468 20204 22520 20256
rect 23848 20204 23900 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 7012 20000 7064 20052
rect 11428 20000 11480 20052
rect 15844 20000 15896 20052
rect 17960 20000 18012 20052
rect 18236 20000 18288 20052
rect 20904 20000 20956 20052
rect 23940 20000 23992 20052
rect 7656 19932 7708 19984
rect 7932 19932 7984 19984
rect 11520 19932 11572 19984
rect 13636 19932 13688 19984
rect 14372 19932 14424 19984
rect 2044 19864 2096 19916
rect 5172 19907 5224 19916
rect 5172 19873 5181 19907
rect 5181 19873 5215 19907
rect 5215 19873 5224 19907
rect 5172 19864 5224 19873
rect 6184 19864 6236 19916
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 4896 19796 4948 19848
rect 7472 19864 7524 19916
rect 10784 19864 10836 19916
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 5356 19660 5408 19712
rect 7840 19796 7892 19848
rect 17132 19932 17184 19984
rect 18788 19932 18840 19984
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18236 19907 18288 19916
rect 18236 19873 18245 19907
rect 18245 19873 18279 19907
rect 18279 19873 18288 19907
rect 18236 19864 18288 19873
rect 18696 19907 18748 19916
rect 18696 19873 18705 19907
rect 18705 19873 18739 19907
rect 18739 19873 18748 19907
rect 18696 19864 18748 19873
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 11428 19728 11480 19780
rect 7472 19660 7524 19712
rect 7656 19660 7708 19712
rect 8208 19660 8260 19712
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 11152 19660 11204 19712
rect 12440 19728 12492 19780
rect 14004 19796 14056 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 14556 19796 14608 19848
rect 19156 19932 19208 19984
rect 20628 19975 20680 19984
rect 20628 19941 20637 19975
rect 20637 19941 20671 19975
rect 20671 19941 20680 19975
rect 20628 19932 20680 19941
rect 13268 19728 13320 19780
rect 14924 19728 14976 19780
rect 15016 19728 15068 19780
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 15936 19728 15988 19780
rect 16764 19728 16816 19780
rect 20720 19864 20772 19916
rect 23296 19864 23348 19916
rect 24400 19864 24452 19916
rect 25044 19907 25096 19916
rect 25044 19873 25053 19907
rect 25053 19873 25087 19907
rect 25087 19873 25096 19907
rect 25044 19864 25096 19873
rect 25136 19907 25188 19916
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 25136 19864 25188 19873
rect 20628 19796 20680 19848
rect 23480 19796 23532 19848
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 14464 19660 14516 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 16856 19660 16908 19712
rect 19524 19728 19576 19780
rect 21824 19728 21876 19780
rect 24124 19728 24176 19780
rect 25044 19728 25096 19780
rect 17224 19660 17276 19712
rect 19708 19660 19760 19712
rect 21640 19660 21692 19712
rect 23480 19660 23532 19712
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 24308 19660 24360 19712
rect 24584 19703 24636 19712
rect 24584 19669 24593 19703
rect 24593 19669 24627 19703
rect 24627 19669 24636 19703
rect 24584 19660 24636 19669
rect 26056 19660 26108 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 4620 19456 4672 19508
rect 6276 19456 6328 19508
rect 7288 19456 7340 19508
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 9680 19456 9732 19508
rect 10876 19456 10928 19508
rect 11060 19499 11112 19508
rect 11060 19465 11069 19499
rect 11069 19465 11103 19499
rect 11103 19465 11112 19499
rect 11060 19456 11112 19465
rect 11612 19456 11664 19508
rect 5908 19388 5960 19440
rect 5448 19320 5500 19372
rect 8300 19388 8352 19440
rect 1860 19252 1912 19304
rect 2872 19252 2924 19304
rect 6552 19252 6604 19304
rect 7748 19320 7800 19372
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 8944 19320 8996 19372
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 13820 19456 13872 19508
rect 14004 19456 14056 19508
rect 14648 19456 14700 19508
rect 14924 19499 14976 19508
rect 14924 19465 14933 19499
rect 14933 19465 14967 19499
rect 14967 19465 14976 19499
rect 14924 19456 14976 19465
rect 15568 19456 15620 19508
rect 17040 19456 17092 19508
rect 18144 19456 18196 19508
rect 20996 19456 21048 19508
rect 21180 19456 21232 19508
rect 22376 19499 22428 19508
rect 22376 19465 22385 19499
rect 22385 19465 22419 19499
rect 22419 19465 22428 19499
rect 22376 19456 22428 19465
rect 25136 19456 25188 19508
rect 25320 19456 25372 19508
rect 12624 19388 12676 19440
rect 13268 19388 13320 19440
rect 14280 19388 14332 19440
rect 14464 19320 14516 19372
rect 15200 19320 15252 19372
rect 16580 19388 16632 19440
rect 19432 19388 19484 19440
rect 23572 19388 23624 19440
rect 24124 19388 24176 19440
rect 16488 19320 16540 19372
rect 6736 19295 6788 19304
rect 6736 19261 6745 19295
rect 6745 19261 6779 19295
rect 6779 19261 6788 19295
rect 6736 19252 6788 19261
rect 10784 19252 10836 19304
rect 11796 19252 11848 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 15108 19252 15160 19304
rect 16028 19252 16080 19304
rect 16396 19252 16448 19304
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 17684 19252 17736 19304
rect 6920 19184 6972 19236
rect 3332 19116 3384 19168
rect 8576 19116 8628 19168
rect 9404 19116 9456 19168
rect 15660 19184 15712 19236
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11428 19116 11480 19168
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 12440 19116 12492 19168
rect 13636 19116 13688 19168
rect 14464 19116 14516 19168
rect 14740 19116 14792 19168
rect 16396 19116 16448 19168
rect 21272 19320 21324 19372
rect 21364 19320 21416 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 20352 19252 20404 19304
rect 21088 19184 21140 19236
rect 22008 19252 22060 19304
rect 21732 19184 21784 19236
rect 25228 19252 25280 19304
rect 24676 19184 24728 19236
rect 25044 19184 25096 19236
rect 19708 19116 19760 19168
rect 20352 19116 20404 19168
rect 20996 19116 21048 19168
rect 22192 19116 22244 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 2412 18912 2464 18964
rect 3608 18912 3660 18964
rect 3700 18912 3752 18964
rect 5540 18912 5592 18964
rect 5908 18912 5960 18964
rect 8576 18912 8628 18964
rect 10692 18912 10744 18964
rect 14188 18912 14240 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 6552 18776 6604 18828
rect 7196 18776 7248 18828
rect 7564 18776 7616 18828
rect 7840 18776 7892 18828
rect 23204 18912 23256 18964
rect 25044 18912 25096 18964
rect 9496 18776 9548 18828
rect 10968 18776 11020 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 5080 18708 5132 18760
rect 6184 18708 6236 18760
rect 4252 18640 4304 18692
rect 3240 18615 3292 18624
rect 3240 18581 3249 18615
rect 3249 18581 3283 18615
rect 3283 18581 3292 18615
rect 3240 18572 3292 18581
rect 5724 18640 5776 18692
rect 9128 18708 9180 18760
rect 11796 18708 11848 18760
rect 14740 18776 14792 18828
rect 14924 18844 14976 18896
rect 17868 18844 17920 18896
rect 19064 18844 19116 18896
rect 21640 18844 21692 18896
rect 15016 18776 15068 18828
rect 17684 18776 17736 18828
rect 18328 18776 18380 18828
rect 22468 18776 22520 18828
rect 9312 18640 9364 18692
rect 13820 18708 13872 18760
rect 14924 18708 14976 18760
rect 18880 18708 18932 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 13728 18640 13780 18692
rect 15016 18640 15068 18692
rect 16028 18640 16080 18692
rect 16304 18640 16356 18692
rect 18328 18640 18380 18692
rect 19248 18640 19300 18692
rect 8208 18572 8260 18624
rect 8576 18572 8628 18624
rect 10508 18572 10560 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13544 18572 13596 18624
rect 15660 18572 15712 18624
rect 17132 18572 17184 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 19708 18572 19760 18624
rect 21088 18640 21140 18692
rect 22100 18708 22152 18760
rect 22192 18708 22244 18760
rect 22192 18572 22244 18624
rect 22836 18708 22888 18760
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 22560 18640 22612 18692
rect 22836 18572 22888 18624
rect 23020 18572 23072 18624
rect 24124 18708 24176 18760
rect 25688 18640 25740 18692
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 2136 18368 2188 18420
rect 2872 18368 2924 18420
rect 4068 18368 4120 18420
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 5816 18411 5868 18420
rect 5816 18377 5825 18411
rect 5825 18377 5859 18411
rect 5859 18377 5868 18411
rect 5816 18368 5868 18377
rect 7012 18368 7064 18420
rect 7656 18411 7708 18420
rect 7656 18377 7665 18411
rect 7665 18377 7699 18411
rect 7699 18377 7708 18411
rect 7656 18368 7708 18377
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 2504 18232 2556 18284
rect 3332 18232 3384 18284
rect 3700 18232 3752 18284
rect 6736 18300 6788 18352
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 6920 18232 6972 18284
rect 9128 18300 9180 18352
rect 10784 18368 10836 18420
rect 12072 18368 12124 18420
rect 13820 18368 13872 18420
rect 14740 18368 14792 18420
rect 15660 18411 15712 18420
rect 15660 18377 15669 18411
rect 15669 18377 15703 18411
rect 15703 18377 15712 18411
rect 15660 18368 15712 18377
rect 10876 18300 10928 18352
rect 10968 18300 11020 18352
rect 11796 18300 11848 18352
rect 18512 18368 18564 18420
rect 20352 18368 20404 18420
rect 17408 18300 17460 18352
rect 17960 18300 18012 18352
rect 20536 18300 20588 18352
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 5540 18164 5592 18216
rect 8760 18164 8812 18216
rect 10508 18232 10560 18284
rect 16304 18232 16356 18284
rect 17132 18232 17184 18284
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18236 18232 18288 18284
rect 2780 18096 2832 18148
rect 2688 18028 2740 18080
rect 8392 18096 8444 18148
rect 9312 18164 9364 18216
rect 3240 18028 3292 18080
rect 6552 18028 6604 18080
rect 7840 18028 7892 18080
rect 9036 18028 9088 18080
rect 9772 18028 9824 18080
rect 10876 18028 10928 18080
rect 11612 18028 11664 18080
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12440 18164 12492 18216
rect 16212 18164 16264 18216
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 17500 18164 17552 18216
rect 12440 18028 12492 18080
rect 20444 18232 20496 18284
rect 18696 18207 18748 18216
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19524 18164 19576 18216
rect 19800 18207 19852 18216
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 20996 18300 21048 18352
rect 23112 18368 23164 18420
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 24124 18368 24176 18420
rect 24676 18368 24728 18420
rect 21456 18300 21508 18352
rect 24308 18300 24360 18352
rect 25872 18300 25924 18352
rect 21824 18232 21876 18284
rect 20720 18164 20772 18216
rect 20996 18207 21048 18216
rect 20996 18173 21005 18207
rect 21005 18173 21039 18207
rect 21039 18173 21048 18207
rect 20996 18164 21048 18173
rect 21272 18164 21324 18216
rect 24676 18164 24728 18216
rect 14740 18028 14792 18080
rect 17500 18028 17552 18080
rect 18236 18028 18288 18080
rect 20536 18096 20588 18148
rect 19248 18071 19300 18080
rect 19248 18037 19257 18071
rect 19257 18037 19291 18071
rect 19291 18037 19300 18071
rect 19248 18028 19300 18037
rect 20720 18028 20772 18080
rect 21824 18096 21876 18148
rect 22100 18096 22152 18148
rect 23388 18096 23440 18148
rect 22560 18028 22612 18080
rect 25504 18164 25556 18216
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 4988 17824 5040 17876
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 7012 17824 7064 17876
rect 7196 17824 7248 17876
rect 7840 17824 7892 17876
rect 8760 17824 8812 17876
rect 9312 17824 9364 17876
rect 11244 17824 11296 17876
rect 8300 17756 8352 17808
rect 11060 17756 11112 17808
rect 13360 17824 13412 17876
rect 13452 17824 13504 17876
rect 18880 17824 18932 17876
rect 19156 17824 19208 17876
rect 19892 17824 19944 17876
rect 20720 17824 20772 17876
rect 22192 17824 22244 17876
rect 22652 17824 22704 17876
rect 22836 17824 22888 17876
rect 17316 17756 17368 17808
rect 24860 17824 24912 17876
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 5264 17688 5316 17740
rect 6000 17688 6052 17740
rect 6368 17688 6420 17740
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 7840 17620 7892 17672
rect 9036 17688 9088 17740
rect 3332 17484 3384 17536
rect 3884 17527 3936 17536
rect 3884 17493 3893 17527
rect 3893 17493 3927 17527
rect 3927 17493 3936 17527
rect 3884 17484 3936 17493
rect 8484 17552 8536 17604
rect 4620 17484 4672 17536
rect 7564 17484 7616 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 11704 17688 11756 17740
rect 12624 17688 12676 17740
rect 13728 17688 13780 17740
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 15660 17688 15712 17740
rect 15844 17688 15896 17740
rect 16396 17688 16448 17740
rect 16764 17688 16816 17740
rect 16304 17620 16356 17672
rect 18604 17620 18656 17672
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 9496 17552 9548 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 11612 17552 11664 17604
rect 12716 17552 12768 17604
rect 13636 17552 13688 17604
rect 15200 17595 15252 17604
rect 15200 17561 15209 17595
rect 15209 17561 15243 17595
rect 15243 17561 15252 17595
rect 15200 17552 15252 17561
rect 11428 17484 11480 17536
rect 11980 17484 12032 17536
rect 12532 17484 12584 17536
rect 17408 17552 17460 17604
rect 16580 17484 16632 17536
rect 17684 17484 17736 17536
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 18788 17484 18840 17536
rect 19616 17484 19668 17536
rect 19892 17731 19944 17740
rect 19892 17697 19901 17731
rect 19901 17697 19935 17731
rect 19935 17697 19944 17731
rect 19892 17688 19944 17697
rect 20352 17688 20404 17740
rect 22560 17688 22612 17740
rect 23204 17688 23256 17740
rect 23940 17731 23992 17740
rect 23940 17697 23949 17731
rect 23949 17697 23983 17731
rect 23983 17697 23992 17731
rect 23940 17688 23992 17697
rect 24308 17688 24360 17740
rect 25780 17688 25832 17740
rect 23388 17620 23440 17672
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 24492 17620 24544 17672
rect 20720 17484 20772 17536
rect 21272 17552 21324 17604
rect 23572 17552 23624 17604
rect 24124 17484 24176 17536
rect 24216 17484 24268 17536
rect 24492 17484 24544 17536
rect 24584 17484 24636 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 6920 17280 6972 17332
rect 8392 17280 8444 17332
rect 16580 17280 16632 17332
rect 16856 17280 16908 17332
rect 23112 17280 23164 17332
rect 4620 17144 4672 17196
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 9128 17212 9180 17264
rect 9772 17212 9824 17264
rect 11612 17212 11664 17264
rect 11980 17255 12032 17264
rect 11980 17221 11989 17255
rect 11989 17221 12023 17255
rect 12023 17221 12032 17255
rect 11980 17212 12032 17221
rect 12716 17212 12768 17264
rect 13452 17212 13504 17264
rect 6920 17144 6972 17196
rect 7288 17144 7340 17196
rect 7564 17144 7616 17196
rect 4712 17076 4764 17128
rect 6552 17076 6604 17128
rect 8300 17144 8352 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9036 17144 9088 17196
rect 11704 17187 11756 17196
rect 7932 17076 7984 17128
rect 9864 17076 9916 17128
rect 10048 17076 10100 17128
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 7472 17008 7524 17060
rect 7564 17008 7616 17060
rect 8576 17051 8628 17060
rect 8576 17017 8585 17051
rect 8585 17017 8619 17051
rect 8619 17017 8628 17051
rect 8576 17008 8628 17017
rect 8852 16940 8904 16992
rect 9036 16940 9088 16992
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 12624 17076 12676 17128
rect 13820 17076 13872 17128
rect 11980 16940 12032 16992
rect 15108 17008 15160 17060
rect 17868 17212 17920 17264
rect 16948 17144 17000 17196
rect 18880 17212 18932 17264
rect 21548 17212 21600 17264
rect 22100 17212 22152 17264
rect 23664 17280 23716 17332
rect 24308 17323 24360 17332
rect 24308 17289 24317 17323
rect 24317 17289 24351 17323
rect 24351 17289 24360 17323
rect 24308 17280 24360 17289
rect 24124 17212 24176 17264
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 17684 17076 17736 17128
rect 19156 17076 19208 17128
rect 19340 17076 19392 17128
rect 20076 17119 20128 17128
rect 20076 17085 20085 17119
rect 20085 17085 20119 17119
rect 20119 17085 20128 17119
rect 20076 17076 20128 17085
rect 22284 17144 22336 17196
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 25136 17212 25188 17264
rect 21272 17076 21324 17128
rect 21824 17076 21876 17128
rect 16488 17008 16540 17060
rect 15016 16940 15068 16992
rect 16580 16940 16632 16992
rect 20628 16940 20680 16992
rect 21272 16940 21324 16992
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 22376 16940 22428 16992
rect 25504 17008 25556 17060
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 4620 16736 4672 16788
rect 4712 16736 4764 16788
rect 7932 16736 7984 16788
rect 8392 16779 8444 16788
rect 8392 16745 8401 16779
rect 8401 16745 8435 16779
rect 8435 16745 8444 16779
rect 8392 16736 8444 16745
rect 9404 16736 9456 16788
rect 6920 16711 6972 16720
rect 6920 16677 6929 16711
rect 6929 16677 6963 16711
rect 6963 16677 6972 16711
rect 6920 16668 6972 16677
rect 11060 16668 11112 16720
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 8668 16600 8720 16652
rect 10048 16600 10100 16652
rect 15016 16736 15068 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 21732 16736 21784 16788
rect 22284 16736 22336 16788
rect 19340 16668 19392 16720
rect 20720 16668 20772 16720
rect 21548 16668 21600 16720
rect 12256 16600 12308 16652
rect 14924 16600 14976 16652
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22652 16600 22704 16652
rect 8760 16532 8812 16584
rect 10968 16532 11020 16584
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11704 16532 11756 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 21272 16532 21324 16584
rect 25228 16532 25280 16584
rect 11796 16464 11848 16516
rect 12532 16464 12584 16516
rect 12716 16464 12768 16516
rect 15016 16464 15068 16516
rect 16304 16464 16356 16516
rect 21824 16464 21876 16516
rect 24124 16464 24176 16516
rect 4712 16439 4764 16448
rect 4712 16405 4721 16439
rect 4721 16405 4755 16439
rect 4755 16405 4764 16439
rect 4712 16396 4764 16405
rect 8852 16396 8904 16448
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 12348 16396 12400 16448
rect 14372 16396 14424 16448
rect 14924 16396 14976 16448
rect 18328 16396 18380 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 19156 16396 19208 16448
rect 21272 16396 21324 16448
rect 21456 16396 21508 16448
rect 23940 16396 23992 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 8300 16192 8352 16244
rect 4712 16124 4764 16176
rect 9680 16192 9732 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 10140 16192 10192 16244
rect 9496 16124 9548 16176
rect 12624 16124 12676 16176
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 14556 16192 14608 16244
rect 15016 16235 15068 16244
rect 15016 16201 15025 16235
rect 15025 16201 15059 16235
rect 15059 16201 15068 16235
rect 15016 16192 15068 16201
rect 16304 16192 16356 16244
rect 18512 16192 18564 16244
rect 19708 16192 19760 16244
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 9404 16056 9456 16108
rect 10048 16056 10100 16108
rect 8392 15988 8444 16040
rect 11520 16056 11572 16108
rect 13912 16056 13964 16108
rect 15568 16056 15620 16108
rect 15752 16056 15804 16108
rect 18972 16056 19024 16108
rect 19708 16099 19760 16108
rect 19708 16065 19717 16099
rect 19717 16065 19751 16099
rect 19751 16065 19760 16099
rect 19708 16056 19760 16065
rect 6092 15920 6144 15972
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 9128 15895 9180 15904
rect 9128 15861 9137 15895
rect 9137 15861 9171 15895
rect 9171 15861 9180 15895
rect 9128 15852 9180 15861
rect 9588 15920 9640 15972
rect 10784 15852 10836 15904
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12348 15988 12400 16040
rect 12440 15988 12492 16040
rect 13360 15988 13412 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 21088 16192 21140 16244
rect 21916 16192 21968 16244
rect 23848 16235 23900 16244
rect 23848 16201 23857 16235
rect 23857 16201 23891 16235
rect 23891 16201 23900 16235
rect 23848 16192 23900 16201
rect 25228 16235 25280 16244
rect 25228 16201 25237 16235
rect 25237 16201 25271 16235
rect 25271 16201 25280 16235
rect 25228 16192 25280 16201
rect 25780 16124 25832 16176
rect 20904 16056 20956 16108
rect 13544 15852 13596 15904
rect 15016 15852 15068 15904
rect 17592 15920 17644 15972
rect 19892 16031 19944 16040
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 17408 15852 17460 15904
rect 20812 15852 20864 15904
rect 21088 15920 21140 15972
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 23756 16099 23808 16108
rect 23756 16065 23765 16099
rect 23765 16065 23799 16099
rect 23799 16065 23808 16099
rect 23756 16056 23808 16065
rect 24032 16056 24084 16108
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 22192 15988 22244 16040
rect 23940 16031 23992 16040
rect 23940 15997 23949 16031
rect 23949 15997 23983 16031
rect 23983 15997 23992 16031
rect 23940 15988 23992 15997
rect 22192 15852 22244 15904
rect 22652 15852 22704 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9956 15648 10008 15700
rect 12164 15648 12216 15700
rect 11796 15580 11848 15632
rect 12532 15648 12584 15700
rect 14096 15648 14148 15700
rect 15200 15648 15252 15700
rect 16672 15691 16724 15700
rect 16672 15657 16681 15691
rect 16681 15657 16715 15691
rect 16715 15657 16724 15691
rect 16672 15648 16724 15657
rect 17960 15648 18012 15700
rect 19800 15648 19852 15700
rect 22192 15648 22244 15700
rect 22744 15648 22796 15700
rect 22928 15648 22980 15700
rect 24124 15691 24176 15700
rect 24124 15657 24133 15691
rect 24133 15657 24167 15691
rect 24167 15657 24176 15691
rect 24124 15648 24176 15657
rect 24584 15648 24636 15700
rect 12348 15580 12400 15632
rect 13544 15580 13596 15632
rect 18328 15580 18380 15632
rect 21640 15580 21692 15632
rect 8944 15512 8996 15564
rect 10416 15512 10468 15564
rect 13268 15512 13320 15564
rect 14188 15512 14240 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 16856 15512 16908 15564
rect 18880 15512 18932 15564
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 24032 15580 24084 15632
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10232 15444 10284 15496
rect 13820 15444 13872 15496
rect 16304 15444 16356 15496
rect 18328 15444 18380 15496
rect 18604 15444 18656 15496
rect 20904 15444 20956 15496
rect 22836 15512 22888 15564
rect 25596 15512 25648 15564
rect 26240 15512 26292 15564
rect 10692 15376 10744 15428
rect 7748 15308 7800 15360
rect 10968 15308 11020 15360
rect 11152 15308 11204 15360
rect 12624 15376 12676 15428
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 12348 15308 12400 15360
rect 14648 15376 14700 15428
rect 16580 15376 16632 15428
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 19248 15308 19300 15360
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 20812 15308 20864 15360
rect 20904 15308 20956 15360
rect 22376 15376 22428 15428
rect 24952 15376 25004 15428
rect 26608 15308 26660 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10232 15104 10284 15156
rect 13820 15104 13872 15156
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12624 15036 12676 15088
rect 14648 15036 14700 15088
rect 16764 15036 16816 15088
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 10324 14875 10376 14884
rect 10324 14841 10333 14875
rect 10333 14841 10367 14875
rect 10367 14841 10376 14875
rect 10324 14832 10376 14841
rect 10692 14900 10744 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 12532 14900 12584 14952
rect 16028 14968 16080 15020
rect 17408 15036 17460 15088
rect 18972 15147 19024 15156
rect 18972 15113 18981 15147
rect 18981 15113 19015 15147
rect 19015 15113 19024 15147
rect 18972 15104 19024 15113
rect 21272 15104 21324 15156
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 21456 15036 21508 15088
rect 21548 15036 21600 15088
rect 22192 15036 22244 15088
rect 23020 15036 23072 15088
rect 23940 15104 23992 15156
rect 24400 15104 24452 15156
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 11152 14832 11204 14884
rect 13544 14832 13596 14884
rect 18236 14968 18288 15020
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 11060 14764 11112 14816
rect 12072 14764 12124 14816
rect 16396 14764 16448 14816
rect 16488 14764 16540 14816
rect 17868 14900 17920 14952
rect 19340 14943 19392 14952
rect 17132 14764 17184 14816
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 20720 14832 20772 14884
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 19800 14764 19852 14816
rect 21732 14900 21784 14952
rect 22284 14968 22336 15020
rect 24216 14968 24268 15020
rect 25136 15011 25188 15020
rect 25136 14977 25145 15011
rect 25145 14977 25179 15011
rect 25179 14977 25188 15011
rect 25136 14968 25188 14977
rect 23204 14900 23256 14952
rect 21272 14832 21324 14884
rect 22100 14832 22152 14884
rect 25320 14875 25372 14884
rect 25320 14841 25329 14875
rect 25329 14841 25363 14875
rect 25363 14841 25372 14875
rect 25320 14832 25372 14841
rect 21456 14764 21508 14816
rect 23296 14764 23348 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10508 14560 10560 14612
rect 12532 14560 12584 14612
rect 13820 14560 13872 14612
rect 24768 14560 24820 14612
rect 25136 14560 25188 14612
rect 15936 14492 15988 14544
rect 16212 14492 16264 14544
rect 18696 14492 18748 14544
rect 20076 14492 20128 14544
rect 20536 14492 20588 14544
rect 21456 14492 21508 14544
rect 21548 14492 21600 14544
rect 12256 14424 12308 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 18604 14424 18656 14476
rect 21916 14424 21968 14476
rect 22284 14424 22336 14476
rect 23848 14492 23900 14544
rect 24216 14492 24268 14544
rect 23480 14424 23532 14476
rect 24584 14424 24636 14476
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 14096 14356 14148 14408
rect 15936 14356 15988 14408
rect 16304 14356 16356 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 19432 14356 19484 14408
rect 21364 14356 21416 14408
rect 24124 14356 24176 14408
rect 12624 14288 12676 14340
rect 13820 14220 13872 14272
rect 14096 14220 14148 14272
rect 14372 14220 14424 14272
rect 18236 14288 18288 14340
rect 16764 14220 16816 14272
rect 17132 14220 17184 14272
rect 18604 14220 18656 14272
rect 23388 14288 23440 14340
rect 25412 14288 25464 14340
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 20904 14220 20956 14272
rect 22008 14220 22060 14272
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 11336 14016 11388 14068
rect 11888 14016 11940 14068
rect 12808 14016 12860 14068
rect 14004 14016 14056 14068
rect 14648 14016 14700 14068
rect 15844 14016 15896 14068
rect 17132 14016 17184 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 13636 13880 13688 13932
rect 14280 13948 14332 14000
rect 15936 13948 15988 14000
rect 18512 13948 18564 14000
rect 19248 14016 19300 14068
rect 20536 14016 20588 14068
rect 20628 14016 20680 14068
rect 22008 14016 22060 14068
rect 22652 14016 22704 14068
rect 19800 13948 19852 14000
rect 16396 13880 16448 13932
rect 14464 13812 14516 13864
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 20904 13948 20956 14000
rect 21732 13948 21784 14000
rect 20720 13880 20772 13932
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 19984 13812 20036 13864
rect 22100 13923 22152 13932
rect 22100 13889 22109 13923
rect 22109 13889 22143 13923
rect 22143 13889 22152 13923
rect 23388 13948 23440 14000
rect 23848 13948 23900 14000
rect 22100 13880 22152 13889
rect 22284 13880 22336 13932
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25872 13880 25924 13932
rect 15568 13744 15620 13796
rect 18512 13744 18564 13796
rect 19524 13744 19576 13796
rect 21456 13812 21508 13864
rect 24400 13812 24452 13864
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 25228 13812 25280 13864
rect 14004 13719 14056 13728
rect 14004 13685 14034 13719
rect 14034 13685 14056 13719
rect 14004 13676 14056 13685
rect 15936 13676 15988 13728
rect 16580 13676 16632 13728
rect 16764 13676 16816 13728
rect 17316 13676 17368 13728
rect 19432 13676 19484 13728
rect 20536 13676 20588 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 22744 13676 22796 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 14004 13472 14056 13524
rect 13360 13404 13412 13456
rect 19708 13472 19760 13524
rect 19800 13472 19852 13524
rect 20996 13472 21048 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 23480 13472 23532 13524
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 11520 13200 11572 13252
rect 10048 13132 10100 13184
rect 10692 13132 10744 13184
rect 13452 13200 13504 13252
rect 14188 13200 14240 13252
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 18696 13336 18748 13388
rect 21916 13379 21968 13388
rect 17868 13268 17920 13320
rect 19524 13268 19576 13320
rect 16764 13200 16816 13252
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 23848 13404 23900 13456
rect 24768 13404 24820 13456
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 24860 13336 24912 13388
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 15936 13132 15988 13184
rect 16304 13132 16356 13184
rect 17592 13132 17644 13184
rect 18880 13132 18932 13184
rect 19892 13200 19944 13252
rect 20996 13200 21048 13252
rect 22192 13243 22244 13252
rect 22192 13209 22201 13243
rect 22201 13209 22235 13243
rect 22235 13209 22244 13243
rect 22192 13200 22244 13209
rect 25596 13200 25648 13252
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 13452 12928 13504 12980
rect 13820 12928 13872 12980
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 17316 12928 17368 12980
rect 15568 12860 15620 12912
rect 19064 12928 19116 12980
rect 19616 12928 19668 12980
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 22192 12928 22244 12980
rect 25136 12928 25188 12980
rect 22560 12860 22612 12912
rect 23848 12860 23900 12912
rect 24032 12860 24084 12912
rect 24768 12860 24820 12912
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18236 12792 18288 12844
rect 18420 12792 18472 12844
rect 21640 12792 21692 12844
rect 21916 12792 21968 12844
rect 24676 12792 24728 12844
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 16672 12724 16724 12776
rect 17500 12724 17552 12776
rect 18328 12724 18380 12776
rect 18788 12724 18840 12776
rect 19064 12724 19116 12776
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 18604 12656 18656 12665
rect 20444 12656 20496 12708
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 15936 12588 15988 12640
rect 16580 12588 16632 12640
rect 17868 12588 17920 12640
rect 18328 12588 18380 12640
rect 18512 12588 18564 12640
rect 19248 12588 19300 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20536 12588 20588 12640
rect 20904 12588 20956 12640
rect 22100 12588 22152 12640
rect 22652 12588 22704 12640
rect 24032 12588 24084 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 14096 12384 14148 12436
rect 15568 12384 15620 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 18236 12384 18288 12436
rect 18788 12384 18840 12436
rect 4068 12248 4120 12300
rect 5724 12044 5776 12096
rect 14372 12044 14424 12096
rect 16764 12248 16816 12300
rect 17408 12248 17460 12300
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 18236 12180 18288 12232
rect 20812 12180 20864 12232
rect 16304 12112 16356 12164
rect 18696 12155 18748 12164
rect 18696 12121 18703 12155
rect 18703 12121 18748 12155
rect 18696 12112 18748 12121
rect 19248 12112 19300 12164
rect 22376 12384 22428 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 21364 12248 21416 12300
rect 21916 12248 21968 12300
rect 24584 12248 24636 12300
rect 22100 12180 22152 12232
rect 24216 12180 24268 12232
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 19340 12044 19392 12096
rect 20352 12044 20404 12096
rect 20444 12044 20496 12096
rect 21272 12044 21324 12096
rect 23940 12044 23992 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 13820 11840 13872 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 14832 11840 14884 11892
rect 13360 11772 13412 11824
rect 14372 11772 14424 11824
rect 14740 11772 14792 11824
rect 17316 11840 17368 11892
rect 19340 11840 19392 11892
rect 19616 11840 19668 11892
rect 15936 11704 15988 11756
rect 18788 11772 18840 11824
rect 16580 11704 16632 11756
rect 19708 11772 19760 11824
rect 20812 11704 20864 11756
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 18604 11636 18656 11688
rect 20444 11636 20496 11688
rect 21180 11883 21232 11892
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 21732 11840 21784 11892
rect 22100 11840 22152 11892
rect 23388 11840 23440 11892
rect 24860 11772 24912 11824
rect 23572 11704 23624 11756
rect 22468 11636 22520 11688
rect 23848 11636 23900 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 25136 11636 25188 11688
rect 26332 11636 26384 11688
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 15568 11500 15620 11552
rect 21272 11568 21324 11620
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 16028 11296 16080 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 16948 11296 17000 11348
rect 17040 11296 17092 11348
rect 18604 11296 18656 11348
rect 14740 11271 14792 11280
rect 14740 11237 14749 11271
rect 14749 11237 14783 11271
rect 14783 11237 14792 11271
rect 14740 11228 14792 11237
rect 15936 11228 15988 11280
rect 18696 11228 18748 11280
rect 24492 11296 24544 11348
rect 26056 11296 26108 11348
rect 18420 11160 18472 11212
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 16396 11092 16448 11144
rect 21456 11160 21508 11212
rect 21640 11203 21692 11212
rect 21640 11169 21649 11203
rect 21649 11169 21683 11203
rect 21683 11169 21692 11203
rect 21640 11160 21692 11169
rect 22192 11203 22244 11212
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 17132 11024 17184 11076
rect 18328 11024 18380 11076
rect 18788 11024 18840 11076
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 19892 11092 19944 11144
rect 20076 11092 20128 11144
rect 23480 11228 23532 11280
rect 25872 11228 25924 11280
rect 24860 11160 24912 11212
rect 22744 11092 22796 11144
rect 18696 10999 18748 11008
rect 18696 10965 18705 10999
rect 18705 10965 18739 10999
rect 18739 10965 18748 10999
rect 18696 10956 18748 10965
rect 20536 11024 20588 11076
rect 24308 11024 24360 11076
rect 20812 10956 20864 11008
rect 21456 10956 21508 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 15660 10752 15712 10804
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 18512 10616 18564 10668
rect 19708 10752 19760 10804
rect 20076 10752 20128 10804
rect 21548 10752 21600 10804
rect 20996 10684 21048 10736
rect 22560 10752 22612 10804
rect 24860 10684 24912 10736
rect 20076 10616 20128 10668
rect 20352 10616 20404 10668
rect 20720 10616 20772 10668
rect 22008 10616 22060 10668
rect 20168 10548 20220 10600
rect 21640 10548 21692 10600
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 17776 10480 17828 10532
rect 23940 10480 23992 10532
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 19708 10412 19760 10464
rect 20352 10412 20404 10464
rect 20812 10412 20864 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 19708 10208 19760 10260
rect 16672 10140 16724 10192
rect 21640 10208 21692 10260
rect 21824 10208 21876 10260
rect 20720 10183 20772 10192
rect 20720 10149 20729 10183
rect 20729 10149 20763 10183
rect 20763 10149 20772 10183
rect 20720 10140 20772 10149
rect 22744 10140 22796 10192
rect 21272 10072 21324 10124
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 19432 10004 19484 10056
rect 19708 10004 19760 10056
rect 20996 10004 21048 10056
rect 24216 10072 24268 10124
rect 24124 10004 24176 10056
rect 25780 10004 25832 10056
rect 19524 9868 19576 9920
rect 21180 9936 21232 9988
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 19708 9664 19760 9716
rect 22100 9664 22152 9716
rect 19432 9596 19484 9648
rect 8484 9528 8536 9580
rect 18880 9571 18932 9580
rect 18880 9537 18889 9571
rect 18889 9537 18923 9571
rect 18923 9537 18932 9571
rect 18880 9528 18932 9537
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 17224 9460 17276 9512
rect 21456 9571 21508 9580
rect 21456 9537 21465 9571
rect 21465 9537 21499 9571
rect 21499 9537 21508 9571
rect 21456 9528 21508 9537
rect 21732 9528 21784 9580
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 18604 9392 18656 9444
rect 19432 9392 19484 9444
rect 22836 9392 22888 9444
rect 15936 9324 15988 9376
rect 20996 9324 21048 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 14924 9120 14976 9172
rect 19524 9120 19576 9172
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 22560 9052 22612 9104
rect 24124 9120 24176 9172
rect 26240 9120 26292 9172
rect 26424 9052 26476 9104
rect 18880 8916 18932 8968
rect 23664 8984 23716 9036
rect 24860 8984 24912 9036
rect 9312 8848 9364 8900
rect 12532 8848 12584 8900
rect 19892 8916 19944 8968
rect 21088 8916 21140 8968
rect 21640 8916 21692 8968
rect 22100 8848 22152 8900
rect 25044 8848 25096 8900
rect 23848 8780 23900 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 19616 8576 19668 8628
rect 20904 8576 20956 8628
rect 19156 8508 19208 8560
rect 15292 8440 15344 8492
rect 20996 8508 21048 8560
rect 21916 8440 21968 8492
rect 24860 8508 24912 8560
rect 24952 8440 25004 8492
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 16212 8304 16264 8356
rect 21732 8304 21784 8356
rect 21548 8236 21600 8288
rect 24032 8236 24084 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 22100 8032 22152 8084
rect 23572 7964 23624 8016
rect 19800 7896 19852 7948
rect 25596 7964 25648 8016
rect 18696 7828 18748 7880
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 24952 7896 25004 7948
rect 24492 7828 24544 7880
rect 25688 7760 25740 7812
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 23480 7692 23532 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 20720 7420 20772 7472
rect 20260 7352 20312 7404
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 24860 7420 24912 7472
rect 25320 7352 25372 7404
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 23296 7148 23348 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 19340 6808 19392 6860
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 23756 6808 23808 6860
rect 24860 6808 24912 6860
rect 22836 6740 22888 6792
rect 25044 6672 25096 6724
rect 21640 6604 21692 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 21456 6400 21508 6452
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 24952 6400 25004 6452
rect 24860 6332 24912 6384
rect 25504 6264 25556 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 15200 5856 15252 5908
rect 24584 5788 24636 5840
rect 21732 5720 21784 5772
rect 21824 5652 21876 5704
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 23480 5652 23532 5704
rect 24952 5584 25004 5636
rect 23480 5516 23532 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 24860 5244 24912 5296
rect 23388 5176 23440 5228
rect 23848 5176 23900 5228
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 19064 4768 19116 4820
rect 22284 4564 22336 4616
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23296 4564 23348 4616
rect 24952 4496 25004 4548
rect 22284 4428 22336 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 19984 4088 20036 4140
rect 18972 4020 19024 4072
rect 20168 4020 20220 4072
rect 22100 4020 22152 4072
rect 25044 4088 25096 4140
rect 26608 4088 26660 4140
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 7472 3476 7524 3528
rect 20536 3476 20588 3528
rect 23480 3476 23532 3528
rect 24584 3476 24636 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24952 3408 25004 3460
rect 7196 3340 7248 3392
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 19248 3068 19300 3120
rect 6736 3000 6788 3052
rect 19800 3000 19852 3052
rect 24860 3068 24912 3120
rect 25136 3111 25188 3120
rect 25136 3077 25145 3111
rect 25145 3077 25179 3111
rect 25179 3077 25188 3111
rect 25136 3068 25188 3077
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 25412 3000 25464 3052
rect 19524 2932 19576 2984
rect 25044 2932 25096 2984
rect 6736 2796 6788 2848
rect 19800 2796 19852 2848
rect 25228 2796 25280 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 8668 2592 8720 2644
rect 19800 2635 19852 2644
rect 19800 2601 19809 2635
rect 19809 2601 19843 2635
rect 19843 2601 19852 2635
rect 19800 2592 19852 2601
rect 19524 2456 19576 2508
rect 22744 2456 22796 2508
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 22652 2388 22704 2440
rect 24584 2388 24636 2440
rect 23388 2320 23440 2372
rect 24952 2320 25004 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 2042 26200 2098 27000
rect 2410 26330 2466 27000
rect 2778 26466 2834 27000
rect 2778 26450 3096 26466
rect 2778 26444 3108 26450
rect 2778 26438 3056 26444
rect 2410 26302 2728 26330
rect 2410 26200 2466 26302
rect 2504 26240 2556 26246
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 1412 21622 1440 25871
rect 1490 24848 1546 24857
rect 1490 24783 1546 24792
rect 1504 22778 1532 24783
rect 1582 24168 1638 24177
rect 1582 24103 1584 24112
rect 1636 24103 1638 24112
rect 1584 24074 1636 24080
rect 1688 23882 1716 26200
rect 1950 24712 2006 24721
rect 1950 24647 2006 24656
rect 1688 23854 1900 23882
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 1688 22681 1716 23666
rect 1674 22672 1730 22681
rect 1674 22607 1730 22616
rect 1688 22098 1716 22607
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1400 21616 1452 21622
rect 1400 21558 1452 21564
rect 1872 19310 1900 23854
rect 1964 23254 1992 24647
rect 1952 23248 2004 23254
rect 1952 23190 2004 23196
rect 2056 19922 2084 26200
rect 2504 26182 2556 26188
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2320 24676 2372 24682
rect 2320 24618 2372 24624
rect 2332 24070 2360 24618
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 2332 23866 2360 24006
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22234 2268 22374
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2148 18766 2176 21830
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2240 19417 2268 19790
rect 2226 19408 2282 19417
rect 2226 19343 2282 19352
rect 2424 18970 2452 24754
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18426 2176 18702
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 2516 18290 2544 26182
rect 2700 23474 2728 26302
rect 2778 26200 2834 26438
rect 3056 26386 3108 26392
rect 3146 26330 3202 27000
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 2884 26302 3202 26330
rect 2700 23446 2820 23474
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2700 18086 2728 21966
rect 2792 21078 2820 23446
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 3344 20398 3372 26386
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3422 23760 3478 23769
rect 3422 23695 3478 23704
rect 3436 20534 3464 23695
rect 3528 21486 3556 26200
rect 3974 25392 4030 25401
rect 3974 25327 4030 25336
rect 3988 24410 4016 25327
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 3620 23322 3648 23666
rect 3608 23316 3660 23322
rect 3608 23258 3660 23264
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 2792 18154 2820 19751
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2884 18426 2912 19246
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 3252 18086 3280 18566
rect 3344 18290 3372 19110
rect 3620 18970 3648 22510
rect 3896 19514 3924 24142
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3988 23225 4016 23258
rect 3974 23216 4030 23225
rect 3974 23151 4030 23160
rect 4080 22094 4108 26302
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4986 26330 5042 27000
rect 4986 26302 5120 26330
rect 4986 26200 5042 26302
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 22506 4200 24142
rect 4264 22710 4292 26200
rect 4632 23186 4660 26200
rect 4986 25800 5042 25809
rect 4986 25735 5042 25744
rect 4804 25016 4856 25022
rect 4804 24958 4856 24964
rect 4816 24206 4844 24958
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4618 23080 4674 23089
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4080 22066 4200 22094
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 20806 4016 21966
rect 4172 21010 4200 22066
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3712 18290 3740 18906
rect 4264 18698 4292 20266
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3330 17912 3386 17921
rect 3330 17847 3386 17856
rect 2226 17776 2282 17785
rect 2226 17711 2228 17720
rect 2280 17711 2282 17720
rect 2228 17682 2280 17688
rect 3344 17542 3372 17847
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3896 17105 3924 17478
rect 3882 17096 3938 17105
rect 3882 17031 3938 17040
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 4080 12306 4108 18362
rect 4356 13977 4384 23054
rect 4618 23015 4674 23024
rect 4528 22636 4580 22642
rect 4528 22578 4580 22584
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4448 15473 4476 21966
rect 4540 18426 4568 22578
rect 4632 19514 4660 23015
rect 4896 20528 4948 20534
rect 4894 20496 4896 20505
rect 4948 20496 4950 20505
rect 4894 20431 4950 20440
rect 4908 19854 4936 20431
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4802 19680 4858 19689
rect 4802 19615 4858 19624
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4710 19136 4766 19145
rect 4710 19071 4766 19080
rect 4724 18766 4752 19071
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4710 17776 4766 17785
rect 4710 17711 4766 17720
rect 4724 17678 4752 17711
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17202 4660 17478
rect 4816 17202 4844 19615
rect 5000 17882 5028 25735
rect 5092 21486 5120 26302
rect 5170 26208 5226 26217
rect 5354 26200 5410 27000
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26330 6882 27000
rect 6564 26302 6882 26330
rect 5170 26143 5226 26152
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5184 21162 5212 26143
rect 5368 23798 5396 26200
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5262 22672 5318 22681
rect 5262 22607 5318 22616
rect 5092 21134 5212 21162
rect 5092 18766 5120 21134
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5184 19922 5212 21014
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5276 17746 5304 22607
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5368 20233 5396 20470
rect 5354 20224 5410 20233
rect 5354 20159 5410 20168
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 18290 5396 19654
rect 5460 19378 5488 23462
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5552 22545 5580 23054
rect 5736 22710 5764 26200
rect 5816 24744 5868 24750
rect 5816 24686 5868 24692
rect 5828 23798 5856 24686
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5920 23594 5948 24550
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 5816 23044 5868 23050
rect 5816 22986 5868 22992
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5538 22536 5594 22545
rect 5538 22471 5594 22480
rect 5644 21049 5672 22578
rect 5828 22438 5856 22986
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 21146 5856 22374
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5630 21040 5686 21049
rect 5630 20975 5686 20984
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20369 5580 20402
rect 5538 20360 5594 20369
rect 5538 20295 5594 20304
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5538 19000 5594 19009
rect 5538 18935 5540 18944
rect 5592 18935 5594 18944
rect 5540 18906 5592 18912
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5540 18216 5592 18222
rect 5538 18184 5540 18193
rect 5592 18184 5594 18193
rect 5538 18119 5594 18128
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4632 16794 4660 17138
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16794 4752 17070
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4724 16182 4752 16390
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4434 15464 4490 15473
rect 4434 15399 4490 15408
rect 4342 13968 4398 13977
rect 4342 13903 4398 13912
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 5736 12102 5764 18634
rect 5828 18426 5856 20878
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5920 18970 5948 19382
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 6012 17746 6040 23598
rect 6104 22098 6132 26200
rect 6472 24274 6500 26200
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6182 23488 6238 23497
rect 6182 23423 6238 23432
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 6104 15978 6132 21490
rect 6196 19922 6224 23423
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6288 19514 6316 23054
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6196 15065 6224 18702
rect 6380 17746 6408 24006
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 17882 6500 21966
rect 6564 21010 6592 26302
rect 6826 26200 6882 26302
rect 7194 26200 7250 27000
rect 7562 26330 7618 27000
rect 7930 26330 7986 27000
rect 7300 26302 7618 26330
rect 6642 26072 6698 26081
rect 6642 26007 6698 26016
rect 6656 21434 6684 26007
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6748 24206 6776 24346
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6840 23769 6868 23802
rect 6826 23760 6882 23769
rect 6736 23724 6788 23730
rect 6826 23695 6882 23704
rect 6920 23724 6972 23730
rect 6736 23666 6788 23672
rect 6920 23666 6972 23672
rect 6748 23322 6776 23666
rect 6932 23633 6960 23666
rect 6918 23624 6974 23633
rect 6918 23559 6974 23568
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6748 21690 6776 22578
rect 6932 22094 6960 22714
rect 6840 22066 6960 22094
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6656 21406 6776 21434
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6552 19304 6604 19310
rect 6550 19272 6552 19281
rect 6604 19272 6606 19281
rect 6550 19207 6606 19216
rect 6564 18834 6592 19207
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6564 17134 6592 18022
rect 6656 17678 6684 21286
rect 6748 19310 6776 21406
rect 6840 20602 6868 22066
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6932 20346 6960 21626
rect 7024 21457 7052 23190
rect 7116 22778 7144 24618
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7208 21468 7236 26200
rect 7300 24750 7328 26302
rect 7562 26200 7618 26302
rect 7668 26302 7986 26330
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7300 21690 7328 24142
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7380 22024 7432 22030
rect 7378 21992 7380 22001
rect 7432 21992 7434 22001
rect 7378 21927 7434 21936
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7010 21448 7066 21457
rect 7208 21440 7288 21468
rect 7288 21422 7340 21428
rect 7010 21383 7066 21392
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6840 20318 6960 20346
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6748 18358 6776 19246
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6840 18170 6868 20318
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19394 6960 20198
rect 7024 20058 7052 20402
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6932 19366 7052 19394
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6932 18290 6960 19178
rect 7024 18426 7052 19366
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6840 18142 6960 18170
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6932 17338 6960 18142
rect 7116 17898 7144 20878
rect 7300 20602 7328 20878
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7208 18834 7236 20198
rect 7286 19952 7342 19961
rect 7286 19887 7342 19896
rect 7300 19514 7328 19887
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7116 17882 7236 17898
rect 7012 17876 7064 17882
rect 7116 17876 7248 17882
rect 7116 17870 7196 17876
rect 7012 17818 7064 17824
rect 7196 17818 7248 17824
rect 7024 17649 7052 17818
rect 7010 17640 7066 17649
rect 7010 17575 7066 17584
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6182 15056 6238 15065
rect 6182 14991 6238 15000
rect 6564 14385 6592 16934
rect 6932 16726 6960 17138
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 7300 16658 7328 17138
rect 7392 16946 7420 21490
rect 7484 19922 7512 24006
rect 7668 23186 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26200 8722 27000
rect 9034 26330 9090 27000
rect 8772 26302 9090 26330
rect 7748 24880 7800 24886
rect 7748 24822 7800 24828
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7484 17066 7512 19654
rect 7576 18834 7604 22986
rect 7760 22094 7788 24822
rect 7838 24304 7894 24313
rect 7838 24239 7894 24248
rect 7668 22066 7788 22094
rect 7668 20992 7696 22066
rect 7668 20964 7788 20992
rect 7654 20904 7710 20913
rect 7654 20839 7656 20848
rect 7708 20839 7710 20848
rect 7656 20810 7708 20816
rect 7654 20088 7710 20097
rect 7654 20023 7710 20032
rect 7668 19990 7696 20023
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7668 18714 7696 19654
rect 7760 19378 7788 20964
rect 7852 20233 7880 24239
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 8036 23662 8064 23802
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22166 8340 26200
rect 8680 24138 8708 26200
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 8300 22160 8352 22166
rect 8206 22128 8262 22137
rect 8300 22102 8352 22108
rect 8206 22063 8262 22072
rect 8220 21894 8248 22063
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 7932 21412 7984 21418
rect 7932 21354 7984 21360
rect 7944 20942 7972 21354
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7838 20224 7894 20233
rect 7838 20159 7894 20168
rect 7944 19990 7972 20334
rect 8022 20224 8078 20233
rect 8022 20159 8078 20168
rect 7932 19984 7984 19990
rect 7932 19926 7984 19932
rect 7840 19848 7892 19854
rect 8036 19825 8064 20159
rect 8312 19938 8340 21422
rect 8220 19910 8340 19938
rect 7840 19790 7892 19796
rect 8022 19816 8078 19825
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7852 18834 7880 19790
rect 8022 19751 8078 19760
rect 8220 19718 8248 19910
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8404 19514 8432 22646
rect 8574 22400 8630 22409
rect 8574 22335 8630 22344
rect 8482 21720 8538 21729
rect 8482 21655 8538 21664
rect 8496 21622 8524 21655
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8588 21486 8616 22335
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7576 18686 7696 18714
rect 7576 17542 7604 18686
rect 7944 18612 7972 19314
rect 8206 18728 8262 18737
rect 8206 18663 8262 18672
rect 8220 18630 8248 18663
rect 7760 18584 7972 18612
rect 8208 18624 8260 18630
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7668 18329 7696 18362
rect 7654 18320 7710 18329
rect 7654 18255 7710 18264
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7562 17232 7618 17241
rect 7562 17167 7564 17176
rect 7616 17167 7618 17176
rect 7564 17138 7616 17144
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16946 7604 17002
rect 7392 16918 7604 16946
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7760 15366 7788 18584
rect 8208 18566 8260 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18426 8340 19382
rect 8390 18864 8446 18873
rect 8390 18799 8446 18808
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 18086 7880 18226
rect 8404 18154 8432 18799
rect 8496 18290 8524 21014
rect 8588 20466 8616 21286
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18970 8616 19110
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7852 17678 7880 17818
rect 8300 17808 8352 17814
rect 8298 17776 8300 17785
rect 8352 17776 8354 17785
rect 8298 17711 8354 17720
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7944 16794 7972 17070
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16250 8340 17138
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8404 16046 8432 16730
rect 8496 16561 8524 17546
rect 8588 17066 8616 18566
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8680 16658 8708 23122
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9692 26302 9826 26330
rect 9128 25084 9180 25090
rect 9128 25026 9180 25032
rect 8942 24984 8998 24993
rect 8942 24919 8998 24928
rect 8850 22808 8906 22817
rect 8850 22743 8906 22752
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8864 22386 8892 22743
rect 8772 22358 8892 22386
rect 8772 18222 8800 22358
rect 8956 22250 8984 24919
rect 9140 24410 9168 25026
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9324 23866 9352 24142
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9220 23520 9272 23526
rect 9220 23462 9272 23468
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 8864 22222 8984 22250
rect 8864 20806 8892 22222
rect 9048 22098 9076 22510
rect 9036 22092 9088 22098
rect 9036 22034 9088 22040
rect 9048 21554 9076 22034
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 9048 20466 9076 21490
rect 9140 21146 9168 23258
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9232 21010 9260 23462
rect 9416 23254 9444 26200
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26200 11298 27000
rect 11610 26200 11666 27000
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26330 12770 27000
rect 13082 26330 13138 27000
rect 12636 26302 12770 26330
rect 12636 26246 12664 26302
rect 12624 26240 12676 26246
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9600 23118 9628 24074
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9770 23896 9826 23905
rect 9770 23831 9826 23840
rect 9784 23730 9812 23831
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9508 22030 9536 22170
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9312 21888 9364 21894
rect 9310 21856 9312 21865
rect 9364 21856 9366 21865
rect 9310 21791 9366 21800
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8850 19544 8906 19553
rect 8850 19479 8906 19488
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 17882 8800 18158
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8758 17368 8814 17377
rect 8758 17303 8814 17312
rect 8772 17202 8800 17303
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8864 16998 8892 19479
rect 9048 19378 9076 20402
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8760 16584 8812 16590
rect 8482 16552 8538 16561
rect 8760 16526 8812 16532
rect 8482 16487 8538 16496
rect 8666 16144 8722 16153
rect 8666 16079 8668 16088
rect 8720 16079 8722 16088
rect 8668 16050 8720 16056
rect 8392 16040 8444 16046
rect 8772 16017 8800 16526
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8392 15982 8444 15988
rect 8758 16008 8814 16017
rect 8758 15943 8814 15952
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 6550 14376 6606 14385
rect 6550 14311 6606 14320
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8496 9586 8524 15846
rect 8772 15706 8800 15943
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8864 14521 8892 16390
rect 8956 15570 8984 19314
rect 9048 18086 9076 19314
rect 9140 18766 9168 19654
rect 9416 19258 9444 21898
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9784 20641 9812 20878
rect 9770 20632 9826 20641
rect 9770 20567 9826 20576
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9232 19230 9444 19258
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9232 18442 9260 19230
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9140 18414 9260 18442
rect 9140 18358 9168 18414
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9324 18222 9352 18634
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9048 17746 9076 18022
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9048 17202 9076 17682
rect 9324 17678 9352 17818
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17270 9168 17478
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9048 16998 9076 17138
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9416 16794 9444 19110
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9508 17610 9536 18770
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9416 16114 9444 16730
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16182 9536 16390
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9600 15978 9628 20470
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9692 16250 9720 19450
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17270 9812 18022
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9876 17134 9904 24006
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9770 16416 9826 16425
rect 9770 16351 9826 16360
rect 9784 16250 9812 16351
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9128 15904 9180 15910
rect 9126 15872 9128 15881
rect 9180 15872 9182 15881
rect 9126 15807 9182 15816
rect 9968 15706 9996 24142
rect 10152 23798 10180 26200
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 10060 23497 10088 23598
rect 10046 23488 10102 23497
rect 10046 23423 10102 23432
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22438 10088 22986
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10060 20602 10088 20946
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10060 17134 10088 17546
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10046 16688 10102 16697
rect 10046 16623 10048 16632
rect 10100 16623 10102 16632
rect 10048 16594 10100 16600
rect 10060 16114 10088 16594
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16250 10180 16390
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9402 15600 9458 15609
rect 8944 15564 8996 15570
rect 9402 15535 9458 15544
rect 8944 15506 8996 15512
rect 9416 15502 9444 15535
rect 10244 15502 10272 24890
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10336 21162 10364 24550
rect 10428 21962 10456 24686
rect 10520 23186 10548 26200
rect 10888 23798 10916 26200
rect 11060 24336 11112 24342
rect 11060 24278 11112 24284
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10980 23526 11008 23734
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10508 21888 10560 21894
rect 10612 21865 10640 22102
rect 10508 21830 10560 21836
rect 10598 21856 10654 21865
rect 10520 21434 10548 21830
rect 10598 21791 10654 21800
rect 10796 21622 10824 22578
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10520 21418 10640 21434
rect 10520 21412 10652 21418
rect 10520 21406 10600 21412
rect 10600 21354 10652 21360
rect 10416 21344 10468 21350
rect 10414 21312 10416 21321
rect 10508 21344 10560 21350
rect 10468 21312 10470 21321
rect 10508 21286 10560 21292
rect 10414 21247 10470 21256
rect 10336 21134 10456 21162
rect 10428 19689 10456 21134
rect 10520 21010 10548 21286
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20398 10548 20946
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10612 20534 10640 20742
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10414 19680 10470 19689
rect 10414 19615 10470 19624
rect 10704 18970 10732 21490
rect 10888 21486 10916 22442
rect 11072 22250 11100 24278
rect 11256 24274 11284 26200
rect 11334 24304 11390 24313
rect 11244 24268 11296 24274
rect 11334 24239 11390 24248
rect 11244 24210 11296 24216
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 10980 22222 11100 22250
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10796 19922 10824 20198
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10796 19310 10824 19858
rect 10888 19514 10916 21286
rect 10980 20602 11008 22222
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11072 21010 11100 22034
rect 11164 21350 11192 22646
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11072 20262 11100 20470
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10784 19168 10836 19174
rect 10980 19156 11008 19858
rect 11072 19514 11100 20198
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10836 19128 11008 19156
rect 10784 19110 10836 19116
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18290 10548 18566
rect 10796 18426 10824 19110
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10980 18358 11008 18770
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10968 18352 11020 18358
rect 10968 18294 11020 18300
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10888 18086 10916 18294
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10980 16590 11008 18294
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11072 16726 11100 17750
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11164 16590 11192 19654
rect 11256 17882 11284 22374
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 15910 10824 16390
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10414 15600 10470 15609
rect 10414 15535 10416 15544
rect 10468 15535 10470 15544
rect 10416 15506 10468 15512
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9416 15162 9444 15438
rect 10244 15162 10272 15438
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10506 15056 10562 15065
rect 10506 14991 10508 15000
rect 10560 14991 10562 15000
rect 10508 14962 10560 14968
rect 10322 14920 10378 14929
rect 10322 14855 10324 14864
rect 10376 14855 10378 14864
rect 10324 14826 10376 14832
rect 10520 14618 10548 14962
rect 10704 14958 10732 15370
rect 10968 15360 11020 15366
rect 10966 15328 10968 15337
rect 11020 15328 11022 15337
rect 10966 15263 11022 15272
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 8850 14512 8906 14521
rect 8850 14447 8906 14456
rect 10704 14414 10732 14894
rect 11072 14822 11100 15982
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 14890 11192 15302
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 13190 10732 14350
rect 10980 13841 11008 14758
rect 11348 14074 11376 24239
rect 11624 23186 11652 26200
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 23866 11744 24550
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11992 23662 12020 26200
rect 12360 24342 12388 26200
rect 12714 26200 12770 26302
rect 12820 26302 13138 26330
rect 12624 26182 12676 26188
rect 12530 24440 12586 24449
rect 12530 24375 12586 24384
rect 12348 24336 12400 24342
rect 12348 24278 12400 24284
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12070 23896 12126 23905
rect 12070 23831 12126 23840
rect 12084 23730 12112 23831
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11886 23352 11942 23361
rect 11886 23287 11942 23296
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11612 21616 11664 21622
rect 11610 21584 11612 21593
rect 11664 21584 11666 21593
rect 11610 21519 11666 21528
rect 11900 20992 11928 23287
rect 12452 23202 12480 24210
rect 12544 24206 12572 24375
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12636 23361 12664 23462
rect 12622 23352 12678 23361
rect 12622 23287 12678 23296
rect 12256 23180 12308 23186
rect 12452 23174 12664 23202
rect 12256 23122 12308 23128
rect 12268 22778 12296 23122
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11978 21856 12034 21865
rect 11978 21791 12034 21800
rect 11808 20964 11928 20992
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11440 19786 11468 19994
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11532 19417 11560 19926
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19514 11652 19790
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11518 19408 11574 19417
rect 11518 19343 11574 19352
rect 11808 19310 11836 20964
rect 11992 20534 12020 21791
rect 12084 21690 12112 21966
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 12084 20097 12112 21286
rect 12070 20088 12126 20097
rect 12070 20023 12126 20032
rect 11886 19408 11942 19417
rect 11886 19343 11942 19352
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11440 17542 11468 19110
rect 11808 18766 11836 19110
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11704 18624 11756 18630
rect 11518 18592 11574 18601
rect 11704 18566 11756 18572
rect 11518 18527 11574 18536
rect 11428 17536 11480 17542
rect 11426 17504 11428 17513
rect 11480 17504 11482 17513
rect 11426 17439 11482 17448
rect 11532 16114 11560 18527
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11624 17610 11652 18022
rect 11716 17746 11744 18566
rect 11808 18358 11836 18702
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11624 17270 11652 17546
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11716 17202 11744 17682
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11716 16046 11744 16526
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11716 14958 11744 15982
rect 11808 15638 11836 16458
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11900 14074 11928 19343
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18426 12112 19246
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12268 17921 12296 22374
rect 12452 22098 12480 22510
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 12360 20777 12388 21354
rect 12452 21321 12480 21354
rect 12438 21312 12494 21321
rect 12438 21247 12494 21256
rect 12440 20800 12492 20806
rect 12346 20768 12402 20777
rect 12440 20742 12492 20748
rect 12346 20703 12402 20712
rect 12452 20602 12480 20742
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 19786 12480 20198
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12438 19680 12494 19689
rect 12438 19615 12494 19624
rect 12452 19174 12480 19615
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12544 19009 12572 22918
rect 12636 19446 12664 23174
rect 12728 22778 12756 23530
rect 12820 22982 12848 26302
rect 13082 26200 13138 26302
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26330 14242 27000
rect 13924 26302 14242 26330
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13360 23520 13412 23526
rect 13358 23488 13360 23497
rect 13412 23488 13414 23497
rect 12950 23420 13258 23429
rect 13358 23423 13414 23432
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 13280 22778 13308 23258
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13004 22438 13032 22578
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 12992 22432 13044 22438
rect 13372 22409 13400 22442
rect 12992 22374 13044 22380
rect 13358 22400 13414 22409
rect 12950 22332 13258 22341
rect 13358 22335 13414 22344
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13464 22234 13492 26200
rect 13832 23905 13860 26200
rect 13818 23896 13874 23905
rect 13818 23831 13874 23840
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22681 13584 22918
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 13634 22128 13690 22137
rect 12728 21894 12756 22102
rect 13556 22072 13634 22094
rect 13556 22066 13690 22072
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12728 21078 12756 21830
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12716 21072 12768 21078
rect 12716 21014 12768 21020
rect 12820 21010 12848 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21049 13400 21830
rect 13464 21350 13492 21966
rect 13556 21962 13584 22066
rect 13634 22063 13690 22066
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13740 21842 13768 23054
rect 13924 23050 13952 26302
rect 14186 26200 14242 26302
rect 14554 26200 14610 27000
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15658 26200 15714 27000
rect 16026 26330 16082 27000
rect 15764 26302 16082 26330
rect 14555 26058 14583 26200
rect 14555 26030 14596 26058
rect 14568 24614 14596 26030
rect 14832 24676 14884 24682
rect 14832 24618 14884 24624
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14016 23866 14044 24142
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14462 23080 14518 23089
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13740 21814 13860 21842
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13634 21448 13690 21457
rect 13544 21412 13596 21418
rect 13634 21383 13690 21392
rect 13544 21354 13596 21360
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13358 21040 13414 21049
rect 12808 21004 12860 21010
rect 13358 20975 13414 20984
rect 12808 20946 12860 20952
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12806 20768 12862 20777
rect 12806 20703 12862 20712
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12530 19000 12586 19009
rect 12530 18935 12586 18944
rect 12728 18714 12756 20334
rect 12636 18686 12756 18714
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12254 17912 12310 17921
rect 12254 17847 12310 17856
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17270 12020 17478
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 16998 12020 17206
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12162 16280 12218 16289
rect 12162 16215 12218 16224
rect 12176 15706 12204 16215
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12268 15366 12296 16594
rect 12360 16454 12388 18158
rect 12452 18086 12480 18158
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12636 17746 12664 18686
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 16522 12572 17478
rect 12636 17134 12664 17682
rect 12728 17610 12756 18566
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 17270 12756 17546
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12728 16522 12756 17206
rect 12532 16516 12584 16522
rect 12716 16516 12768 16522
rect 12532 16458 12584 16464
rect 12636 16476 12716 16504
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12360 16046 12388 16390
rect 12636 16182 12664 16476
rect 12716 16458 12768 16464
rect 12624 16176 12676 16182
rect 12438 16144 12494 16153
rect 12624 16118 12676 16124
rect 12438 16079 12494 16088
rect 12452 16046 12480 16079
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12348 15632 12400 15638
rect 12346 15600 12348 15609
rect 12544 15609 12572 15642
rect 12400 15600 12402 15609
rect 12346 15535 12402 15544
rect 12530 15600 12586 15609
rect 12530 15535 12586 15544
rect 12636 15434 12664 16118
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12256 15360 12308 15366
rect 12348 15360 12400 15366
rect 12256 15302 12308 15308
rect 12346 15328 12348 15337
rect 12400 15328 12402 15337
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 10966 13832 11022 13841
rect 10966 13767 11022 13776
rect 12084 13394 12112 14758
rect 12268 14482 12296 15302
rect 12346 15263 12402 15272
rect 12636 15094 12664 15370
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12544 14618 12572 14894
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12636 14346 12664 15030
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 10060 9042 10088 13126
rect 11532 12986 11560 13194
rect 12636 12986 12664 14282
rect 12820 14074 12848 20703
rect 12912 20262 12940 20810
rect 13188 20641 13216 20878
rect 13464 20874 13492 21286
rect 13556 20874 13584 21354
rect 13648 21146 13676 21383
rect 13740 21146 13768 21626
rect 13832 21418 13860 21814
rect 14016 21570 14044 22986
rect 14200 22710 14228 23054
rect 14462 23015 14518 23024
rect 14556 23044 14608 23050
rect 14476 22982 14504 23015
rect 14556 22986 14608 22992
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14568 22778 14596 22986
rect 14752 22778 14780 23598
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14094 22400 14150 22409
rect 14094 22335 14150 22344
rect 13924 21542 14044 21570
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13818 21312 13874 21321
rect 13818 21247 13874 21256
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 21026 13860 21247
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13740 20998 13860 21026
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13360 20800 13412 20806
rect 13358 20768 13360 20777
rect 13556 20777 13584 20810
rect 13412 20768 13414 20777
rect 13358 20703 13414 20712
rect 13542 20768 13598 20777
rect 13542 20703 13598 20712
rect 13174 20632 13230 20641
rect 13174 20567 13176 20576
rect 13228 20567 13230 20576
rect 13358 20632 13414 20641
rect 13358 20567 13414 20576
rect 13176 20538 13228 20544
rect 13372 20330 13400 20567
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 13358 20224 13414 20233
rect 12950 20156 13258 20165
rect 13358 20159 13414 20168
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 19446 13308 19722
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17882 13400 20159
rect 13648 19990 13676 20946
rect 13740 20806 13768 20998
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 19174 13676 19654
rect 13832 19514 13860 20538
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13648 18952 13676 19110
rect 13556 18924 13676 18952
rect 13556 18630 13584 18924
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13464 17882 13492 18566
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13648 17610 13676 18770
rect 13832 18766 13860 19450
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 17746 13768 18634
rect 13832 18426 13860 18702
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13464 16250 13492 17206
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15745 13400 15982
rect 13358 15736 13414 15745
rect 13358 15671 13414 15680
rect 13464 15586 13492 16186
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15638 13584 15846
rect 13280 15570 13492 15586
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13268 15564 13492 15570
rect 13320 15558 13492 15564
rect 13268 15506 13320 15512
rect 13832 15502 13860 17070
rect 13924 16289 13952 21542
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 14016 21049 14044 21422
rect 14002 21040 14058 21049
rect 14108 21010 14136 22335
rect 14200 22030 14228 22646
rect 14370 22536 14426 22545
rect 14370 22471 14426 22480
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14002 20975 14058 20984
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14200 20602 14228 21966
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14094 20088 14150 20097
rect 14094 20023 14150 20032
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 19514 14044 19790
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14002 18048 14058 18057
rect 14002 17983 14058 17992
rect 13910 16280 13966 16289
rect 13910 16215 13966 16224
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13924 15162 13952 16050
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13556 14482 13584 14826
rect 13832 14618 13860 15098
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13636 13932 13688 13938
rect 13832 13920 13860 14214
rect 14016 14074 14044 17983
rect 14108 16810 14136 20023
rect 14292 19854 14320 21558
rect 14384 19990 14412 22471
rect 14752 22234 14780 22714
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14844 22094 14872 24618
rect 14936 23186 14964 26200
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 23798 15240 24754
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 15304 22710 15332 26200
rect 15382 24168 15438 24177
rect 15382 24103 15438 24112
rect 15396 23798 15424 24103
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15672 23322 15700 26200
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15764 23202 15792 26302
rect 16026 26200 16082 26302
rect 16394 26200 16450 27000
rect 16762 26200 16818 27000
rect 17130 26200 17186 27000
rect 17498 26200 17554 27000
rect 17866 26330 17922 27000
rect 17696 26302 17922 26330
rect 16408 24993 16436 26200
rect 16394 24984 16450 24993
rect 16394 24919 16450 24928
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15856 23730 15884 24142
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15396 23174 15792 23202
rect 15396 23050 15424 23174
rect 15384 23044 15436 23050
rect 15384 22986 15436 22992
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15212 22094 15240 22442
rect 14752 22066 14872 22094
rect 15120 22066 15240 22094
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14462 20904 14518 20913
rect 14462 20839 14518 20848
rect 14476 20806 14504 20839
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14568 20398 14596 21830
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14370 19408 14426 19417
rect 14292 18970 14320 19382
rect 14476 19378 14504 19654
rect 14370 19343 14426 19352
rect 14464 19372 14516 19378
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14200 18850 14228 18906
rect 14384 18850 14412 19343
rect 14464 19314 14516 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14200 18822 14412 18850
rect 14384 17202 14412 18822
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14108 16782 14320 16810
rect 14094 16688 14150 16697
rect 14094 16623 14150 16632
rect 14108 15706 14136 16623
rect 14292 15722 14320 16782
rect 14384 16454 14412 17138
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14096 15700 14148 15706
rect 14292 15694 14412 15722
rect 14096 15642 14148 15648
rect 14108 14414 14136 15642
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13688 13892 13860 13920
rect 13636 13874 13688 13880
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 11520 12980 11572 12986
rect 12624 12980 12676 12986
rect 11520 12922 11572 12928
rect 12544 12940 12624 12968
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 12544 8906 12572 12940
rect 12624 12922 12676 12928
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 11830 13400 13398
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 12986 13492 13194
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13832 11898 13860 12922
rect 14108 12442 14136 14214
rect 14200 13258 14228 15506
rect 14292 14482 14320 15506
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14006 14320 14418
rect 14384 14278 14412 15694
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14292 13394 14320 13942
rect 14476 13870 14504 19110
rect 14568 16250 14596 19790
rect 14660 19514 14688 20810
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14752 19174 14780 22066
rect 15120 21729 15148 22066
rect 15580 22030 15608 22578
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15106 21720 15162 21729
rect 15106 21655 15162 21664
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14752 18426 14780 18770
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14646 17776 14702 17785
rect 14646 17711 14702 17720
rect 14660 16969 14688 17711
rect 14752 17105 14780 18022
rect 14738 17096 14794 17105
rect 14738 17031 14794 17040
rect 14646 16960 14702 16969
rect 14646 16895 14702 16904
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 14482 14596 15982
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14660 15094 14688 15370
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14056 14596 14418
rect 14648 14068 14700 14074
rect 14568 14028 14648 14056
rect 14648 14010 14700 14016
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14292 12986 14320 13330
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14384 11830 14412 12038
rect 14568 11898 14596 13194
rect 14844 11898 14872 20878
rect 15014 20496 15070 20505
rect 15014 20431 15070 20440
rect 15028 20398 15056 20431
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15120 20330 15148 21422
rect 15396 20806 15424 21490
rect 15580 21350 15608 21966
rect 15672 21486 15700 22918
rect 16028 22704 16080 22710
rect 16028 22646 16080 22652
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15290 20496 15346 20505
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14936 19514 14964 19722
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14922 19408 14978 19417
rect 14922 19343 14978 19352
rect 14936 18902 14964 19343
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 15028 18834 15056 19722
rect 15120 19310 15148 20266
rect 15212 19378 15240 20470
rect 15290 20431 15346 20440
rect 15304 20097 15332 20431
rect 15290 20088 15346 20097
rect 15290 20023 15346 20032
rect 15396 19786 15424 20742
rect 15580 20534 15608 21286
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19553 15332 19654
rect 15290 19544 15346 19553
rect 15290 19479 15346 19488
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14936 17746 14964 18702
rect 15028 18698 15056 18770
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15014 17776 15070 17785
rect 14924 17740 14976 17746
rect 15014 17711 15070 17720
rect 14924 17682 14976 17688
rect 14936 16658 14964 17682
rect 15028 17202 15056 17711
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16794 15056 16934
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 14752 11286 14780 11766
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 14936 9178 14964 16390
rect 15028 16250 15056 16458
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15028 15026 15056 15846
rect 15120 15314 15148 17002
rect 15212 15706 15240 17546
rect 15382 16824 15438 16833
rect 15382 16759 15438 16768
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15120 15286 15332 15314
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 15120 11558 15148 11727
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 9324 6458 9352 8842
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6748 2854 6776 2994
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6748 800 6776 2790
rect 7208 2446 7236 3334
rect 7484 3194 7512 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 8680 2650 8708 6258
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 15212 5914 15240 12718
rect 15304 8498 15332 15286
rect 15396 14958 15424 16759
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15488 10305 15516 20402
rect 15566 19544 15622 19553
rect 15566 19479 15568 19488
rect 15620 19479 15622 19488
rect 15568 19450 15620 19456
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15672 18630 15700 19178
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 18426 15700 18566
rect 15660 18420 15712 18426
rect 15580 18380 15660 18408
rect 15580 16114 15608 18380
rect 15660 18362 15712 18368
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 12918 15608 13738
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15580 12442 15608 12854
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15672 12322 15700 17682
rect 15764 17592 15792 22510
rect 15934 21856 15990 21865
rect 15934 21791 15990 21800
rect 15948 21486 15976 21791
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 20942 15976 21422
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15948 20806 15976 20878
rect 15844 20800 15896 20806
rect 15842 20768 15844 20777
rect 15936 20800 15988 20806
rect 15896 20768 15898 20777
rect 15936 20742 15988 20748
rect 15842 20703 15898 20712
rect 15934 20360 15990 20369
rect 15934 20295 15990 20304
rect 15948 20262 15976 20295
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15856 20058 15884 20198
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 16040 19938 16068 22646
rect 15856 19910 16068 19938
rect 15856 17746 15884 19910
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15764 17564 15884 17592
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15580 12294 15700 12322
rect 15580 11558 15608 12294
rect 15660 11688 15712 11694
rect 15658 11656 15660 11665
rect 15712 11656 15714 11665
rect 15658 11591 15714 11600
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15658 11248 15714 11257
rect 15658 11183 15714 11192
rect 15672 11150 15700 11183
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15672 10810 15700 11086
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15474 10296 15530 10305
rect 15474 10231 15530 10240
rect 15764 9674 15792 16050
rect 15856 14074 15884 17564
rect 15948 14550 15976 19722
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18698 16068 19246
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 16040 16794 16068 18634
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15026 16068 15982
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15948 14006 15976 14350
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 15948 13734 15976 13942
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12646 15976 13126
rect 15936 12640 15988 12646
rect 16132 12594 16160 23734
rect 16224 22710 16252 24006
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16316 23254 16344 23598
rect 16304 23248 16356 23254
rect 16304 23190 16356 23196
rect 16316 22982 16344 23190
rect 16408 23118 16436 24006
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16684 23118 16712 23462
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16212 22704 16264 22710
rect 16212 22646 16264 22652
rect 16408 22506 16436 23054
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16500 22545 16528 22714
rect 16592 22642 16620 22918
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16486 22536 16542 22545
rect 16396 22500 16448 22506
rect 16486 22471 16542 22480
rect 16396 22442 16448 22448
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16316 22166 16344 22374
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16408 22098 16436 22442
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 16500 22066 16620 22094
rect 16500 21622 16528 22066
rect 16592 21962 16620 22066
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16224 18222 16252 20742
rect 16316 19961 16344 21422
rect 16408 21350 16436 21490
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16408 20806 16436 21286
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16302 19952 16358 19961
rect 16302 19887 16358 19896
rect 16302 19816 16358 19825
rect 16302 19751 16358 19760
rect 16316 19718 16344 19751
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16408 19310 16436 20742
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 19378 16528 20402
rect 16592 19446 16620 21286
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16316 18290 16344 18634
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16316 17678 16344 18226
rect 16408 17746 16436 19110
rect 16486 18320 16542 18329
rect 16486 18255 16542 18264
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 16522 16344 17614
rect 16500 17066 16528 18255
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17338 16620 17478
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16250 16344 16458
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16316 15502 16344 16186
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 15366 16344 15438
rect 16592 15434 16620 16934
rect 16684 16590 16712 22374
rect 16776 21350 16804 26200
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23905 16896 24006
rect 16854 23896 16910 23905
rect 16854 23831 16910 23840
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16868 23322 16896 23462
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17052 22710 17080 23190
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16868 22137 16896 22442
rect 17038 22400 17094 22409
rect 17038 22335 17094 22344
rect 16854 22128 16910 22137
rect 16854 22063 16910 22072
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16868 21146 16896 21830
rect 16960 21729 16988 21830
rect 16946 21720 17002 21729
rect 16946 21655 17002 21664
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16764 21072 16816 21078
rect 16960 21026 16988 21655
rect 17052 21078 17080 22335
rect 16764 21014 16816 21020
rect 16776 20398 16804 21014
rect 16868 20998 16988 21026
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16868 20641 16896 20998
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16854 20632 16910 20641
rect 16854 20567 16910 20576
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 18057 16804 19722
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 19417 16896 19654
rect 16854 19408 16910 19417
rect 16854 19343 16910 19352
rect 16762 18048 16818 18057
rect 16762 17983 16818 17992
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16684 15706 16712 16526
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 15936 12582 15988 12588
rect 15948 11762 15976 12582
rect 16040 12566 16160 12594
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 11286 15976 11698
rect 16040 11354 16068 12566
rect 16118 11384 16174 11393
rect 16028 11348 16080 11354
rect 16118 11319 16120 11328
rect 16028 11290 16080 11296
rect 16172 11319 16174 11328
rect 16120 11290 16172 11296
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15764 9646 15976 9674
rect 15948 9382 15976 9646
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 16224 8362 16252 14486
rect 16316 14414 16344 15302
rect 16776 15094 16804 17682
rect 16854 17504 16910 17513
rect 16854 17439 16910 17448
rect 16868 17338 16896 17439
rect 16856 17332 16908 17338
rect 16960 17320 16988 20878
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 19514 17080 20198
rect 17144 19990 17172 26200
rect 17512 25809 17540 26200
rect 17498 25800 17554 25809
rect 17498 25735 17554 25744
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17236 23526 17264 24006
rect 17328 23730 17356 24346
rect 17420 24274 17448 24754
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17314 23080 17370 23089
rect 17314 23015 17370 23024
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17236 22817 17264 22918
rect 17222 22808 17278 22817
rect 17222 22743 17278 22752
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21865 17264 22034
rect 17222 21856 17278 21865
rect 17222 21791 17278 21800
rect 17328 21690 17356 23015
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17420 21554 17448 23734
rect 17512 21622 17540 24210
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17420 20913 17448 21490
rect 17604 21468 17632 24074
rect 17696 22438 17724 26302
rect 17866 26200 17922 26302
rect 18234 26200 18290 27000
rect 18602 26330 18658 27000
rect 18432 26302 18658 26330
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17788 23662 17816 24754
rect 18248 24138 18276 26200
rect 18432 24886 18460 26302
rect 18602 26200 18658 26302
rect 18970 26200 19026 27000
rect 19338 26330 19394 27000
rect 19260 26302 19394 26330
rect 18984 25945 19012 26200
rect 18970 25936 19026 25945
rect 18970 25871 19026 25880
rect 18696 25016 18748 25022
rect 18696 24958 18748 24964
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18524 23905 18552 24210
rect 18510 23896 18566 23905
rect 18510 23831 18566 23840
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17868 23112 17920 23118
rect 17774 23080 17830 23089
rect 17830 23060 17868 23066
rect 17972 23089 18000 23530
rect 18064 23118 18092 23598
rect 18052 23112 18104 23118
rect 17830 23054 17920 23060
rect 17958 23080 18014 23089
rect 17830 23038 17908 23054
rect 17774 23015 17830 23024
rect 18052 23054 18104 23060
rect 17958 23015 18014 23024
rect 17776 22976 17828 22982
rect 18064 22964 18092 23054
rect 17776 22918 17828 22924
rect 17880 22936 18092 22964
rect 17788 22438 17816 22918
rect 17880 22778 17908 22936
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18432 22710 18460 23734
rect 18708 23186 18736 24958
rect 19260 24750 19288 26302
rect 19338 26200 19394 26302
rect 19706 26200 19762 27000
rect 20074 26200 20130 27000
rect 20442 26330 20498 27000
rect 20180 26302 20498 26330
rect 20180 26217 20208 26302
rect 20166 26208 20222 26217
rect 19720 26081 19748 26200
rect 19706 26072 19762 26081
rect 19706 26007 19762 26016
rect 20088 25673 20116 26200
rect 20442 26200 20498 26302
rect 20810 26200 20866 27000
rect 21178 26200 21234 27000
rect 21546 26200 21602 27000
rect 21914 26200 21970 27000
rect 22282 26200 22338 27000
rect 22650 26330 22706 27000
rect 23018 26330 23074 27000
rect 23386 26330 23442 27000
rect 24490 26330 24546 27000
rect 22388 26302 22706 26330
rect 20166 26143 20222 26152
rect 20074 25664 20130 25673
rect 20074 25599 20130 25608
rect 20536 24880 20588 24886
rect 20536 24822 20588 24828
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 18972 24064 19024 24070
rect 18972 24006 19024 24012
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18524 22778 18552 23122
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18696 22976 18748 22982
rect 18616 22936 18696 22964
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17696 21729 17724 22102
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18420 22092 18472 22098
rect 18616 22094 18644 22936
rect 18800 22953 18828 22986
rect 18696 22918 18748 22924
rect 18786 22944 18842 22953
rect 18786 22879 18842 22888
rect 18892 22642 18920 23734
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18892 22438 18920 22578
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18892 22234 18920 22374
rect 18880 22228 18932 22234
rect 18800 22188 18880 22216
rect 18800 22137 18828 22188
rect 18880 22170 18932 22176
rect 18420 22034 18472 22040
rect 18524 22066 18644 22094
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17682 21720 17738 21729
rect 17788 21690 17816 21898
rect 18156 21894 18184 22034
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17682 21655 17738 21664
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17512 21440 17632 21468
rect 17684 21480 17736 21486
rect 17406 20904 17462 20913
rect 17316 20868 17368 20874
rect 17406 20839 17462 20848
rect 17316 20810 17368 20816
rect 17222 20632 17278 20641
rect 17222 20567 17224 20576
rect 17276 20567 17278 20576
rect 17224 20538 17276 20544
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17328 19802 17356 20810
rect 17144 19774 17356 19802
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17144 19334 17172 19774
rect 17512 19768 17540 21440
rect 17684 21422 17736 21428
rect 17512 19740 17632 19768
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 19553 17264 19654
rect 17222 19544 17278 19553
rect 17604 19496 17632 19740
rect 17222 19479 17278 19488
rect 17512 19468 17632 19496
rect 17406 19348 17462 19357
rect 17144 19306 17264 19334
rect 17236 19145 17264 19306
rect 17316 19304 17368 19310
rect 17406 19283 17462 19292
rect 17316 19246 17368 19252
rect 17222 19136 17278 19145
rect 17222 19071 17278 19080
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 18290 17172 18566
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 16960 17292 17080 17320
rect 16856 17274 16908 17280
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16408 13938 16436 14758
rect 16500 14414 16528 14758
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12170 16344 13126
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16408 11150 16436 13631
rect 16500 13394 16528 14350
rect 16776 14278 16804 15030
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16500 12434 16528 13330
rect 16592 12646 16620 13670
rect 16776 13258 16804 13670
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16868 12850 16896 15506
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16500 12406 16620 12434
rect 16592 11762 16620 12406
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 10810 16436 11086
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16684 10198 16712 12718
rect 16868 12434 16896 12786
rect 16776 12406 16896 12434
rect 16776 12306 16804 12406
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16960 11354 16988 17138
rect 17052 11354 17080 17292
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17144 14822 17172 16594
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17236 14464 17264 18226
rect 17328 17814 17356 19246
rect 17420 18358 17448 19283
rect 17512 18578 17540 19468
rect 17696 19310 17724 21422
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17788 21146 17816 21354
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17696 18630 17724 18770
rect 17684 18624 17736 18630
rect 17512 18550 17632 18578
rect 17684 18566 17736 18572
rect 17498 18456 17554 18465
rect 17498 18391 17554 18400
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17512 18222 17540 18391
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17420 17610 17448 18158
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 15994 17448 17070
rect 17144 14436 17264 14464
rect 17328 15966 17448 15994
rect 17144 14278 17172 14436
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17144 11200 17172 14010
rect 17328 13734 17356 15966
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15094 17448 15846
rect 17408 15088 17460 15094
rect 17408 15030 17460 15036
rect 17512 14074 17540 18022
rect 17604 15978 17632 18550
rect 17696 17542 17724 18566
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17134 17724 17478
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17328 11898 17356 12922
rect 17420 12306 17448 13874
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17604 13190 17632 13806
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17144 11172 17264 11200
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10810 17172 11018
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 17236 9518 17264 11172
rect 17590 10568 17646 10577
rect 17788 10538 17816 20946
rect 17880 20942 17908 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18432 20942 18460 22034
rect 18524 21894 18552 22066
rect 18616 22030 18644 22066
rect 18786 22128 18842 22137
rect 18786 22063 18842 22072
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18512 21888 18564 21894
rect 18512 21830 18564 21836
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17972 19700 18000 19994
rect 18156 19922 18184 20538
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18248 20058 18276 20334
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18236 19916 18288 19922
rect 18288 19876 18368 19904
rect 18236 19858 18288 19864
rect 17880 19672 18000 19700
rect 17880 19496 17908 19672
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 19530 18368 19876
rect 18144 19508 18196 19514
rect 17880 19468 18000 19496
rect 17972 19394 18000 19468
rect 18340 19502 18460 19530
rect 18144 19450 18196 19456
rect 17880 19366 18000 19394
rect 17880 18902 17908 19366
rect 17868 18896 17920 18902
rect 18156 18873 18184 19450
rect 18432 19334 18460 19502
rect 18340 19306 18460 19334
rect 18340 18952 18368 19306
rect 18248 18924 18368 18952
rect 17868 18838 17920 18844
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18248 18612 18276 18924
rect 18328 18828 18380 18834
rect 18380 18788 18460 18816
rect 18328 18770 18380 18776
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 17880 18584 18276 18612
rect 17880 17270 17908 18584
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17972 17649 18000 18294
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 18086 18276 18226
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 18340 17202 18368 18634
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 15348 18000 15642
rect 18340 15638 18368 16390
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17880 15320 18000 15348
rect 17880 14958 17908 15320
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18236 15020 18288 15026
rect 18340 15008 18368 15438
rect 18288 14980 18368 15008
rect 18236 14962 18288 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18248 14346 18276 14962
rect 18236 14340 18288 14346
rect 18236 14282 18288 14288
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17880 12832 17908 13262
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18432 12968 18460 18788
rect 18524 18426 18552 21558
rect 18800 21078 18828 22063
rect 18878 21448 18934 21457
rect 18878 21383 18934 21392
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 20602 18736 20946
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18800 20534 18828 21014
rect 18892 20913 18920 21383
rect 18878 20904 18934 20913
rect 18878 20839 18934 20848
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 19428 18736 19858
rect 18616 19400 18736 19428
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18524 16250 18552 18362
rect 18616 17678 18644 19400
rect 18694 19348 18750 19357
rect 18694 19283 18750 19292
rect 18708 18329 18736 19283
rect 18694 18320 18750 18329
rect 18694 18255 18750 18264
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18524 14006 18552 16186
rect 18616 15502 18644 17478
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14482 18644 14758
rect 18708 14550 18736 18158
rect 18800 17678 18828 19926
rect 18892 18766 18920 20538
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18984 18601 19012 24006
rect 19062 23080 19118 23089
rect 19062 23015 19118 23024
rect 19076 21690 19104 23015
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19168 21418 19196 24074
rect 19340 24064 19392 24070
rect 19338 24032 19340 24041
rect 19524 24064 19576 24070
rect 19392 24032 19394 24041
rect 19394 24012 19524 24018
rect 19394 24006 19576 24012
rect 19394 23990 19564 24006
rect 19338 23967 19394 23976
rect 20548 23746 20576 24822
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20640 23866 20668 24006
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20626 23760 20682 23769
rect 20548 23718 20626 23746
rect 20732 23730 20760 24210
rect 20626 23695 20682 23704
rect 20720 23724 20772 23730
rect 20640 23662 20668 23695
rect 20720 23666 20772 23672
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 19800 23520 19852 23526
rect 19444 23468 19800 23474
rect 19444 23462 19852 23468
rect 19444 23446 19840 23462
rect 19444 23254 19472 23446
rect 19432 23248 19484 23254
rect 19246 23216 19302 23225
rect 19432 23190 19484 23196
rect 19246 23151 19302 23160
rect 19260 22778 19288 23151
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19352 22030 19380 23054
rect 19996 23050 20024 23598
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 20088 23032 20116 23462
rect 20168 23044 20220 23050
rect 20088 23004 20168 23032
rect 20088 22556 20116 23004
rect 20168 22986 20220 22992
rect 20732 22982 20760 23666
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20824 22681 20852 26200
rect 20904 25084 20956 25090
rect 20904 25026 20956 25032
rect 20810 22672 20866 22681
rect 20628 22636 20680 22642
rect 20810 22607 20866 22616
rect 20628 22578 20680 22584
rect 20168 22568 20220 22574
rect 20088 22528 20168 22556
rect 20088 22438 20116 22528
rect 20168 22510 20220 22516
rect 20534 22536 20590 22545
rect 20534 22471 20590 22480
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19340 22024 19392 22030
rect 19444 22001 19472 22170
rect 19340 21966 19392 21972
rect 19430 21992 19486 22001
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19260 20806 19288 21966
rect 19352 21350 19380 21966
rect 19430 21927 19486 21936
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19352 20618 19380 20878
rect 19260 20590 19380 20618
rect 19260 20398 19288 20590
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18970 18592 19026 18601
rect 18970 18527 19026 18536
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18524 13802 18552 13942
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18340 12940 18460 12968
rect 18236 12844 18288 12850
rect 17880 12804 18236 12832
rect 17880 12646 17908 12804
rect 18236 12786 18288 12792
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 18248 12442 18276 12786
rect 18340 12782 18368 12940
rect 18616 12866 18644 14214
rect 18708 13394 18736 14486
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18524 12838 18644 12866
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18248 12238 18276 12378
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11082 18368 12582
rect 18432 11218 18460 12786
rect 18524 12646 18552 12838
rect 18800 12782 18828 17478
rect 18892 17270 18920 17818
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 15570 18920 16390
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18984 15162 19012 16050
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18510 12472 18566 12481
rect 18510 12407 18566 12416
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18064 10713 18092 10746
rect 18050 10704 18106 10713
rect 18524 10674 18552 12407
rect 18616 11694 18644 12650
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18050 10639 18106 10648
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 17590 10503 17646 10512
rect 17776 10532 17828 10538
rect 17604 10062 17632 10503
rect 17776 10474 17828 10480
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 18616 9450 18644 11290
rect 18708 11286 18736 12106
rect 18800 11830 18828 12378
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18800 11082 18828 11766
rect 18892 11150 18920 13126
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 18708 7886 18736 10950
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 8974 18920 9522
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18984 4078 19012 15098
rect 19076 12986 19104 18838
rect 19168 17882 19196 19926
rect 19260 18698 19288 20334
rect 19444 19446 19472 21422
rect 19536 20777 19564 21898
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19800 20800 19852 20806
rect 19522 20768 19578 20777
rect 19800 20742 19852 20748
rect 19522 20703 19578 20712
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19536 18222 19564 19722
rect 19628 18766 19656 20198
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19417 19748 19654
rect 19706 19408 19762 19417
rect 19706 19343 19762 19352
rect 19706 19272 19762 19281
rect 19706 19207 19762 19216
rect 19720 19174 19748 19207
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19708 18624 19760 18630
rect 19812 18612 19840 20742
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19904 19310 19932 20334
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19904 18873 19932 19246
rect 19890 18864 19946 18873
rect 19890 18799 19946 18808
rect 19760 18584 19840 18612
rect 19708 18566 19760 18572
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16454 19196 17070
rect 19260 16574 19288 18022
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 16726 19380 17070
rect 19536 16969 19564 18158
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19522 16960 19578 16969
rect 19522 16895 19578 16904
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19260 16546 19472 16574
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19154 15192 19210 15201
rect 19154 15127 19210 15136
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 4826 19104 12718
rect 19168 12481 19196 15127
rect 19260 14074 19288 15302
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19352 13988 19380 14894
rect 19444 14414 19472 16546
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19536 14113 19564 15302
rect 19522 14104 19578 14113
rect 19522 14039 19578 14048
rect 19352 13960 19472 13988
rect 19444 13734 19472 13960
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19154 12472 19210 12481
rect 19154 12407 19210 12416
rect 19260 12322 19288 12582
rect 19168 12294 19288 12322
rect 19444 12306 19472 13670
rect 19536 13326 19564 13738
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 12300 19484 12306
rect 19168 8566 19196 12294
rect 19432 12242 19484 12248
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 19260 3126 19288 12106
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11898 19380 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19536 11150 19564 13262
rect 19628 12986 19656 17478
rect 19720 16250 19748 18566
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19720 13530 19748 16050
rect 19812 15706 19840 18158
rect 19890 18048 19946 18057
rect 19890 17983 19946 17992
rect 19904 17882 19932 17983
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 19904 17746 19932 17818
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19812 14006 19840 14758
rect 19800 14000 19852 14006
rect 19800 13942 19852 13948
rect 19812 13530 19840 13942
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19522 10704 19578 10713
rect 19522 10639 19578 10648
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19352 6866 19380 10406
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19444 9654 19472 9998
rect 19536 9926 19564 10639
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19430 9480 19486 9489
rect 19430 9415 19432 9424
rect 19484 9415 19486 9424
rect 19432 9386 19484 9392
rect 19536 9178 19564 9522
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19628 8634 19656 11834
rect 19720 11830 19748 13262
rect 19904 13258 19932 15982
rect 19996 15366 20024 21286
rect 20088 17134 20116 21830
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20180 16640 20208 20334
rect 20088 16612 20208 16640
rect 20088 16153 20116 16612
rect 20166 16416 20222 16425
rect 20166 16351 20222 16360
rect 20074 16144 20130 16153
rect 20074 16079 20130 16088
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19798 12472 19854 12481
rect 19798 12407 19854 12416
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19706 11112 19762 11121
rect 19706 11047 19762 11056
rect 19720 10810 19748 11047
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19720 10266 19748 10406
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9722 19748 9998
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19812 7954 19840 12407
rect 19890 12336 19946 12345
rect 19890 12271 19946 12280
rect 19904 11150 19932 12271
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 8974 19932 11086
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19996 4146 20024 13806
rect 20088 11150 20116 14486
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20088 10674 20116 10746
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20180 10606 20208 16351
rect 20272 13705 20300 22374
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20456 20641 20484 21490
rect 20442 20632 20498 20641
rect 20442 20567 20498 20576
rect 20548 20262 20576 22471
rect 20640 21593 20668 22578
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20732 21060 20760 21626
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20640 21032 20760 21060
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20640 19990 20668 21032
rect 20824 20369 20852 21490
rect 20916 20618 20944 25026
rect 21192 23361 21220 26200
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 21178 23352 21234 23361
rect 21178 23287 21234 23296
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20996 22500 21048 22506
rect 20996 22442 21048 22448
rect 21008 21486 21036 22442
rect 21100 21962 21128 22510
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21100 20874 21128 21898
rect 21192 21078 21220 23122
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21088 20868 21140 20874
rect 21140 20828 21220 20856
rect 21088 20810 21140 20816
rect 20916 20590 21036 20618
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20810 20360 20866 20369
rect 20720 20324 20772 20330
rect 20810 20295 20866 20304
rect 20720 20266 20772 20272
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20732 19922 20760 20266
rect 20916 20058 20944 20470
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20718 19816 20774 19825
rect 20352 19304 20404 19310
rect 20350 19272 20352 19281
rect 20404 19272 20406 19281
rect 20350 19207 20406 19216
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18426 20392 19110
rect 20534 18456 20590 18465
rect 20352 18420 20404 18426
rect 20534 18391 20590 18400
rect 20352 18362 20404 18368
rect 20548 18358 20576 18391
rect 20536 18352 20588 18358
rect 20442 18320 20498 18329
rect 20536 18294 20588 18300
rect 20442 18255 20444 18264
rect 20496 18255 20498 18264
rect 20444 18226 20496 18232
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20258 13696 20314 13705
rect 20258 13631 20314 13640
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 9489 20208 9522
rect 20166 9480 20222 9489
rect 20166 9415 20222 9424
rect 20272 7410 20300 12582
rect 20364 12102 20392 17682
rect 20548 14634 20576 18090
rect 20640 16998 20668 19790
rect 20718 19751 20774 19760
rect 20732 18222 20760 19751
rect 21008 19666 21036 20590
rect 21192 20346 21220 20828
rect 21284 20602 21312 22170
rect 21376 21690 21404 23462
rect 21468 21706 21496 24142
rect 21560 22409 21588 26200
rect 21928 23497 21956 26200
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 21914 23488 21970 23497
rect 21914 23423 21970 23432
rect 21730 23080 21786 23089
rect 21730 23015 21786 23024
rect 21916 23044 21968 23050
rect 21546 22400 21602 22409
rect 21546 22335 21602 22344
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21364 21684 21416 21690
rect 21468 21678 21588 21706
rect 21364 21626 21416 21632
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21376 20602 21404 20742
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21192 20318 21404 20346
rect 21376 20262 21404 20318
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 20916 19638 21036 19666
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17882 20760 18022
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20810 17640 20866 17649
rect 20810 17575 20866 17584
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20732 16726 20760 17478
rect 20720 16720 20772 16726
rect 20824 16697 20852 17575
rect 20720 16662 20772 16668
rect 20810 16688 20866 16697
rect 20810 16623 20866 16632
rect 20810 16144 20866 16153
rect 20916 16114 20944 19638
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21008 19174 21036 19450
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18442 21036 19110
rect 21100 18698 21128 19178
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21008 18414 21128 18442
rect 20996 18352 21048 18358
rect 20994 18320 20996 18329
rect 21048 18320 21050 18329
rect 20994 18255 21050 18264
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20810 16079 20866 16088
rect 20904 16108 20956 16114
rect 20824 15910 20852 16079
rect 20904 16050 20956 16056
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 15366 20944 15438
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20548 14606 20668 14634
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20548 14278 20576 14486
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20548 14074 20576 14214
rect 20640 14074 20668 14606
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20548 13734 20576 14010
rect 20732 13938 20760 14826
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 12102 20484 12650
rect 20548 12646 20576 13670
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11694 20484 12038
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20364 10470 20392 10610
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 19536 2514 19564 2926
rect 19812 2854 19840 2994
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19812 2650 19840 2790
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 4014
rect 20548 3534 20576 11018
rect 20732 10674 20760 13670
rect 20824 12345 20852 15302
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 14006 20944 14214
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21008 13530 21036 18158
rect 21100 16250 21128 18414
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20996 13252 21048 13258
rect 20916 13212 20996 13240
rect 20916 12646 20944 13212
rect 20996 13194 21048 13200
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20812 12232 20864 12238
rect 20916 12220 20944 12582
rect 21100 12458 21128 15914
rect 21192 15570 21220 19450
rect 21376 19378 21404 20198
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21284 18222 21312 19314
rect 21362 19272 21418 19281
rect 21362 19207 21418 19216
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21376 17921 21404 19207
rect 21468 18358 21496 21558
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21362 17912 21418 17921
rect 21362 17847 21418 17856
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21284 17134 21312 17546
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16590 21312 16934
rect 21272 16584 21324 16590
rect 21468 16538 21496 18294
rect 21560 17270 21588 21678
rect 21652 21622 21680 21830
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 19718 21680 20946
rect 21744 20777 21772 23015
rect 21916 22986 21968 22992
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21836 22574 21864 22918
rect 21824 22568 21876 22574
rect 21824 22510 21876 22516
rect 21928 21962 21956 22986
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 20942 21956 21286
rect 22020 21162 22048 24006
rect 22112 23662 22140 24346
rect 22296 24290 22324 26200
rect 22388 24954 22416 26302
rect 22650 26200 22706 26302
rect 22756 26302 23074 26330
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22204 24262 22324 24290
rect 22560 24268 22612 24274
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22112 21298 22140 22442
rect 22204 22273 22232 24262
rect 22560 24210 22612 24216
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23662 22324 24142
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22296 23186 22324 23598
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22190 22264 22246 22273
rect 22190 22199 22246 22208
rect 22388 22166 22416 23462
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22204 21418 22232 21626
rect 22192 21412 22244 21418
rect 22192 21354 22244 21360
rect 22112 21270 22232 21298
rect 22020 21134 22140 21162
rect 22112 21049 22140 21134
rect 22098 21040 22154 21049
rect 22098 20975 22154 20984
rect 22112 20942 22140 20975
rect 21916 20936 21968 20942
rect 21836 20896 21916 20924
rect 21730 20768 21786 20777
rect 21730 20703 21786 20712
rect 21836 20346 21864 20896
rect 21916 20878 21968 20884
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21744 20318 21864 20346
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 18902 21680 19654
rect 21744 19334 21772 20318
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 19786 21864 20198
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21744 19306 21864 19334
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21638 17912 21694 17921
rect 21638 17847 21694 17856
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21272 16526 21324 16532
rect 21376 16510 21496 16538
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15570 21312 16390
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21376 15162 21404 16510
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21284 14890 21312 15098
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21376 14414 21404 15098
rect 21468 15094 21496 16390
rect 21560 15094 21588 16662
rect 21652 15638 21680 17847
rect 21744 16794 21772 19178
rect 21836 18290 21864 19306
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21836 17134 21864 18090
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21836 16998 21864 17070
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21468 14822 21496 15030
rect 21744 14958 21772 16730
rect 21836 16522 21864 16934
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21928 16250 21956 20538
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14550 21496 14758
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21376 12986 21404 14350
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21468 13530 21496 13806
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21100 12430 21220 12458
rect 21086 12336 21142 12345
rect 21086 12271 21142 12280
rect 20864 12192 20944 12220
rect 20812 12174 20864 12180
rect 20824 11762 20852 12174
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20824 11014 20852 11698
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20718 10296 20774 10305
rect 20718 10231 20774 10240
rect 20732 10198 20760 10231
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 7478 20760 7686
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20824 6798 20852 10406
rect 21008 10062 21036 10678
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21008 9466 21036 9998
rect 20916 9438 21036 9466
rect 20916 8634 20944 9438
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 21008 8566 21036 9318
rect 21100 8974 21128 12271
rect 21192 11898 21220 12430
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 9994 21220 11834
rect 21284 11626 21312 12038
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10130 21312 10406
rect 21376 10130 21404 12242
rect 21454 11928 21510 11937
rect 21454 11863 21510 11872
rect 21468 11558 21496 11863
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21468 11218 21496 11494
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21468 9586 21496 10950
rect 21560 10810 21588 14486
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21652 11218 21680 12786
rect 21744 12345 21772 13942
rect 21928 13394 21956 14418
rect 22020 14278 22048 19246
rect 22204 19174 22232 21270
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 18766 22232 19110
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22112 18154 22140 18702
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22204 17882 22232 18566
rect 22296 17921 22324 21626
rect 22388 21554 22416 21966
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22480 21146 22508 24074
rect 22572 23662 22600 24210
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 21350 22600 23462
rect 22664 22438 22692 24550
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22388 20942 22416 21082
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22664 20754 22692 22102
rect 22388 20726 22692 20754
rect 22388 20466 22416 20726
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22388 19514 22416 20402
rect 22480 20262 22508 20538
rect 22572 20398 22600 20538
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22558 19136 22614 19145
rect 22558 19071 22614 19080
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22282 17912 22338 17921
rect 22192 17876 22244 17882
rect 22282 17847 22338 17856
rect 22192 17818 22244 17824
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22112 14890 22140 17206
rect 22204 16046 22232 17818
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22296 16794 22324 17138
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15706 22232 15846
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 22098 14376 22154 14385
rect 22098 14311 22154 14320
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21822 13016 21878 13025
rect 21822 12951 21878 12960
rect 21730 12336 21786 12345
rect 21730 12271 21786 12280
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21652 10266 21680 10542
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21744 9586 21772 11834
rect 21836 10418 21864 12951
rect 21928 12850 21956 13330
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 12306 21956 12786
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22020 10674 22048 14010
rect 22112 13938 22140 14311
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22204 13376 22232 15030
rect 22296 15026 22324 16594
rect 22388 16114 22416 16934
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15609 22416 16050
rect 22374 15600 22430 15609
rect 22374 15535 22430 15544
rect 22374 15464 22430 15473
rect 22374 15399 22376 15408
rect 22428 15399 22430 15408
rect 22376 15370 22428 15376
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14482 22324 14962
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22296 13938 22324 14418
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22480 13682 22508 18770
rect 22572 18698 22600 19071
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22558 18592 22614 18601
rect 22558 18527 22614 18536
rect 22572 18086 22600 18527
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22664 17882 22692 20334
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 17202 22600 17682
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22664 16658 22692 17818
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22756 15994 22784 26302
rect 23018 26200 23074 26302
rect 23124 26302 23442 26330
rect 22836 24676 22888 24682
rect 22836 24618 22888 24624
rect 22848 23633 22876 24618
rect 23124 24614 23152 26302
rect 23386 26200 23442 26302
rect 24044 26302 24546 26330
rect 23386 25664 23442 25673
rect 23386 25599 23442 25608
rect 23294 25528 23350 25537
rect 23294 25463 23350 25472
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24426 23336 25463
rect 23400 24886 23428 25599
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23386 24440 23442 24449
rect 23308 24398 23386 24426
rect 23386 24375 23442 24384
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22940 23866 22968 24006
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 23296 23656 23348 23662
rect 22834 23624 22890 23633
rect 23348 23604 23428 23610
rect 23296 23598 23428 23604
rect 23308 23582 23428 23598
rect 22834 23559 22890 23568
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23400 23254 23428 23582
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23308 22574 23336 23122
rect 23756 23044 23808 23050
rect 23756 22986 23808 22992
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 21554 23336 22510
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 18766 22876 21286
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23112 20936 23164 20942
rect 23204 20936 23256 20942
rect 23112 20878 23164 20884
rect 23202 20904 23204 20913
rect 23256 20904 23258 20913
rect 23124 20806 23152 20878
rect 23202 20839 23258 20848
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23308 20466 23336 21490
rect 23386 21448 23442 21457
rect 23386 21383 23442 21392
rect 23400 20874 23428 21383
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19922 23336 20402
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19378 23336 19858
rect 23492 19854 23520 22034
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 22926 18864 22982 18873
rect 23110 18864 23166 18873
rect 22982 18822 23060 18850
rect 22926 18799 22982 18808
rect 22836 18760 22888 18766
rect 22834 18728 22836 18737
rect 22888 18728 22890 18737
rect 22834 18663 22890 18672
rect 23032 18630 23060 18822
rect 23110 18799 23166 18808
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22848 17882 22876 18566
rect 23124 18426 23152 18799
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23216 18329 23244 18906
rect 23308 18426 23336 19314
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23202 18320 23258 18329
rect 23202 18255 23258 18264
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 23308 17762 23336 18362
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23400 17785 23428 18090
rect 23216 17746 23336 17762
rect 23204 17740 23336 17746
rect 23256 17734 23336 17740
rect 23386 17776 23442 17785
rect 23386 17711 23442 17720
rect 23204 17682 23256 17688
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23110 17504 23166 17513
rect 23110 17439 23166 17448
rect 23124 17338 23152 17439
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16776 23428 17614
rect 23308 16748 23428 16776
rect 22834 16552 22890 16561
rect 22834 16487 22890 16496
rect 22112 13348 22232 13376
rect 22296 13654 22508 13682
rect 22572 15966 22784 15994
rect 22112 12646 22140 13348
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22204 12986 22232 13194
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22190 12880 22246 12889
rect 22190 12815 22246 12824
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11898 22140 12174
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11336 22232 12815
rect 22296 12782 22324 13654
rect 22572 13512 22600 15966
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22664 14074 22692 15846
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22756 15450 22784 15642
rect 22848 15570 22876 16487
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22756 15422 22876 15450
rect 22742 14512 22798 14521
rect 22742 14447 22798 14456
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22650 13832 22706 13841
rect 22650 13767 22706 13776
rect 22480 13484 22600 13512
rect 22480 12889 22508 13484
rect 22558 13424 22614 13433
rect 22558 13359 22614 13368
rect 22572 12918 22600 13359
rect 22560 12912 22612 12918
rect 22466 12880 22522 12889
rect 22560 12854 22612 12860
rect 22466 12815 22522 12824
rect 22284 12776 22336 12782
rect 22664 12730 22692 13767
rect 22756 13734 22784 14447
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22848 13546 22876 15422
rect 22940 15337 22968 15642
rect 23018 15464 23074 15473
rect 23018 15399 23074 15408
rect 22926 15328 22982 15337
rect 22926 15263 22982 15272
rect 23032 15094 23060 15399
rect 23308 15314 23336 16748
rect 23386 16688 23442 16697
rect 23386 16623 23442 16632
rect 23216 15286 23336 15314
rect 23020 15088 23072 15094
rect 23216 15065 23244 15286
rect 23400 15144 23428 16623
rect 23308 15116 23428 15144
rect 23020 15030 23072 15036
rect 23202 15056 23258 15065
rect 23202 14991 23258 15000
rect 23204 14952 23256 14958
rect 23308 14940 23336 15116
rect 23386 15056 23442 15065
rect 23386 14991 23442 15000
rect 23256 14912 23336 14940
rect 23204 14894 23256 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22284 12718 22336 12724
rect 22296 12594 22324 12718
rect 22572 12702 22692 12730
rect 22756 13518 22876 13546
rect 22296 12566 22416 12594
rect 22388 12442 22416 12566
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22112 11308 22232 11336
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21836 10390 21956 10418
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21454 8392 21510 8401
rect 21454 8327 21510 8336
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 21284 7546 21312 7783
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21468 7410 21496 8327
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 7886 21588 8230
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 21468 6458 21496 7346
rect 21652 6662 21680 8910
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21744 5778 21772 8298
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21836 5710 21864 10202
rect 21928 8498 21956 10390
rect 22112 9722 22140 11308
rect 22190 11248 22246 11257
rect 22190 11183 22192 11192
rect 22244 11183 22246 11192
rect 22192 11154 22244 11160
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22112 8090 22140 8842
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22480 6914 22508 11630
rect 22572 10810 22600 12702
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22664 9738 22692 12582
rect 22756 11150 22784 13518
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 23308 10826 23336 14758
rect 23400 14346 23428 14991
rect 23492 14482 23520 19654
rect 23584 19446 23612 22918
rect 23768 22778 23796 22986
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23676 21622 23704 22374
rect 23860 22234 23888 24210
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23952 23798 23980 24074
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23952 22778 23980 23734
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23952 21622 23980 22714
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23676 20534 23704 20946
rect 23768 20641 23796 21286
rect 23952 21078 23980 21558
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23754 20632 23810 20641
rect 23754 20567 23810 20576
rect 23768 20534 23796 20567
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23676 19292 23704 19790
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19417 23796 19654
rect 23754 19408 23810 19417
rect 23754 19343 23810 19352
rect 23584 19264 23704 19292
rect 23584 17610 23612 19264
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23676 17338 23704 17614
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23570 16280 23626 16289
rect 23860 16250 23888 20198
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23952 17746 23980 19994
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23570 16215 23626 16224
rect 23848 16244 23900 16250
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23388 14000 23440 14006
rect 23440 13948 23520 13954
rect 23388 13942 23520 13948
rect 23400 13926 23520 13942
rect 23492 13530 23520 13926
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23584 12730 23612 16215
rect 23848 16186 23900 16192
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23400 12702 23612 12730
rect 23400 11898 23428 12702
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23308 10798 23428 10826
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22572 9710 22692 9738
rect 22572 9110 22600 9710
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22296 6886 22508 6914
rect 22190 6352 22246 6361
rect 22190 6287 22246 6296
rect 22204 5710 22232 6287
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22296 4622 22324 6886
rect 22664 4622 22692 9551
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 1170 22048 3402
rect 22112 1601 22140 4014
rect 22296 3058 22324 4422
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22756 2666 22784 10134
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22848 6798 22876 9386
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23308 4622 23336 7142
rect 23400 5234 23428 10798
rect 23492 9489 23520 11222
rect 23478 9480 23534 9489
rect 23478 9415 23534 9424
rect 23584 8022 23612 11698
rect 23676 9042 23704 14214
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 5710 23520 7686
rect 23768 6866 23796 16050
rect 23952 16046 23980 16390
rect 24044 16114 24072 26302
rect 24490 26200 24546 26302
rect 24858 26200 24914 27000
rect 25226 26200 25282 27000
rect 25318 26480 25374 26489
rect 25318 26415 25374 26424
rect 24214 26072 24270 26081
rect 24214 26007 24270 26016
rect 24124 24812 24176 24818
rect 24124 24754 24176 24760
rect 24136 24070 24164 24754
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 22574 24164 24006
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24228 22030 24256 26007
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25148 24721 25176 25191
rect 25134 24712 25190 24721
rect 25134 24647 25190 24656
rect 25044 24200 25096 24206
rect 25042 24168 25044 24177
rect 25096 24168 25098 24177
rect 25042 24103 25098 24112
rect 24860 24064 24912 24070
rect 24912 24024 25084 24052
rect 24860 24006 24912 24012
rect 24858 23896 24914 23905
rect 24858 23831 24914 23840
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24136 19786 24164 21014
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24136 19446 24164 19722
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24122 18864 24178 18873
rect 24122 18799 24178 18808
rect 24136 18766 24164 18799
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 24136 17542 24164 18362
rect 24228 17542 24256 21966
rect 24320 19718 24348 23598
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22137 24624 22918
rect 24780 22438 24808 23054
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24582 22128 24638 22137
rect 24582 22063 24638 22072
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24412 20534 24440 21014
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 24320 18193 24348 18294
rect 24306 18184 24362 18193
rect 24306 18119 24362 18128
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24136 17270 24164 17478
rect 24320 17338 24348 17682
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24136 16522 24164 17206
rect 24124 16516 24176 16522
rect 24176 16476 24256 16504
rect 24124 16458 24176 16464
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 24122 16008 24178 16017
rect 23952 15162 23980 15982
rect 24122 15943 24178 15952
rect 24136 15706 24164 15943
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23860 14006 23888 14486
rect 23938 14240 23994 14249
rect 23938 14175 23994 14184
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23860 13462 23888 13942
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23860 12918 23888 13398
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23952 12186 23980 14175
rect 24044 12918 24072 15574
rect 24136 14414 24164 15642
rect 24228 15026 24256 16476
rect 24306 15872 24362 15881
rect 24306 15807 24362 15816
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14550 24256 14962
rect 24216 14544 24268 14550
rect 24216 14486 24268 14492
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24320 14226 24348 15807
rect 24412 15162 24440 19858
rect 24504 17678 24532 21830
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24688 20942 24716 21422
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24872 20806 24900 23831
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24766 20496 24822 20505
rect 24766 20431 24822 20440
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24596 19553 24624 19654
rect 24780 19553 24808 20431
rect 24858 19952 24914 19961
rect 24858 19887 24914 19896
rect 24582 19544 24638 19553
rect 24582 19479 24638 19488
rect 24766 19544 24822 19553
rect 24766 19479 24822 19488
rect 24872 19394 24900 19887
rect 24780 19366 24900 19394
rect 24676 19236 24728 19242
rect 24676 19178 24728 19184
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18057 24624 18566
rect 24688 18426 24716 19178
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24492 17536 24544 17542
rect 24492 17478 24544 17484
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24136 14198 24348 14226
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 23860 12158 23980 12186
rect 23860 11694 23888 12158
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23952 10674 23980 12038
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23846 10024 23902 10033
rect 23846 9959 23902 9968
rect 23860 9926 23888 9959
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23952 9586 23980 10474
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23492 3534 23520 5510
rect 23860 5234 23888 8774
rect 24044 8294 24072 12582
rect 24136 10062 24164 14198
rect 24412 13870 24440 15098
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24504 13682 24532 17478
rect 24596 16425 24624 17478
rect 24582 16416 24638 16425
rect 24582 16351 24638 16360
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24596 15706 24624 16050
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24596 13870 24624 14418
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24320 13654 24532 13682
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24228 10130 24256 12174
rect 24320 11082 24348 13654
rect 24596 12306 24624 13806
rect 24688 12850 24716 18158
rect 24780 14618 24808 19366
rect 24964 19258 24992 22918
rect 25056 19922 25084 24024
rect 25148 23798 25176 24647
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25332 23050 25360 26415
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25148 19922 25176 21898
rect 25424 21434 25452 22102
rect 25332 21406 25452 21434
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 24872 19230 24992 19258
rect 25056 19242 25084 19722
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25044 19236 25096 19242
rect 24872 17882 24900 19230
rect 25044 19178 25096 19184
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24964 16153 24992 18566
rect 24950 16144 25006 16153
rect 24950 16079 25006 16088
rect 25056 15722 25084 18906
rect 25148 17270 25176 19450
rect 25240 19310 25268 20198
rect 25332 19514 25360 21406
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 25424 20602 25452 21286
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25240 18834 25268 19246
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25516 18222 25544 23802
rect 25872 23588 25924 23594
rect 25872 23530 25924 23536
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 16250 25268 16526
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 24872 15694 25084 15722
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24780 12918 24808 13398
rect 24872 13394 24900 15694
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24780 12696 24808 12854
rect 24688 12668 24808 12696
rect 24688 12442 24716 12668
rect 24766 12608 24822 12617
rect 24766 12543 24822 12552
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24674 12200 24730 12209
rect 24674 12135 24730 12144
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24308 11076 24360 11082
rect 24308 11018 24360 11024
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 9178 24164 9998
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24504 7886 24532 11290
rect 24688 10606 24716 12135
rect 24780 11694 24808 12543
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24872 11218 24900 11319
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24582 10160 24638 10169
rect 24582 10095 24638 10104
rect 24596 8430 24624 10095
rect 24780 9518 24808 10911
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24872 10577 24900 10678
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24872 9042 24900 9279
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24688 7342 24716 8871
rect 24860 8560 24912 8566
rect 24858 8528 24860 8537
rect 24912 8528 24914 8537
rect 24964 8498 24992 15370
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25148 14929 25176 14962
rect 25134 14920 25190 14929
rect 25134 14855 25190 14864
rect 25320 14884 25372 14890
rect 25148 14618 25176 14855
rect 25320 14826 25372 14832
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25134 13968 25190 13977
rect 25134 13903 25136 13912
rect 25188 13903 25190 13912
rect 25136 13874 25188 13880
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25148 12986 25176 13330
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25042 12336 25098 12345
rect 25042 12271 25044 12280
rect 25096 12271 25098 12280
rect 25044 12242 25096 12248
rect 25136 11688 25188 11694
rect 25134 11656 25136 11665
rect 25188 11656 25190 11665
rect 25134 11591 25190 11600
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 24858 8463 24914 8472
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24950 8120 25006 8129
rect 24950 8055 25006 8064
rect 24964 7954 24992 8055
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 24596 3534 24624 5782
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 25056 6914 25084 8842
rect 24858 6896 24914 6905
rect 24858 6831 24860 6840
rect 24912 6831 24914 6840
rect 24964 6886 25084 6914
rect 24860 6802 24912 6808
rect 24964 6458 24992 6886
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24950 5672 25006 5681
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24860 5296 24912 5302
rect 24766 5264 24822 5273
rect 24860 5238 24912 5244
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24780 4078 24808 5199
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 25056 4146 25084 6666
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25134 4040 25190 4049
rect 24952 4004 25004 4010
rect 25134 3975 25190 3984
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22664 2638 22784 2666
rect 22664 2446 22692 2638
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22756 2009 22784 2450
rect 24596 2446 24624 3334
rect 24964 3233 24992 3402
rect 24950 3224 25006 3233
rect 24950 3159 25006 3168
rect 25148 3126 25176 3975
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24950 2408 25006 2417
rect 23388 2372 23440 2378
rect 24950 2343 24952 2352
rect 23388 2314 23440 2320
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 22742 2000 22798 2009
rect 22742 1935 22798 1944
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2314
rect 25056 785 25084 2926
rect 25240 2854 25268 13806
rect 25332 7410 25360 14826
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25424 3058 25452 14282
rect 25516 6322 25544 17002
rect 25608 15609 25636 21830
rect 25700 18873 25728 22374
rect 25686 18864 25742 18873
rect 25686 18799 25742 18808
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25594 15600 25650 15609
rect 25594 15535 25596 15544
rect 25648 15535 25650 15544
rect 25596 15506 25648 15512
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 8022 25636 13194
rect 25596 8016 25648 8022
rect 25596 7958 25648 7964
rect 25700 7818 25728 18634
rect 25792 17746 25820 22510
rect 25884 18358 25912 23530
rect 26054 22808 26110 22817
rect 26054 22743 26110 22752
rect 26068 22094 26096 22743
rect 26068 22066 26372 22094
rect 26054 21176 26110 21185
rect 26054 21111 26110 21120
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 25872 18352 25924 18358
rect 25872 18294 25924 18300
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25780 16176 25832 16182
rect 25780 16118 25832 16124
rect 25792 10062 25820 16118
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25884 11286 25912 13874
rect 25872 11280 25924 11286
rect 25872 11222 25924 11228
rect 25976 10713 26004 20742
rect 26068 20738 26096 21111
rect 26056 20732 26108 20738
rect 26056 20674 26108 20680
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26068 17241 26096 19654
rect 26054 17232 26110 17241
rect 26054 17167 26110 17176
rect 26068 11354 26096 17167
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 25962 10704 26018 10713
rect 25962 10639 26018 10648
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 26252 9178 26280 15506
rect 26344 11694 26372 22066
rect 26424 20732 26476 20738
rect 26424 20674 26476 20680
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26436 9110 26464 20674
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 26620 4146 26648 15302
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 1398 25880 1454 25936
rect 1490 24792 1546 24848
rect 1582 24132 1638 24168
rect 1582 24112 1584 24132
rect 1584 24112 1636 24132
rect 1636 24112 1638 24132
rect 1950 24656 2006 24712
rect 1674 22616 1730 22672
rect 2226 19352 2282 19408
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 3422 23704 3478 23760
rect 3974 25336 4030 25392
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 19760 2834 19816
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3974 23160 4030 23216
rect 4986 25744 5042 25800
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3330 17856 3386 17912
rect 2226 17740 2282 17776
rect 2226 17720 2228 17740
rect 2228 17720 2280 17740
rect 2280 17720 2282 17740
rect 3882 17040 3938 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 4618 23024 4674 23080
rect 4894 20476 4896 20496
rect 4896 20476 4948 20496
rect 4948 20476 4950 20496
rect 4894 20440 4950 20476
rect 4802 19624 4858 19680
rect 4710 19080 4766 19136
rect 4710 17720 4766 17776
rect 5170 26152 5226 26208
rect 5262 22616 5318 22672
rect 5354 20168 5410 20224
rect 5538 22480 5594 22536
rect 5630 20984 5686 21040
rect 5538 20304 5594 20360
rect 5538 18964 5594 19000
rect 5538 18944 5540 18964
rect 5540 18944 5592 18964
rect 5592 18944 5594 18964
rect 5538 18164 5540 18184
rect 5540 18164 5592 18184
rect 5592 18164 5594 18184
rect 5538 18128 5594 18164
rect 4434 15408 4490 15464
rect 4342 13912 4398 13968
rect 6182 23432 6238 23488
rect 6642 26016 6698 26072
rect 6826 23704 6882 23760
rect 6918 23568 6974 23624
rect 6550 19252 6552 19272
rect 6552 19252 6604 19272
rect 6604 19252 6606 19272
rect 6550 19216 6606 19252
rect 7378 21972 7380 21992
rect 7380 21972 7432 21992
rect 7432 21972 7434 21992
rect 7378 21936 7434 21972
rect 7010 21392 7066 21448
rect 7286 19896 7342 19952
rect 7010 17584 7066 17640
rect 6182 15000 6238 15056
rect 7838 24248 7894 24304
rect 7654 20868 7710 20904
rect 7654 20848 7656 20868
rect 7656 20848 7708 20868
rect 7708 20848 7710 20868
rect 7654 20032 7710 20088
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 8206 22072 8262 22128
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7838 20168 7894 20224
rect 8022 20168 8078 20224
rect 8022 19760 8078 19816
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8574 22344 8630 22400
rect 8482 21664 8538 21720
rect 8206 18672 8262 18728
rect 7654 18264 7710 18320
rect 7562 17196 7618 17232
rect 7562 17176 7564 17196
rect 7564 17176 7616 17196
rect 7616 17176 7618 17196
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8390 18808 8446 18864
rect 8298 17756 8300 17776
rect 8300 17756 8352 17776
rect 8352 17756 8354 17776
rect 8298 17720 8354 17756
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8942 24928 8998 24984
rect 8850 22752 8906 22808
rect 9770 23840 9826 23896
rect 9310 21836 9312 21856
rect 9312 21836 9364 21856
rect 9364 21836 9366 21856
rect 9310 21800 9366 21836
rect 8850 19488 8906 19544
rect 8758 17312 8814 17368
rect 8482 16496 8538 16552
rect 8666 16108 8722 16144
rect 8666 16088 8668 16108
rect 8668 16088 8720 16108
rect 8720 16088 8722 16108
rect 8758 15952 8814 16008
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 6550 14320 6606 14376
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 9770 20576 9826 20632
rect 9770 16360 9826 16416
rect 9126 15852 9128 15872
rect 9128 15852 9180 15872
rect 9180 15852 9182 15872
rect 9126 15816 9182 15852
rect 10046 23432 10102 23488
rect 10046 16652 10102 16688
rect 10046 16632 10048 16652
rect 10048 16632 10100 16652
rect 10100 16632 10102 16652
rect 9402 15544 9458 15600
rect 10598 21800 10654 21856
rect 10414 21292 10416 21312
rect 10416 21292 10468 21312
rect 10468 21292 10470 21312
rect 10414 21256 10470 21292
rect 10414 19624 10470 19680
rect 11334 24248 11390 24304
rect 10414 15564 10470 15600
rect 10414 15544 10416 15564
rect 10416 15544 10468 15564
rect 10468 15544 10470 15564
rect 10506 15020 10562 15056
rect 10506 15000 10508 15020
rect 10508 15000 10560 15020
rect 10560 15000 10562 15020
rect 10322 14884 10378 14920
rect 10322 14864 10324 14884
rect 10324 14864 10376 14884
rect 10376 14864 10378 14884
rect 10966 15308 10968 15328
rect 10968 15308 11020 15328
rect 11020 15308 11022 15328
rect 10966 15272 11022 15308
rect 8850 14456 8906 14512
rect 12530 24384 12586 24440
rect 12070 23840 12126 23896
rect 11886 23296 11942 23352
rect 11610 21564 11612 21584
rect 11612 21564 11664 21584
rect 11664 21564 11666 21584
rect 11610 21528 11666 21564
rect 12622 23296 12678 23352
rect 11978 21800 12034 21856
rect 11518 19352 11574 19408
rect 12070 20032 12126 20088
rect 11886 19352 11942 19408
rect 11518 18536 11574 18592
rect 11426 17484 11428 17504
rect 11428 17484 11480 17504
rect 11480 17484 11482 17504
rect 11426 17448 11482 17484
rect 12438 21256 12494 21312
rect 12346 20712 12402 20768
rect 12438 19624 12494 19680
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 13358 23468 13360 23488
rect 13360 23468 13412 23488
rect 13412 23468 13414 23488
rect 13358 23432 13414 23468
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13358 22344 13414 22400
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13818 23840 13874 23896
rect 13542 22616 13598 22672
rect 13634 22072 13690 22128
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13634 21392 13690 21448
rect 13358 20984 13414 21040
rect 12806 20712 12862 20768
rect 12530 18944 12586 19000
rect 12254 17856 12310 17912
rect 12162 16224 12218 16280
rect 12438 16088 12494 16144
rect 12346 15580 12348 15600
rect 12348 15580 12400 15600
rect 12400 15580 12402 15600
rect 12346 15544 12402 15580
rect 12530 15544 12586 15600
rect 12346 15308 12348 15328
rect 12348 15308 12400 15328
rect 12400 15308 12402 15328
rect 10966 13776 11022 13832
rect 12346 15272 12402 15308
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 14462 23024 14518 23080
rect 14094 22344 14150 22400
rect 13818 21256 13874 21312
rect 13358 20748 13360 20768
rect 13360 20748 13412 20768
rect 13412 20748 13414 20768
rect 13358 20712 13414 20748
rect 13542 20712 13598 20768
rect 13174 20596 13230 20632
rect 13174 20576 13176 20596
rect 13176 20576 13228 20596
rect 13228 20576 13230 20596
rect 13358 20576 13414 20632
rect 13358 20168 13414 20224
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13358 15680 13414 15736
rect 14002 20984 14058 21040
rect 14370 22480 14426 22536
rect 14094 20032 14150 20088
rect 14002 17992 14058 18048
rect 13910 16224 13966 16280
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 15382 24112 15438 24168
rect 16394 24928 16450 24984
rect 14462 20848 14518 20904
rect 14370 19352 14426 19408
rect 14094 16632 14150 16688
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 15106 21664 15162 21720
rect 14646 17720 14702 17776
rect 14738 17040 14794 17096
rect 14646 16904 14702 16960
rect 15014 20440 15070 20496
rect 14922 19352 14978 19408
rect 15290 20440 15346 20496
rect 15290 20032 15346 20088
rect 15290 19488 15346 19544
rect 15014 17720 15070 17776
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 15382 16768 15438 16824
rect 15106 11736 15162 11792
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 15566 19508 15622 19544
rect 15566 19488 15568 19508
rect 15568 19488 15620 19508
rect 15620 19488 15622 19508
rect 15934 21800 15990 21856
rect 15842 20748 15844 20768
rect 15844 20748 15896 20768
rect 15896 20748 15898 20768
rect 15842 20712 15898 20748
rect 15934 20304 15990 20360
rect 15658 11636 15660 11656
rect 15660 11636 15712 11656
rect 15712 11636 15714 11656
rect 15658 11600 15714 11636
rect 15658 11192 15714 11248
rect 15474 10240 15530 10296
rect 16486 22480 16542 22536
rect 16302 19896 16358 19952
rect 16302 19760 16358 19816
rect 16486 18264 16542 18320
rect 16854 23840 16910 23896
rect 17038 22344 17094 22400
rect 16854 22072 16910 22128
rect 16946 21664 17002 21720
rect 16854 20576 16910 20632
rect 16854 19352 16910 19408
rect 16762 17992 16818 18048
rect 16118 11348 16174 11384
rect 16118 11328 16120 11348
rect 16120 11328 16172 11348
rect 16172 11328 16174 11348
rect 16854 17448 16910 17504
rect 17498 25744 17554 25800
rect 17314 23024 17370 23080
rect 17222 22752 17278 22808
rect 17222 21800 17278 21856
rect 18970 25880 19026 25936
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 18510 23840 18566 23896
rect 17774 23024 17830 23080
rect 17958 23024 18014 23080
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 19706 26016 19762 26072
rect 20166 26152 20222 26208
rect 20074 25608 20130 25664
rect 18786 22888 18842 22944
rect 17682 21664 17738 21720
rect 17406 20848 17462 20904
rect 17222 20596 17278 20632
rect 17222 20576 17224 20596
rect 17224 20576 17276 20596
rect 17276 20576 17278 20596
rect 17222 19488 17278 19544
rect 17406 19292 17462 19348
rect 17222 19080 17278 19136
rect 16394 13640 16450 13696
rect 17498 18400 17554 18456
rect 17590 10512 17646 10568
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18786 22072 18842 22128
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18142 18808 18198 18864
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17958 17584 18014 17640
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18878 21392 18934 21448
rect 18878 20848 18934 20904
rect 18694 19292 18750 19348
rect 18694 18264 18750 18320
rect 19062 23024 19118 23080
rect 19338 24012 19340 24032
rect 19340 24012 19392 24032
rect 19392 24012 19394 24032
rect 19338 23976 19394 24012
rect 20626 23704 20682 23760
rect 19246 23160 19302 23216
rect 20810 22616 20866 22672
rect 20534 22480 20590 22536
rect 19430 21936 19486 21992
rect 18970 18536 19026 18592
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18510 12416 18566 12472
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18050 10648 18106 10704
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19522 20712 19578 20768
rect 19706 19352 19762 19408
rect 19706 19216 19762 19272
rect 19890 18808 19946 18864
rect 19522 16904 19578 16960
rect 19154 15136 19210 15192
rect 19522 14048 19578 14104
rect 19154 12416 19210 12472
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19890 17992 19946 18048
rect 19522 10648 19578 10704
rect 19430 9444 19486 9480
rect 19430 9424 19432 9444
rect 19432 9424 19484 9444
rect 19484 9424 19486 9444
rect 20166 16360 20222 16416
rect 20074 16088 20130 16144
rect 19798 12416 19854 12472
rect 19706 11056 19762 11112
rect 19890 12280 19946 12336
rect 20442 20576 20498 20632
rect 20626 21528 20682 21584
rect 21178 23296 21234 23352
rect 20810 20304 20866 20360
rect 20350 19252 20352 19272
rect 20352 19252 20404 19272
rect 20404 19252 20406 19272
rect 20350 19216 20406 19252
rect 20534 18400 20590 18456
rect 20442 18284 20498 18320
rect 20442 18264 20444 18284
rect 20444 18264 20496 18284
rect 20496 18264 20498 18284
rect 20258 13640 20314 13696
rect 20166 9424 20222 9480
rect 20718 19760 20774 19816
rect 21914 23432 21970 23488
rect 21730 23024 21786 23080
rect 21546 22344 21602 22400
rect 20810 17584 20866 17640
rect 20810 16632 20866 16688
rect 20810 16088 20866 16144
rect 20994 18300 20996 18320
rect 20996 18300 21048 18320
rect 21048 18300 21050 18320
rect 20994 18264 21050 18300
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20810 12280 20866 12336
rect 21362 19216 21418 19272
rect 21362 17856 21418 17912
rect 22190 22208 22246 22264
rect 22098 20984 22154 21040
rect 21730 20712 21786 20768
rect 21638 17856 21694 17912
rect 21086 12280 21142 12336
rect 20718 10240 20774 10296
rect 21454 11872 21510 11928
rect 22558 19080 22614 19136
rect 22282 17856 22338 17912
rect 22098 14320 22154 14376
rect 21822 12960 21878 13016
rect 21730 12280 21786 12336
rect 22374 15544 22430 15600
rect 22374 15428 22430 15464
rect 22374 15408 22376 15428
rect 22376 15408 22428 15428
rect 22428 15408 22430 15428
rect 22558 18536 22614 18592
rect 23386 25608 23442 25664
rect 23294 25472 23350 25528
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 23386 24384 23442 24440
rect 22834 23568 22890 23624
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23202 20884 23204 20904
rect 23204 20884 23256 20904
rect 23256 20884 23258 20904
rect 23202 20848 23258 20884
rect 23386 21392 23442 21448
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22926 18808 22982 18864
rect 22834 18708 22836 18728
rect 22836 18708 22888 18728
rect 22888 18708 22890 18728
rect 22834 18672 22890 18708
rect 23110 18808 23166 18864
rect 23202 18264 23258 18320
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17720 23442 17776
rect 23110 17448 23166 17504
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22834 16496 22890 16552
rect 22190 12824 22246 12880
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22742 14456 22798 14512
rect 22650 13776 22706 13832
rect 22558 13368 22614 13424
rect 22466 12824 22522 12880
rect 23018 15408 23074 15464
rect 22926 15272 22982 15328
rect 23386 16632 23442 16688
rect 23202 15000 23258 15056
rect 23386 15000 23442 15056
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 21454 8336 21510 8392
rect 21270 7792 21326 7848
rect 22190 11212 22246 11248
rect 22190 11192 22192 11212
rect 22192 11192 22244 11212
rect 22244 11192 22246 11212
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23754 20576 23810 20632
rect 23754 19352 23810 19408
rect 23570 16224 23626 16280
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22650 9560 22706 9616
rect 22190 6296 22246 6352
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23478 9424 23534 9480
rect 25318 26424 25374 26480
rect 24214 26016 24270 26072
rect 25134 25200 25190 25256
rect 25134 24656 25190 24712
rect 25042 24148 25044 24168
rect 25044 24148 25096 24168
rect 25096 24148 25098 24168
rect 25042 24112 25098 24148
rect 24858 23840 24914 23896
rect 24122 18808 24178 18864
rect 24582 22072 24638 22128
rect 24306 18128 24362 18184
rect 24122 15952 24178 16008
rect 23938 14184 23994 14240
rect 24306 15816 24362 15872
rect 24766 20440 24822 20496
rect 24858 19896 24914 19952
rect 24582 19488 24638 19544
rect 24766 19488 24822 19544
rect 24582 17992 24638 18048
rect 23846 9968 23902 10024
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24582 16360 24638 16416
rect 24950 16088 25006 16144
rect 24766 12552 24822 12608
rect 24674 12144 24730 12200
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24858 11328 24914 11384
rect 24766 10920 24822 10976
rect 24582 10104 24638 10160
rect 24858 10512 24914 10568
rect 24858 9288 24914 9344
rect 24674 8880 24730 8936
rect 24858 8508 24860 8528
rect 24860 8508 24912 8528
rect 24912 8508 24914 8528
rect 24858 8472 24914 8508
rect 25134 14864 25190 14920
rect 25134 13932 25190 13968
rect 25134 13912 25136 13932
rect 25136 13912 25188 13932
rect 25188 13912 25190 13932
rect 25042 12300 25098 12336
rect 25042 12280 25044 12300
rect 25044 12280 25096 12300
rect 25096 12280 25098 12300
rect 25134 11636 25136 11656
rect 25136 11636 25188 11656
rect 25188 11636 25190 11656
rect 25134 11600 25190 11636
rect 24950 8064 25006 8120
rect 24766 7656 24822 7712
rect 24674 6432 24730 6488
rect 24858 7248 24914 7304
rect 24858 6860 24914 6896
rect 24858 6840 24860 6860
rect 24860 6840 24912 6860
rect 24912 6840 24914 6860
rect 24858 6024 24914 6080
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24766 5208 24822 5264
rect 24858 4800 24914 4856
rect 24950 4392 25006 4448
rect 25134 3984 25190 4040
rect 24950 3576 25006 3632
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24950 3168 25006 3224
rect 24858 2760 24914 2816
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 22742 1944 22798 2000
rect 22098 1536 22154 1592
rect 22098 1128 22154 1184
rect 25686 18808 25742 18864
rect 25594 15564 25650 15600
rect 25594 15544 25596 15564
rect 25596 15544 25648 15564
rect 25648 15544 25650 15564
rect 26054 22752 26110 22808
rect 26054 21120 26110 21176
rect 26054 17176 26110 17232
rect 25962 10648 26018 10704
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 25313 26482 25379 26485
rect 26200 26482 27000 26512
rect 25313 26480 27000 26482
rect 25313 26424 25318 26480
rect 25374 26424 27000 26480
rect 25313 26422 27000 26424
rect 25313 26419 25379 26422
rect 26200 26392 27000 26422
rect 5165 26210 5231 26213
rect 20161 26210 20227 26213
rect 5165 26208 20227 26210
rect 5165 26152 5170 26208
rect 5226 26152 20166 26208
rect 20222 26152 20227 26208
rect 5165 26150 20227 26152
rect 5165 26147 5231 26150
rect 20161 26147 20227 26150
rect 6637 26074 6703 26077
rect 19701 26074 19767 26077
rect 6637 26072 19767 26074
rect 6637 26016 6642 26072
rect 6698 26016 19706 26072
rect 19762 26016 19767 26072
rect 6637 26014 19767 26016
rect 6637 26011 6703 26014
rect 19701 26011 19767 26014
rect 24209 26074 24275 26077
rect 26200 26074 27000 26104
rect 24209 26072 27000 26074
rect 24209 26016 24214 26072
rect 24270 26016 27000 26072
rect 24209 26014 27000 26016
rect 24209 26011 24275 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 6678 25876 6684 25940
rect 6748 25938 6754 25940
rect 18965 25938 19031 25941
rect 6748 25936 19031 25938
rect 6748 25880 18970 25936
rect 19026 25880 19031 25936
rect 6748 25878 19031 25880
rect 6748 25876 6754 25878
rect 18965 25875 19031 25878
rect 4981 25802 5047 25805
rect 17493 25802 17559 25805
rect 4981 25800 17559 25802
rect 4981 25744 4986 25800
rect 5042 25744 17498 25800
rect 17554 25744 17559 25800
rect 4981 25742 17559 25744
rect 4981 25739 5047 25742
rect 17493 25739 17559 25742
rect 4838 25604 4844 25668
rect 4908 25666 4914 25668
rect 20069 25666 20135 25669
rect 4908 25664 20135 25666
rect 4908 25608 20074 25664
rect 20130 25608 20135 25664
rect 4908 25606 20135 25608
rect 4908 25604 4914 25606
rect 20069 25603 20135 25606
rect 23381 25666 23447 25669
rect 26200 25666 27000 25696
rect 23381 25664 27000 25666
rect 23381 25608 23386 25664
rect 23442 25608 27000 25664
rect 23381 25606 27000 25608
rect 23381 25603 23447 25606
rect 26200 25576 27000 25606
rect 10542 25468 10548 25532
rect 10612 25530 10618 25532
rect 23289 25530 23355 25533
rect 10612 25528 23355 25530
rect 10612 25472 23294 25528
rect 23350 25472 23355 25528
rect 10612 25470 23355 25472
rect 10612 25468 10618 25470
rect 23289 25467 23355 25470
rect 3969 25394 4035 25397
rect 19742 25394 19748 25396
rect 3969 25392 19748 25394
rect 3969 25336 3974 25392
rect 4030 25336 19748 25392
rect 3969 25334 19748 25336
rect 3969 25331 4035 25334
rect 19742 25332 19748 25334
rect 19812 25332 19818 25396
rect 7598 25196 7604 25260
rect 7668 25258 7674 25260
rect 22134 25258 22140 25260
rect 7668 25198 22140 25258
rect 7668 25196 7674 25198
rect 22134 25196 22140 25198
rect 22204 25196 22210 25260
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 9438 25060 9444 25124
rect 9508 25122 9514 25124
rect 9508 25062 17280 25122
rect 9508 25060 9514 25062
rect 8937 24986 9003 24989
rect 16389 24986 16455 24989
rect 8937 24984 16455 24986
rect 8937 24928 8942 24984
rect 8998 24928 16394 24984
rect 16450 24928 16455 24984
rect 8937 24926 16455 24928
rect 17220 24986 17280 25062
rect 17220 24926 22110 24986
rect 8937 24923 9003 24926
rect 16389 24923 16455 24926
rect 0 24850 800 24880
rect 1485 24850 1551 24853
rect 0 24848 1551 24850
rect 0 24792 1490 24848
rect 1546 24792 1551 24848
rect 0 24790 1551 24792
rect 22050 24850 22110 24926
rect 26200 24850 27000 24880
rect 22050 24790 27000 24850
rect 0 24760 800 24790
rect 1485 24787 1551 24790
rect 26200 24760 27000 24790
rect 1945 24714 2011 24717
rect 25129 24714 25195 24717
rect 1945 24712 25195 24714
rect 1945 24656 1950 24712
rect 2006 24656 25134 24712
rect 25190 24656 25195 24712
rect 1945 24654 25195 24656
rect 1945 24651 2011 24654
rect 25129 24651 25195 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 5390 24380 5396 24444
rect 5460 24442 5466 24444
rect 12525 24442 12591 24445
rect 5460 24440 12591 24442
rect 5460 24384 12530 24440
rect 12586 24384 12591 24440
rect 5460 24382 12591 24384
rect 5460 24380 5466 24382
rect 12525 24379 12591 24382
rect 23381 24442 23447 24445
rect 26200 24442 27000 24472
rect 23381 24440 27000 24442
rect 23381 24384 23386 24440
rect 23442 24384 27000 24440
rect 23381 24382 27000 24384
rect 23381 24379 23447 24382
rect 26200 24352 27000 24382
rect 7833 24306 7899 24309
rect 11329 24306 11395 24309
rect 7833 24304 8540 24306
rect 7833 24248 7838 24304
rect 7894 24248 8540 24304
rect 7833 24246 8540 24248
rect 7833 24243 7899 24246
rect 1577 24170 1643 24173
rect 8480 24170 8540 24246
rect 11329 24304 25330 24306
rect 11329 24248 11334 24304
rect 11390 24248 25330 24304
rect 11329 24246 25330 24248
rect 11329 24243 11395 24246
rect 15377 24170 15443 24173
rect 1577 24168 8402 24170
rect 1577 24112 1582 24168
rect 1638 24112 8402 24168
rect 1577 24110 8402 24112
rect 8480 24168 15443 24170
rect 8480 24112 15382 24168
rect 15438 24112 15443 24168
rect 8480 24110 15443 24112
rect 1577 24107 1643 24110
rect 8342 24034 8402 24110
rect 15377 24107 15443 24110
rect 16246 24108 16252 24172
rect 16316 24170 16322 24172
rect 25037 24170 25103 24173
rect 16316 24168 25103 24170
rect 16316 24112 25042 24168
rect 25098 24112 25103 24168
rect 16316 24110 25103 24112
rect 16316 24108 16322 24110
rect 16254 24034 16314 24108
rect 25037 24107 25103 24110
rect 8342 23974 16314 24034
rect 19190 23972 19196 24036
rect 19260 24034 19266 24036
rect 19333 24034 19399 24037
rect 19260 24032 19399 24034
rect 19260 23976 19338 24032
rect 19394 23976 19399 24032
rect 19260 23974 19399 23976
rect 25270 24034 25330 24246
rect 26200 24034 27000 24064
rect 25270 23974 27000 24034
rect 19260 23972 19266 23974
rect 19333 23971 19399 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 9765 23898 9831 23901
rect 12065 23898 12131 23901
rect 9765 23896 12131 23898
rect 9765 23840 9770 23896
rect 9826 23840 12070 23896
rect 12126 23840 12131 23896
rect 9765 23838 12131 23840
rect 9765 23835 9831 23838
rect 12065 23835 12131 23838
rect 13813 23898 13879 23901
rect 14038 23898 14044 23900
rect 13813 23896 14044 23898
rect 13813 23840 13818 23896
rect 13874 23840 14044 23896
rect 13813 23838 14044 23840
rect 13813 23835 13879 23838
rect 14038 23836 14044 23838
rect 14108 23836 14114 23900
rect 16849 23898 16915 23901
rect 17534 23898 17540 23900
rect 16849 23896 17540 23898
rect 16849 23840 16854 23896
rect 16910 23840 17540 23896
rect 16849 23838 17540 23840
rect 16849 23835 16915 23838
rect 17534 23836 17540 23838
rect 17604 23836 17610 23900
rect 18505 23898 18571 23901
rect 24853 23898 24919 23901
rect 18505 23896 24919 23898
rect 18505 23840 18510 23896
rect 18566 23840 24858 23896
rect 24914 23840 24919 23896
rect 18505 23838 24919 23840
rect 18505 23835 18571 23838
rect 24853 23835 24919 23838
rect 0 23762 800 23792
rect 3417 23762 3483 23765
rect 0 23760 3483 23762
rect 0 23704 3422 23760
rect 3478 23704 3483 23760
rect 0 23702 3483 23704
rect 0 23672 800 23702
rect 3417 23699 3483 23702
rect 6821 23762 6887 23765
rect 20621 23762 20687 23765
rect 6821 23760 20687 23762
rect 6821 23704 6826 23760
rect 6882 23704 20626 23760
rect 20682 23704 20687 23760
rect 6821 23702 20687 23704
rect 6821 23699 6887 23702
rect 20621 23699 20687 23702
rect 6913 23626 6979 23629
rect 18638 23626 18644 23628
rect 6913 23624 18644 23626
rect 6913 23568 6918 23624
rect 6974 23568 18644 23624
rect 6913 23566 18644 23568
rect 6913 23563 6979 23566
rect 18638 23564 18644 23566
rect 18708 23564 18714 23628
rect 22829 23626 22895 23629
rect 26200 23626 27000 23656
rect 22829 23624 27000 23626
rect 22829 23568 22834 23624
rect 22890 23568 27000 23624
rect 22829 23566 27000 23568
rect 22829 23563 22895 23566
rect 26200 23536 27000 23566
rect 6177 23490 6243 23493
rect 10041 23490 10107 23493
rect 6177 23488 10107 23490
rect 6177 23432 6182 23488
rect 6238 23432 10046 23488
rect 10102 23432 10107 23488
rect 6177 23430 10107 23432
rect 6177 23427 6243 23430
rect 10041 23427 10107 23430
rect 13353 23490 13419 23493
rect 21909 23490 21975 23493
rect 13353 23488 21975 23490
rect 13353 23432 13358 23488
rect 13414 23432 21914 23488
rect 21970 23432 21975 23488
rect 13353 23430 21975 23432
rect 13353 23427 13419 23430
rect 21909 23427 21975 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 11881 23354 11947 23357
rect 12617 23354 12683 23357
rect 11881 23352 12683 23354
rect 11881 23296 11886 23352
rect 11942 23296 12622 23352
rect 12678 23296 12683 23352
rect 11881 23294 12683 23296
rect 11881 23291 11947 23294
rect 12617 23291 12683 23294
rect 13854 23292 13860 23356
rect 13924 23354 13930 23356
rect 21173 23354 21239 23357
rect 13924 23352 21239 23354
rect 13924 23296 21178 23352
rect 21234 23296 21239 23352
rect 13924 23294 21239 23296
rect 13924 23292 13930 23294
rect 21173 23291 21239 23294
rect 3969 23218 4035 23221
rect 19241 23218 19307 23221
rect 26200 23218 27000 23248
rect 3969 23216 19307 23218
rect 3969 23160 3974 23216
rect 4030 23160 19246 23216
rect 19302 23160 19307 23216
rect 3969 23158 19307 23160
rect 3969 23155 4035 23158
rect 19241 23155 19307 23158
rect 22050 23158 27000 23218
rect 4613 23082 4679 23085
rect 14457 23082 14523 23085
rect 4613 23080 14523 23082
rect 4613 23024 4618 23080
rect 4674 23024 14462 23080
rect 14518 23024 14523 23080
rect 4613 23022 14523 23024
rect 4613 23019 4679 23022
rect 14457 23019 14523 23022
rect 17309 23082 17375 23085
rect 17769 23082 17835 23085
rect 17309 23080 17835 23082
rect 17309 23024 17314 23080
rect 17370 23024 17774 23080
rect 17830 23024 17835 23080
rect 17309 23022 17835 23024
rect 17309 23019 17375 23022
rect 17769 23019 17835 23022
rect 17953 23082 18019 23085
rect 19057 23082 19123 23085
rect 17953 23080 19123 23082
rect 17953 23024 17958 23080
rect 18014 23024 19062 23080
rect 19118 23024 19123 23080
rect 17953 23022 19123 23024
rect 17953 23019 18019 23022
rect 19057 23019 19123 23022
rect 21725 23082 21791 23085
rect 22050 23082 22110 23158
rect 26200 23128 27000 23158
rect 21725 23080 22110 23082
rect 21725 23024 21730 23080
rect 21786 23024 22110 23080
rect 21725 23022 22110 23024
rect 21725 23019 21791 23022
rect 18781 22948 18847 22949
rect 18781 22946 18828 22948
rect 12574 22886 17418 22946
rect 18736 22944 18828 22946
rect 18736 22888 18786 22944
rect 18736 22886 18828 22888
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 8845 22810 8911 22813
rect 12574 22810 12634 22886
rect 8845 22808 12634 22810
rect 8845 22752 8850 22808
rect 8906 22752 12634 22808
rect 8845 22750 12634 22752
rect 8845 22747 8911 22750
rect 12750 22748 12756 22812
rect 12820 22810 12826 22812
rect 17217 22810 17283 22813
rect 12820 22808 17283 22810
rect 12820 22752 17222 22808
rect 17278 22752 17283 22808
rect 12820 22750 17283 22752
rect 12820 22748 12826 22750
rect 17217 22747 17283 22750
rect 0 22674 800 22704
rect 1669 22674 1735 22677
rect 0 22672 1735 22674
rect 0 22616 1674 22672
rect 1730 22616 1735 22672
rect 0 22614 1735 22616
rect 0 22584 800 22614
rect 1669 22611 1735 22614
rect 5257 22674 5323 22677
rect 13537 22674 13603 22677
rect 5257 22672 13603 22674
rect 5257 22616 5262 22672
rect 5318 22616 13542 22672
rect 13598 22616 13603 22672
rect 5257 22614 13603 22616
rect 17358 22674 17418 22886
rect 18781 22884 18828 22886
rect 18892 22884 18898 22948
rect 18781 22883 18847 22884
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 26049 22810 26115 22813
rect 26200 22810 27000 22840
rect 26049 22808 27000 22810
rect 26049 22752 26054 22808
rect 26110 22752 27000 22808
rect 26049 22750 27000 22752
rect 26049 22747 26115 22750
rect 26200 22720 27000 22750
rect 20805 22674 20871 22677
rect 17358 22672 20871 22674
rect 17358 22616 20810 22672
rect 20866 22616 20871 22672
rect 17358 22614 20871 22616
rect 5257 22611 5323 22614
rect 13537 22611 13603 22614
rect 20805 22611 20871 22614
rect 5533 22538 5599 22541
rect 14365 22538 14431 22541
rect 5533 22536 14431 22538
rect 5533 22480 5538 22536
rect 5594 22480 14370 22536
rect 14426 22480 14431 22536
rect 5533 22478 14431 22480
rect 5533 22475 5599 22478
rect 14365 22475 14431 22478
rect 16481 22538 16547 22541
rect 20529 22538 20595 22541
rect 16481 22536 20595 22538
rect 16481 22480 16486 22536
rect 16542 22480 20534 22536
rect 20590 22480 20595 22536
rect 16481 22478 20595 22480
rect 16481 22475 16547 22478
rect 20529 22475 20595 22478
rect 21582 22476 21588 22540
rect 21652 22538 21658 22540
rect 21652 22478 24226 22538
rect 21652 22476 21658 22478
rect 8569 22402 8635 22405
rect 12750 22402 12756 22404
rect 8569 22400 12756 22402
rect 8569 22344 8574 22400
rect 8630 22344 12756 22400
rect 8569 22342 12756 22344
rect 8569 22339 8635 22342
rect 12750 22340 12756 22342
rect 12820 22340 12826 22404
rect 13353 22402 13419 22405
rect 14089 22402 14155 22405
rect 13353 22400 14155 22402
rect 13353 22344 13358 22400
rect 13414 22344 14094 22400
rect 14150 22344 14155 22400
rect 13353 22342 14155 22344
rect 13353 22339 13419 22342
rect 14089 22339 14155 22342
rect 17033 22402 17099 22405
rect 21541 22402 21607 22405
rect 17033 22400 21607 22402
rect 17033 22344 17038 22400
rect 17094 22344 21546 22400
rect 21602 22344 21607 22400
rect 17033 22342 21607 22344
rect 24166 22402 24226 22478
rect 26200 22402 27000 22432
rect 24166 22342 27000 22402
rect 17033 22339 17099 22342
rect 21541 22339 21607 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 26200 22312 27000 22342
rect 22946 22271 23262 22272
rect 22185 22266 22251 22269
rect 13494 22264 22251 22266
rect 13494 22208 22190 22264
rect 22246 22208 22251 22264
rect 13494 22206 22251 22208
rect 8201 22130 8267 22133
rect 13494 22130 13554 22206
rect 22185 22203 22251 22206
rect 8201 22128 13554 22130
rect 8201 22072 8206 22128
rect 8262 22072 13554 22128
rect 8201 22070 13554 22072
rect 13629 22132 13695 22133
rect 13629 22128 13676 22132
rect 13740 22130 13746 22132
rect 16849 22130 16915 22133
rect 18781 22130 18847 22133
rect 13629 22072 13634 22128
rect 8201 22067 8267 22070
rect 13629 22068 13676 22072
rect 13740 22070 13786 22130
rect 16849 22128 18847 22130
rect 16849 22072 16854 22128
rect 16910 22072 18786 22128
rect 18842 22072 18847 22128
rect 16849 22070 18847 22072
rect 13740 22068 13746 22070
rect 13629 22067 13695 22068
rect 16849 22067 16915 22070
rect 18781 22067 18847 22070
rect 21398 22068 21404 22132
rect 21468 22130 21474 22132
rect 24577 22130 24643 22133
rect 21468 22128 24643 22130
rect 21468 22072 24582 22128
rect 24638 22072 24643 22128
rect 21468 22070 24643 22072
rect 21468 22068 21474 22070
rect 24577 22067 24643 22070
rect 7373 21994 7439 21997
rect 19425 21994 19491 21997
rect 7373 21992 19491 21994
rect 7373 21936 7378 21992
rect 7434 21936 19430 21992
rect 19486 21936 19491 21992
rect 7373 21934 19491 21936
rect 7373 21931 7439 21934
rect 19425 21931 19491 21934
rect 22318 21932 22324 21996
rect 22388 21994 22394 21996
rect 26200 21994 27000 22024
rect 22388 21934 27000 21994
rect 22388 21932 22394 21934
rect 26200 21904 27000 21934
rect 9305 21858 9371 21861
rect 9622 21858 9628 21860
rect 9305 21856 9628 21858
rect 9305 21800 9310 21856
rect 9366 21800 9628 21856
rect 9305 21798 9628 21800
rect 9305 21795 9371 21798
rect 9622 21796 9628 21798
rect 9692 21796 9698 21860
rect 10593 21858 10659 21861
rect 11973 21858 12039 21861
rect 15929 21858 15995 21861
rect 17217 21858 17283 21861
rect 10593 21856 17283 21858
rect 10593 21800 10598 21856
rect 10654 21800 11978 21856
rect 12034 21800 15934 21856
rect 15990 21800 17222 21856
rect 17278 21800 17283 21856
rect 10593 21798 17283 21800
rect 10593 21795 10659 21798
rect 11973 21795 12039 21798
rect 15929 21795 15995 21798
rect 17217 21795 17283 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 8477 21722 8543 21725
rect 15101 21722 15167 21725
rect 8477 21720 15167 21722
rect 8477 21664 8482 21720
rect 8538 21664 15106 21720
rect 15162 21664 15167 21720
rect 8477 21662 15167 21664
rect 8477 21659 8543 21662
rect 15101 21659 15167 21662
rect 16941 21722 17007 21725
rect 17677 21722 17743 21725
rect 16941 21720 17743 21722
rect 16941 21664 16946 21720
rect 17002 21664 17682 21720
rect 17738 21664 17743 21720
rect 16941 21662 17743 21664
rect 16941 21659 17007 21662
rect 17677 21659 17743 21662
rect 11605 21586 11671 21589
rect 20621 21586 20687 21589
rect 11605 21584 20687 21586
rect 11605 21528 11610 21584
rect 11666 21528 20626 21584
rect 20682 21528 20687 21584
rect 11605 21526 20687 21528
rect 11605 21523 11671 21526
rect 20621 21523 20687 21526
rect 22502 21524 22508 21588
rect 22572 21586 22578 21588
rect 26200 21586 27000 21616
rect 22572 21526 27000 21586
rect 22572 21524 22578 21526
rect 26200 21496 27000 21526
rect 7005 21450 7071 21453
rect 13629 21450 13695 21453
rect 18873 21450 18939 21453
rect 23381 21450 23447 21453
rect 7005 21448 13695 21450
rect 7005 21392 7010 21448
rect 7066 21392 13634 21448
rect 13690 21392 13695 21448
rect 7005 21390 13695 21392
rect 7005 21387 7071 21390
rect 13629 21387 13695 21390
rect 13862 21448 18939 21450
rect 13862 21392 18878 21448
rect 18934 21392 18939 21448
rect 13862 21390 18939 21392
rect 13862 21317 13922 21390
rect 18873 21387 18939 21390
rect 22050 21448 23447 21450
rect 22050 21392 23386 21448
rect 23442 21392 23447 21448
rect 22050 21390 23447 21392
rect 10409 21314 10475 21317
rect 12433 21314 12499 21317
rect 10409 21312 12499 21314
rect 10409 21256 10414 21312
rect 10470 21256 12438 21312
rect 12494 21256 12499 21312
rect 10409 21254 12499 21256
rect 10409 21251 10475 21254
rect 12433 21251 12499 21254
rect 13813 21312 13922 21317
rect 13813 21256 13818 21312
rect 13874 21256 13922 21312
rect 13813 21254 13922 21256
rect 13813 21251 13879 21254
rect 14222 21252 14228 21316
rect 14292 21314 14298 21316
rect 22050 21314 22110 21390
rect 23381 21387 23447 21390
rect 14292 21254 22110 21314
rect 14292 21252 14298 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 26049 21178 26115 21181
rect 26200 21178 27000 21208
rect 26049 21176 27000 21178
rect 26049 21120 26054 21176
rect 26110 21120 27000 21176
rect 26049 21118 27000 21120
rect 26049 21115 26115 21118
rect 26200 21088 27000 21118
rect 5625 21042 5691 21045
rect 13353 21042 13419 21045
rect 5625 21040 13419 21042
rect 5625 20984 5630 21040
rect 5686 20984 13358 21040
rect 13414 20984 13419 21040
rect 5625 20982 13419 20984
rect 5625 20979 5691 20982
rect 13353 20979 13419 20982
rect 13997 21042 14063 21045
rect 22093 21042 22159 21045
rect 13997 21040 22159 21042
rect 13997 20984 14002 21040
rect 14058 20984 22098 21040
rect 22154 20984 22159 21040
rect 13997 20982 22159 20984
rect 13997 20979 14063 20982
rect 22093 20979 22159 20982
rect 7649 20906 7715 20909
rect 14457 20906 14523 20909
rect 17401 20908 17467 20909
rect 7649 20904 14523 20906
rect 7649 20848 7654 20904
rect 7710 20848 14462 20904
rect 14518 20848 14523 20904
rect 7649 20846 14523 20848
rect 7649 20843 7715 20846
rect 14457 20843 14523 20846
rect 17350 20844 17356 20908
rect 17420 20906 17467 20908
rect 18873 20906 18939 20909
rect 23197 20906 23263 20909
rect 17420 20904 17512 20906
rect 17462 20848 17512 20904
rect 17420 20846 17512 20848
rect 18873 20904 23263 20906
rect 18873 20848 18878 20904
rect 18934 20848 23202 20904
rect 23258 20848 23263 20904
rect 18873 20846 23263 20848
rect 17420 20844 17467 20846
rect 17401 20843 17467 20844
rect 18873 20843 18939 20846
rect 23197 20843 23263 20846
rect 12341 20770 12407 20773
rect 12801 20770 12867 20773
rect 13353 20770 13419 20773
rect 13537 20772 13603 20773
rect 12341 20768 13419 20770
rect 12341 20712 12346 20768
rect 12402 20712 12806 20768
rect 12862 20712 13358 20768
rect 13414 20712 13419 20768
rect 12341 20710 13419 20712
rect 12341 20707 12407 20710
rect 12801 20707 12867 20710
rect 13353 20707 13419 20710
rect 13486 20708 13492 20772
rect 13556 20770 13603 20772
rect 15837 20772 15903 20773
rect 19517 20772 19583 20773
rect 13556 20768 13648 20770
rect 13598 20712 13648 20768
rect 13556 20710 13648 20712
rect 15837 20768 15884 20772
rect 15948 20770 15954 20772
rect 15837 20712 15842 20768
rect 13556 20708 13603 20710
rect 13537 20707 13603 20708
rect 15837 20708 15884 20712
rect 15948 20710 15994 20770
rect 19517 20768 19564 20772
rect 19628 20770 19634 20772
rect 19517 20712 19522 20768
rect 15948 20708 15954 20710
rect 19517 20708 19564 20712
rect 19628 20710 19674 20770
rect 19628 20708 19634 20710
rect 20662 20708 20668 20772
rect 20732 20770 20738 20772
rect 21725 20770 21791 20773
rect 20732 20768 21791 20770
rect 20732 20712 21730 20768
rect 21786 20712 21791 20768
rect 20732 20710 21791 20712
rect 20732 20708 20738 20710
rect 15837 20707 15903 20708
rect 19517 20707 19583 20708
rect 21725 20707 21791 20710
rect 22134 20708 22140 20772
rect 22204 20770 22210 20772
rect 26200 20770 27000 20800
rect 22204 20710 27000 20770
rect 22204 20708 22210 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 26200 20680 27000 20710
rect 17946 20639 18262 20640
rect 9765 20634 9831 20637
rect 13169 20634 13235 20637
rect 9765 20632 13235 20634
rect 9765 20576 9770 20632
rect 9826 20576 13174 20632
rect 13230 20576 13235 20632
rect 9765 20574 13235 20576
rect 9765 20571 9831 20574
rect 13169 20571 13235 20574
rect 13353 20634 13419 20637
rect 16849 20634 16915 20637
rect 17217 20634 17283 20637
rect 13353 20632 17283 20634
rect 13353 20576 13358 20632
rect 13414 20576 16854 20632
rect 16910 20576 17222 20632
rect 17278 20576 17283 20632
rect 13353 20574 17283 20576
rect 13353 20571 13419 20574
rect 16849 20571 16915 20574
rect 17217 20571 17283 20574
rect 20437 20634 20503 20637
rect 23749 20634 23815 20637
rect 20437 20632 23815 20634
rect 20437 20576 20442 20632
rect 20498 20576 23754 20632
rect 23810 20576 23815 20632
rect 20437 20574 23815 20576
rect 20437 20571 20503 20574
rect 23749 20571 23815 20574
rect 4889 20498 4955 20501
rect 15009 20498 15075 20501
rect 4889 20496 15075 20498
rect 4889 20440 4894 20496
rect 4950 20440 15014 20496
rect 15070 20440 15075 20496
rect 4889 20438 15075 20440
rect 4889 20435 4955 20438
rect 15009 20435 15075 20438
rect 15285 20498 15351 20501
rect 24761 20498 24827 20501
rect 15285 20496 24827 20498
rect 15285 20440 15290 20496
rect 15346 20440 24766 20496
rect 24822 20440 24827 20496
rect 15285 20438 24827 20440
rect 15285 20435 15351 20438
rect 24761 20435 24827 20438
rect 5533 20362 5599 20365
rect 15929 20362 15995 20365
rect 5533 20360 15995 20362
rect 5533 20304 5538 20360
rect 5594 20304 15934 20360
rect 15990 20304 15995 20360
rect 5533 20302 15995 20304
rect 5533 20299 5599 20302
rect 15929 20299 15995 20302
rect 20110 20300 20116 20364
rect 20180 20362 20186 20364
rect 20805 20362 20871 20365
rect 26200 20362 27000 20392
rect 20180 20360 20871 20362
rect 20180 20304 20810 20360
rect 20866 20304 20871 20360
rect 20180 20302 20871 20304
rect 20180 20300 20186 20302
rect 20805 20299 20871 20302
rect 22050 20302 27000 20362
rect 5349 20226 5415 20229
rect 7833 20226 7899 20229
rect 5349 20224 7899 20226
rect 5349 20168 5354 20224
rect 5410 20168 7838 20224
rect 7894 20168 7899 20224
rect 5349 20166 7899 20168
rect 5349 20163 5415 20166
rect 7833 20163 7899 20166
rect 8017 20226 8083 20229
rect 13353 20226 13419 20229
rect 14038 20226 14044 20228
rect 8017 20224 12818 20226
rect 8017 20168 8022 20224
rect 8078 20168 12818 20224
rect 8017 20166 12818 20168
rect 8017 20163 8083 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 7649 20090 7715 20093
rect 12065 20090 12131 20093
rect 7649 20088 12131 20090
rect 7649 20032 7654 20088
rect 7710 20032 12070 20088
rect 12126 20032 12131 20088
rect 7649 20030 12131 20032
rect 7649 20027 7715 20030
rect 12065 20027 12131 20030
rect 7281 19954 7347 19957
rect 12566 19954 12572 19956
rect 7281 19952 12572 19954
rect 7281 19896 7286 19952
rect 7342 19896 12572 19952
rect 7281 19894 12572 19896
rect 7281 19891 7347 19894
rect 12566 19892 12572 19894
rect 12636 19892 12642 19956
rect 12758 19954 12818 20166
rect 13353 20224 14044 20226
rect 13353 20168 13358 20224
rect 13414 20168 14044 20224
rect 13353 20166 14044 20168
rect 13353 20163 13419 20166
rect 14038 20164 14044 20166
rect 14108 20164 14114 20228
rect 15142 20164 15148 20228
rect 15212 20226 15218 20228
rect 22050 20226 22110 20302
rect 26200 20272 27000 20302
rect 15212 20166 22110 20226
rect 15212 20164 15218 20166
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 14089 20090 14155 20093
rect 15285 20090 15351 20093
rect 14089 20088 15351 20090
rect 14089 20032 14094 20088
rect 14150 20032 15290 20088
rect 15346 20032 15351 20088
rect 14089 20030 15351 20032
rect 14089 20027 14155 20030
rect 15285 20027 15351 20030
rect 16297 19954 16363 19957
rect 12758 19952 16363 19954
rect 12758 19896 16302 19952
rect 16358 19896 16363 19952
rect 12758 19894 16363 19896
rect 16297 19891 16363 19894
rect 17166 19892 17172 19956
rect 17236 19954 17242 19956
rect 18454 19954 18460 19956
rect 17236 19894 18460 19954
rect 17236 19892 17242 19894
rect 18454 19892 18460 19894
rect 18524 19892 18530 19956
rect 24853 19954 24919 19957
rect 26200 19954 27000 19984
rect 24853 19952 27000 19954
rect 24853 19896 24858 19952
rect 24914 19896 27000 19952
rect 24853 19894 27000 19896
rect 24853 19891 24919 19894
rect 26200 19864 27000 19894
rect 2773 19818 2839 19821
rect 8017 19818 8083 19821
rect 16297 19818 16363 19821
rect 20713 19818 20779 19821
rect 2773 19816 8083 19818
rect 2773 19760 2778 19816
rect 2834 19760 8022 19816
rect 8078 19760 8083 19816
rect 2773 19758 8083 19760
rect 2773 19755 2839 19758
rect 8017 19755 8083 19758
rect 8342 19816 16363 19818
rect 8342 19760 16302 19816
rect 16358 19760 16363 19816
rect 8342 19758 16363 19760
rect 4797 19682 4863 19685
rect 5390 19682 5396 19684
rect 4797 19680 5396 19682
rect 4797 19624 4802 19680
rect 4858 19624 5396 19680
rect 4797 19622 5396 19624
rect 4797 19619 4863 19622
rect 5390 19620 5396 19622
rect 5460 19620 5466 19684
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 2221 19410 2287 19413
rect 8342 19410 8402 19758
rect 16297 19755 16363 19758
rect 16438 19816 20779 19818
rect 16438 19760 20718 19816
rect 20774 19760 20779 19816
rect 16438 19758 20779 19760
rect 10409 19682 10475 19685
rect 12433 19682 12499 19685
rect 10409 19680 12499 19682
rect 10409 19624 10414 19680
rect 10470 19624 12438 19680
rect 12494 19624 12499 19680
rect 10409 19622 12499 19624
rect 10409 19619 10475 19622
rect 12433 19619 12499 19622
rect 12566 19620 12572 19684
rect 12636 19682 12642 19684
rect 16438 19682 16498 19758
rect 20713 19755 20779 19758
rect 12636 19622 16498 19682
rect 12636 19620 12642 19622
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 8845 19546 8911 19549
rect 15285 19546 15351 19549
rect 8845 19544 15351 19546
rect 8845 19488 8850 19544
rect 8906 19488 15290 19544
rect 15346 19488 15351 19544
rect 8845 19486 15351 19488
rect 8845 19483 8911 19486
rect 15285 19483 15351 19486
rect 15561 19546 15627 19549
rect 17217 19546 17283 19549
rect 15561 19544 17283 19546
rect 15561 19488 15566 19544
rect 15622 19488 17222 19544
rect 17278 19488 17283 19544
rect 15561 19486 17283 19488
rect 15561 19483 15627 19486
rect 17217 19483 17283 19486
rect 18454 19484 18460 19548
rect 18524 19546 18530 19548
rect 24577 19546 24643 19549
rect 18524 19544 24643 19546
rect 18524 19488 24582 19544
rect 24638 19488 24643 19544
rect 18524 19486 24643 19488
rect 18524 19484 18530 19486
rect 24577 19483 24643 19486
rect 24761 19546 24827 19549
rect 26200 19546 27000 19576
rect 24761 19544 27000 19546
rect 24761 19488 24766 19544
rect 24822 19488 27000 19544
rect 24761 19486 27000 19488
rect 24761 19483 24827 19486
rect 26200 19456 27000 19486
rect 2221 19408 8402 19410
rect 2221 19352 2226 19408
rect 2282 19352 8402 19408
rect 2221 19350 8402 19352
rect 11513 19410 11579 19413
rect 11881 19410 11947 19413
rect 14222 19410 14228 19412
rect 11513 19408 14228 19410
rect 11513 19352 11518 19408
rect 11574 19352 11886 19408
rect 11942 19352 14228 19408
rect 11513 19350 14228 19352
rect 2221 19347 2287 19350
rect 11513 19347 11579 19350
rect 11881 19347 11947 19350
rect 14222 19348 14228 19350
rect 14292 19348 14298 19412
rect 14365 19410 14431 19413
rect 14917 19410 14983 19413
rect 16849 19410 16915 19413
rect 14365 19408 16915 19410
rect 14365 19352 14370 19408
rect 14426 19352 14922 19408
rect 14978 19352 16854 19408
rect 16910 19352 16915 19408
rect 14365 19350 16915 19352
rect 14365 19347 14431 19350
rect 14917 19347 14983 19350
rect 16849 19347 16915 19350
rect 17166 19348 17172 19412
rect 17236 19348 17242 19412
rect 17350 19348 17356 19412
rect 17420 19353 17426 19412
rect 17420 19348 17467 19353
rect 17534 19348 17540 19412
rect 17604 19348 17610 19412
rect 18822 19410 18828 19412
rect 18646 19350 18828 19410
rect 18646 19348 18755 19350
rect 18822 19348 18828 19350
rect 18892 19348 18898 19412
rect 19374 19348 19380 19412
rect 19444 19410 19450 19412
rect 19701 19410 19767 19413
rect 23749 19410 23815 19413
rect 19444 19408 19767 19410
rect 19444 19352 19706 19408
rect 19762 19352 19767 19408
rect 19444 19350 19767 19352
rect 19444 19348 19450 19350
rect 6545 19274 6611 19277
rect 6678 19274 6684 19276
rect 6545 19272 6684 19274
rect 6545 19216 6550 19272
rect 6606 19216 6684 19272
rect 6545 19214 6684 19216
rect 6545 19211 6611 19214
rect 6678 19212 6684 19214
rect 6748 19212 6754 19276
rect 17174 19274 17234 19348
rect 17358 19292 17406 19348
rect 17462 19292 17467 19348
rect 17358 19290 17467 19292
rect 17401 19287 17467 19290
rect 12390 19214 17234 19274
rect 17542 19274 17602 19348
rect 18646 19292 18694 19348
rect 18750 19292 18755 19348
rect 19701 19347 19767 19350
rect 23614 19408 23815 19410
rect 23614 19352 23754 19408
rect 23810 19352 23815 19408
rect 23614 19350 23815 19352
rect 18646 19290 18755 19292
rect 18689 19287 18755 19290
rect 19701 19274 19767 19277
rect 20345 19274 20411 19277
rect 17542 19214 17970 19274
rect 4705 19138 4771 19141
rect 12390 19138 12450 19214
rect 4705 19136 12450 19138
rect 4705 19080 4710 19136
rect 4766 19080 12450 19136
rect 4705 19078 12450 19080
rect 17217 19138 17283 19141
rect 17718 19138 17724 19140
rect 17217 19136 17724 19138
rect 17217 19080 17222 19136
rect 17278 19080 17724 19136
rect 17217 19078 17724 19080
rect 4705 19075 4771 19078
rect 17217 19075 17283 19078
rect 17718 19076 17724 19078
rect 17788 19076 17794 19140
rect 17910 19138 17970 19214
rect 19701 19272 20411 19274
rect 19701 19216 19706 19272
rect 19762 19216 20350 19272
rect 20406 19216 20411 19272
rect 19701 19214 20411 19216
rect 19701 19211 19767 19214
rect 20345 19211 20411 19214
rect 21357 19274 21423 19277
rect 23614 19274 23674 19350
rect 23749 19347 23815 19350
rect 21357 19272 23674 19274
rect 21357 19216 21362 19272
rect 21418 19216 23674 19272
rect 21357 19214 23674 19216
rect 21357 19211 21423 19214
rect 22553 19138 22619 19141
rect 26200 19138 27000 19168
rect 17910 19136 22619 19138
rect 17910 19080 22558 19136
rect 22614 19080 22619 19136
rect 17910 19078 22619 19080
rect 22553 19075 22619 19078
rect 23614 19078 27000 19138
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 5533 19002 5599 19005
rect 12525 19002 12591 19005
rect 5533 19000 12591 19002
rect 5533 18944 5538 19000
rect 5594 18944 12530 19000
rect 12586 18944 12591 19000
rect 5533 18942 12591 18944
rect 5533 18939 5599 18942
rect 12525 18939 12591 18942
rect 17174 18942 22110 19002
rect 8385 18866 8451 18869
rect 17174 18866 17234 18942
rect 8385 18864 17234 18866
rect 8385 18808 8390 18864
rect 8446 18808 17234 18864
rect 8385 18806 17234 18808
rect 18137 18866 18203 18869
rect 19885 18866 19951 18869
rect 18137 18864 19951 18866
rect 18137 18808 18142 18864
rect 18198 18808 19890 18864
rect 19946 18808 19951 18864
rect 18137 18806 19951 18808
rect 22050 18866 22110 18942
rect 22921 18866 22987 18869
rect 22050 18864 22987 18866
rect 22050 18808 22926 18864
rect 22982 18808 22987 18864
rect 22050 18806 22987 18808
rect 8385 18803 8451 18806
rect 18137 18803 18203 18806
rect 19885 18803 19951 18806
rect 22921 18803 22987 18806
rect 23105 18866 23171 18869
rect 23614 18866 23674 19078
rect 26200 19048 27000 19078
rect 23105 18864 23674 18866
rect 23105 18808 23110 18864
rect 23166 18808 23674 18864
rect 23105 18806 23674 18808
rect 24117 18866 24183 18869
rect 25681 18866 25747 18869
rect 24117 18864 25747 18866
rect 24117 18808 24122 18864
rect 24178 18808 25686 18864
rect 25742 18808 25747 18864
rect 24117 18806 25747 18808
rect 23105 18803 23171 18806
rect 24117 18803 24183 18806
rect 25681 18803 25747 18806
rect 8201 18730 8267 18733
rect 22829 18730 22895 18733
rect 26200 18730 27000 18760
rect 8201 18728 22895 18730
rect 8201 18672 8206 18728
rect 8262 18672 22834 18728
rect 22890 18672 22895 18728
rect 8201 18670 22895 18672
rect 8201 18667 8267 18670
rect 22829 18667 22895 18670
rect 23016 18670 27000 18730
rect 11513 18594 11579 18597
rect 18965 18594 19031 18597
rect 22553 18594 22619 18597
rect 11513 18592 17786 18594
rect 11513 18536 11518 18592
rect 11574 18536 17786 18592
rect 11513 18534 17786 18536
rect 11513 18531 11579 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 15510 18396 15516 18460
rect 15580 18458 15586 18460
rect 17493 18458 17559 18461
rect 15580 18456 17559 18458
rect 15580 18400 17498 18456
rect 17554 18400 17559 18456
rect 15580 18398 17559 18400
rect 15580 18396 15586 18398
rect 17493 18395 17559 18398
rect 7649 18322 7715 18325
rect 16481 18322 16547 18325
rect 7649 18320 16547 18322
rect 7649 18264 7654 18320
rect 7710 18264 16486 18320
rect 16542 18264 16547 18320
rect 7649 18262 16547 18264
rect 17726 18322 17786 18534
rect 18965 18592 22619 18594
rect 18965 18536 18970 18592
rect 19026 18536 22558 18592
rect 22614 18536 22619 18592
rect 18965 18534 22619 18536
rect 18965 18531 19031 18534
rect 22553 18531 22619 18534
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 20529 18458 20595 18461
rect 23016 18458 23076 18670
rect 26200 18640 27000 18670
rect 20529 18456 23076 18458
rect 20529 18400 20534 18456
rect 20590 18400 23076 18456
rect 20529 18398 23076 18400
rect 20529 18395 20595 18398
rect 18689 18322 18755 18325
rect 17726 18320 18755 18322
rect 17726 18264 18694 18320
rect 18750 18264 18755 18320
rect 17726 18262 18755 18264
rect 7649 18259 7715 18262
rect 16481 18259 16547 18262
rect 18689 18259 18755 18262
rect 20437 18322 20503 18325
rect 20989 18322 21055 18325
rect 20437 18320 21055 18322
rect 20437 18264 20442 18320
rect 20498 18264 20994 18320
rect 21050 18264 21055 18320
rect 20437 18262 21055 18264
rect 20437 18259 20503 18262
rect 20989 18259 21055 18262
rect 23197 18322 23263 18325
rect 26200 18322 27000 18352
rect 23197 18320 27000 18322
rect 23197 18264 23202 18320
rect 23258 18264 27000 18320
rect 23197 18262 27000 18264
rect 23197 18259 23263 18262
rect 26200 18232 27000 18262
rect 5533 18186 5599 18189
rect 24301 18186 24367 18189
rect 5533 18184 24367 18186
rect 5533 18128 5538 18184
rect 5594 18128 24306 18184
rect 24362 18128 24367 18184
rect 5533 18126 24367 18128
rect 5533 18123 5599 18126
rect 24301 18123 24367 18126
rect 13997 18050 14063 18053
rect 16757 18050 16823 18053
rect 13997 18048 16823 18050
rect 13997 17992 14002 18048
rect 14058 17992 16762 18048
rect 16818 17992 16823 18048
rect 13997 17990 16823 17992
rect 13997 17987 14063 17990
rect 16757 17987 16823 17990
rect 19742 17988 19748 18052
rect 19812 18050 19818 18052
rect 19885 18050 19951 18053
rect 19812 18048 19951 18050
rect 19812 17992 19890 18048
rect 19946 17992 19951 18048
rect 19812 17990 19951 17992
rect 19812 17988 19818 17990
rect 19885 17987 19951 17990
rect 23422 17988 23428 18052
rect 23492 18050 23498 18052
rect 24577 18050 24643 18053
rect 23492 18048 24643 18050
rect 23492 17992 24582 18048
rect 24638 17992 24643 18048
rect 23492 17990 24643 17992
rect 23492 17988 23498 17990
rect 24577 17987 24643 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 3325 17914 3391 17917
rect 12249 17914 12315 17917
rect 21357 17914 21423 17917
rect 3325 17912 12315 17914
rect 3325 17856 3330 17912
rect 3386 17856 12254 17912
rect 12310 17856 12315 17912
rect 3325 17854 12315 17856
rect 3325 17851 3391 17854
rect 12249 17851 12315 17854
rect 14782 17912 21423 17914
rect 14782 17856 21362 17912
rect 21418 17856 21423 17912
rect 14782 17854 21423 17856
rect 2221 17778 2287 17781
rect 4705 17778 4771 17781
rect 4838 17778 4844 17780
rect 2221 17776 2790 17778
rect 2221 17720 2226 17776
rect 2282 17720 2790 17776
rect 2221 17718 2790 17720
rect 2221 17715 2287 17718
rect 2730 17370 2790 17718
rect 4705 17776 4844 17778
rect 4705 17720 4710 17776
rect 4766 17720 4844 17776
rect 4705 17718 4844 17720
rect 4705 17715 4771 17718
rect 4838 17716 4844 17718
rect 4908 17716 4914 17780
rect 8293 17778 8359 17781
rect 14641 17778 14707 17781
rect 8293 17776 14707 17778
rect 8293 17720 8298 17776
rect 8354 17720 14646 17776
rect 14702 17720 14707 17776
rect 8293 17718 14707 17720
rect 8293 17715 8359 17718
rect 14641 17715 14707 17718
rect 7005 17642 7071 17645
rect 14782 17642 14842 17854
rect 21357 17851 21423 17854
rect 21633 17914 21699 17917
rect 22277 17914 22343 17917
rect 26200 17914 27000 17944
rect 21633 17912 22343 17914
rect 21633 17856 21638 17912
rect 21694 17856 22282 17912
rect 22338 17856 22343 17912
rect 21633 17854 22343 17856
rect 21633 17851 21699 17854
rect 22277 17851 22343 17854
rect 24166 17854 27000 17914
rect 15009 17778 15075 17781
rect 23381 17778 23447 17781
rect 15009 17776 23447 17778
rect 15009 17720 15014 17776
rect 15070 17720 23386 17776
rect 23442 17720 23447 17776
rect 15009 17718 23447 17720
rect 15009 17715 15075 17718
rect 23381 17715 23447 17718
rect 17953 17642 18019 17645
rect 7005 17640 14842 17642
rect 7005 17584 7010 17640
rect 7066 17584 14842 17640
rect 7005 17582 14842 17584
rect 17174 17640 18019 17642
rect 17174 17584 17958 17640
rect 18014 17584 18019 17640
rect 17174 17582 18019 17584
rect 7005 17579 7071 17582
rect 11421 17506 11487 17509
rect 16849 17506 16915 17509
rect 11421 17504 16915 17506
rect 11421 17448 11426 17504
rect 11482 17448 16854 17504
rect 16910 17448 16915 17504
rect 11421 17446 16915 17448
rect 11421 17443 11487 17446
rect 16849 17443 16915 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 8753 17370 8819 17373
rect 17174 17370 17234 17582
rect 17953 17579 18019 17582
rect 20805 17642 20871 17645
rect 24166 17642 24226 17854
rect 26200 17824 27000 17854
rect 20805 17640 24226 17642
rect 20805 17584 20810 17640
rect 20866 17584 24226 17640
rect 20805 17582 24226 17584
rect 20805 17579 20871 17582
rect 23105 17506 23171 17509
rect 26200 17506 27000 17536
rect 23105 17504 27000 17506
rect 23105 17448 23110 17504
rect 23166 17448 27000 17504
rect 23105 17446 27000 17448
rect 23105 17443 23171 17446
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 26200 17416 27000 17446
rect 17946 17375 18262 17376
rect 2730 17310 7850 17370
rect 7557 17236 7623 17237
rect 7557 17234 7604 17236
rect 7512 17232 7604 17234
rect 7512 17176 7562 17232
rect 7512 17174 7604 17176
rect 7557 17172 7604 17174
rect 7668 17172 7674 17236
rect 7790 17234 7850 17310
rect 8753 17368 17234 17370
rect 8753 17312 8758 17368
rect 8814 17312 17234 17368
rect 8753 17310 17234 17312
rect 8753 17307 8819 17310
rect 26049 17234 26115 17237
rect 7790 17232 26115 17234
rect 7790 17176 26054 17232
rect 26110 17176 26115 17232
rect 7790 17174 26115 17176
rect 7557 17171 7623 17172
rect 26049 17171 26115 17174
rect 3877 17098 3943 17101
rect 14733 17098 14799 17101
rect 3877 17096 14799 17098
rect 3877 17040 3882 17096
rect 3938 17040 14738 17096
rect 14794 17040 14799 17096
rect 3877 17038 14799 17040
rect 3877 17035 3943 17038
rect 14733 17035 14799 17038
rect 21950 17036 21956 17100
rect 22020 17098 22026 17100
rect 26200 17098 27000 17128
rect 22020 17038 27000 17098
rect 22020 17036 22026 17038
rect 26200 17008 27000 17038
rect 14641 16962 14707 16965
rect 19517 16962 19583 16965
rect 14641 16960 19583 16962
rect 14641 16904 14646 16960
rect 14702 16904 19522 16960
rect 19578 16904 19583 16960
rect 14641 16902 19583 16904
rect 14641 16899 14707 16902
rect 19517 16899 19583 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 15377 16826 15443 16829
rect 19190 16826 19196 16828
rect 15377 16824 19196 16826
rect 15377 16768 15382 16824
rect 15438 16768 19196 16824
rect 15377 16766 19196 16768
rect 15377 16763 15443 16766
rect 19190 16764 19196 16766
rect 19260 16764 19266 16828
rect 10041 16690 10107 16693
rect 13854 16690 13860 16692
rect 10041 16688 13860 16690
rect 10041 16632 10046 16688
rect 10102 16632 13860 16688
rect 10041 16630 13860 16632
rect 10041 16627 10107 16630
rect 13854 16628 13860 16630
rect 13924 16628 13930 16692
rect 14089 16690 14155 16693
rect 20805 16690 20871 16693
rect 14089 16688 20871 16690
rect 14089 16632 14094 16688
rect 14150 16632 20810 16688
rect 20866 16632 20871 16688
rect 14089 16630 20871 16632
rect 14089 16627 14155 16630
rect 20805 16627 20871 16630
rect 23381 16690 23447 16693
rect 26200 16690 27000 16720
rect 23381 16688 27000 16690
rect 23381 16632 23386 16688
rect 23442 16632 27000 16688
rect 23381 16630 27000 16632
rect 23381 16627 23447 16630
rect 26200 16600 27000 16630
rect 8477 16554 8543 16557
rect 22829 16554 22895 16557
rect 8477 16552 22895 16554
rect 8477 16496 8482 16552
rect 8538 16496 22834 16552
rect 22890 16496 22895 16552
rect 8477 16494 22895 16496
rect 8477 16491 8543 16494
rect 22829 16491 22895 16494
rect 9765 16418 9831 16421
rect 20161 16418 20227 16421
rect 24577 16418 24643 16421
rect 9765 16416 17234 16418
rect 9765 16360 9770 16416
rect 9826 16360 17234 16416
rect 9765 16358 17234 16360
rect 9765 16355 9831 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 12157 16282 12223 16285
rect 13905 16282 13971 16285
rect 12157 16280 13971 16282
rect 12157 16224 12162 16280
rect 12218 16224 13910 16280
rect 13966 16224 13971 16280
rect 12157 16222 13971 16224
rect 12157 16219 12223 16222
rect 13905 16219 13971 16222
rect 8661 16146 8727 16149
rect 12433 16146 12499 16149
rect 15142 16146 15148 16148
rect 8661 16144 12499 16146
rect 8661 16088 8666 16144
rect 8722 16088 12438 16144
rect 12494 16088 12499 16144
rect 8661 16086 12499 16088
rect 8661 16083 8727 16086
rect 12433 16083 12499 16086
rect 12574 16086 15148 16146
rect 8753 16010 8819 16013
rect 12574 16010 12634 16086
rect 15142 16084 15148 16086
rect 15212 16084 15218 16148
rect 17174 16146 17234 16358
rect 20161 16416 24643 16418
rect 20161 16360 20166 16416
rect 20222 16360 24582 16416
rect 24638 16360 24643 16416
rect 20161 16358 24643 16360
rect 20161 16355 20227 16358
rect 24577 16355 24643 16358
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 23565 16282 23631 16285
rect 26200 16282 27000 16312
rect 23565 16280 27000 16282
rect 23565 16224 23570 16280
rect 23626 16224 27000 16280
rect 23565 16222 27000 16224
rect 23565 16219 23631 16222
rect 26200 16192 27000 16222
rect 20069 16146 20135 16149
rect 17174 16144 20135 16146
rect 17174 16088 20074 16144
rect 20130 16088 20135 16144
rect 17174 16086 20135 16088
rect 20069 16083 20135 16086
rect 20805 16146 20871 16149
rect 24945 16146 25011 16149
rect 20805 16144 25011 16146
rect 20805 16088 20810 16144
rect 20866 16088 24950 16144
rect 25006 16088 25011 16144
rect 20805 16086 25011 16088
rect 20805 16083 20871 16086
rect 24945 16083 25011 16086
rect 8753 16008 12634 16010
rect 8753 15952 8758 16008
rect 8814 15952 12634 16008
rect 8753 15950 12634 15952
rect 12712 15950 13554 16010
rect 8753 15947 8819 15950
rect 9121 15874 9187 15877
rect 12712 15874 12772 15950
rect 9121 15872 12772 15874
rect 9121 15816 9126 15872
rect 9182 15816 12772 15872
rect 9121 15814 12772 15816
rect 13494 15874 13554 15950
rect 18638 15948 18644 16012
rect 18708 16010 18714 16012
rect 24117 16010 24183 16013
rect 18708 16008 24183 16010
rect 18708 15952 24122 16008
rect 24178 15952 24183 16008
rect 18708 15950 24183 15952
rect 18708 15948 18714 15950
rect 24117 15947 24183 15950
rect 24301 15874 24367 15877
rect 26200 15874 27000 15904
rect 13494 15814 22754 15874
rect 9121 15811 9187 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 13353 15738 13419 15741
rect 21398 15738 21404 15740
rect 13353 15736 21404 15738
rect 13353 15680 13358 15736
rect 13414 15680 21404 15736
rect 13353 15678 21404 15680
rect 13353 15675 13419 15678
rect 21398 15676 21404 15678
rect 21468 15676 21474 15740
rect 9397 15604 9463 15605
rect 9397 15602 9444 15604
rect 9352 15600 9444 15602
rect 9352 15544 9402 15600
rect 9352 15542 9444 15544
rect 9397 15540 9444 15542
rect 9508 15540 9514 15604
rect 10409 15602 10475 15605
rect 12341 15602 12407 15605
rect 10409 15600 12407 15602
rect 10409 15544 10414 15600
rect 10470 15544 12346 15600
rect 12402 15544 12407 15600
rect 10409 15542 12407 15544
rect 9397 15539 9463 15540
rect 10409 15539 10475 15542
rect 12341 15539 12407 15542
rect 12525 15602 12591 15605
rect 22369 15602 22435 15605
rect 12525 15600 22435 15602
rect 12525 15544 12530 15600
rect 12586 15544 22374 15600
rect 22430 15544 22435 15600
rect 12525 15542 22435 15544
rect 22694 15602 22754 15814
rect 24301 15872 27000 15874
rect 24301 15816 24306 15872
rect 24362 15816 27000 15872
rect 24301 15814 27000 15816
rect 24301 15811 24367 15814
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 25589 15602 25655 15605
rect 22694 15600 25655 15602
rect 22694 15544 25594 15600
rect 25650 15544 25655 15600
rect 22694 15542 25655 15544
rect 12525 15539 12591 15542
rect 22369 15539 22435 15542
rect 25589 15539 25655 15542
rect 4429 15466 4495 15469
rect 22369 15466 22435 15469
rect 4429 15464 22435 15466
rect 4429 15408 4434 15464
rect 4490 15408 22374 15464
rect 22430 15408 22435 15464
rect 4429 15406 22435 15408
rect 4429 15403 4495 15406
rect 22369 15403 22435 15406
rect 23013 15466 23079 15469
rect 26200 15466 27000 15496
rect 23013 15464 27000 15466
rect 23013 15408 23018 15464
rect 23074 15408 27000 15464
rect 23013 15406 27000 15408
rect 23013 15403 23079 15406
rect 26200 15376 27000 15406
rect 10961 15330 11027 15333
rect 12341 15330 12407 15333
rect 10961 15328 12407 15330
rect 10961 15272 10966 15328
rect 11022 15272 12346 15328
rect 12402 15272 12407 15328
rect 10961 15270 12407 15272
rect 10961 15267 11027 15270
rect 12341 15267 12407 15270
rect 22686 15268 22692 15332
rect 22756 15330 22762 15332
rect 22921 15330 22987 15333
rect 22756 15328 22987 15330
rect 22756 15272 22926 15328
rect 22982 15272 22987 15328
rect 22756 15270 22987 15272
rect 22756 15268 22762 15270
rect 22921 15267 22987 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 19149 15194 19215 15197
rect 22134 15194 22140 15196
rect 10182 15134 12450 15194
rect 6177 15058 6243 15061
rect 10182 15058 10242 15134
rect 10501 15060 10567 15061
rect 10501 15058 10548 15060
rect 6177 15056 10242 15058
rect 6177 15000 6182 15056
rect 6238 15000 10242 15056
rect 6177 14998 10242 15000
rect 10456 15056 10548 15058
rect 10456 15000 10506 15056
rect 10456 14998 10548 15000
rect 6177 14995 6243 14998
rect 10501 14996 10548 14998
rect 10612 14996 10618 15060
rect 12390 15058 12450 15134
rect 19149 15192 22140 15194
rect 19149 15136 19154 15192
rect 19210 15136 22140 15192
rect 19149 15134 22140 15136
rect 19149 15131 19215 15134
rect 22134 15132 22140 15134
rect 22204 15132 22210 15196
rect 12390 14998 22110 15058
rect 10501 14995 10567 14996
rect 10317 14922 10383 14925
rect 19374 14922 19380 14924
rect 10317 14920 19380 14922
rect 10317 14864 10322 14920
rect 10378 14864 19380 14920
rect 10317 14862 19380 14864
rect 10317 14859 10383 14862
rect 19374 14860 19380 14862
rect 19444 14860 19450 14924
rect 22050 14922 22110 14998
rect 22318 14996 22324 15060
rect 22388 15058 22394 15060
rect 23197 15058 23263 15061
rect 22388 15056 23263 15058
rect 22388 15000 23202 15056
rect 23258 15000 23263 15056
rect 22388 14998 23263 15000
rect 22388 14996 22394 14998
rect 23197 14995 23263 14998
rect 23381 15058 23447 15061
rect 26200 15058 27000 15088
rect 23381 15056 27000 15058
rect 23381 15000 23386 15056
rect 23442 15000 27000 15056
rect 23381 14998 27000 15000
rect 23381 14995 23447 14998
rect 26200 14968 27000 14998
rect 25129 14922 25195 14925
rect 22050 14920 25195 14922
rect 22050 14864 25134 14920
rect 25190 14864 25195 14920
rect 22050 14862 25195 14864
rect 25129 14859 25195 14862
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 26200 14650 27000 14680
rect 23430 14590 27000 14650
rect 8845 14514 8911 14517
rect 15510 14514 15516 14516
rect 8845 14512 15516 14514
rect 8845 14456 8850 14512
rect 8906 14456 15516 14512
rect 8845 14454 15516 14456
rect 8845 14451 8911 14454
rect 15510 14452 15516 14454
rect 15580 14452 15586 14516
rect 22737 14514 22803 14517
rect 23430 14514 23490 14590
rect 26200 14560 27000 14590
rect 22737 14512 23490 14514
rect 22737 14456 22742 14512
rect 22798 14456 23490 14512
rect 22737 14454 23490 14456
rect 22737 14451 22803 14454
rect 6545 14378 6611 14381
rect 22093 14378 22159 14381
rect 6545 14376 22159 14378
rect 6545 14320 6550 14376
rect 6606 14320 22098 14376
rect 22154 14320 22159 14376
rect 6545 14318 22159 14320
rect 6545 14315 6611 14318
rect 22093 14315 22159 14318
rect 23933 14242 23999 14245
rect 26200 14242 27000 14272
rect 23933 14240 27000 14242
rect 23933 14184 23938 14240
rect 23994 14184 27000 14240
rect 23933 14182 27000 14184
rect 23933 14179 23999 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 19517 14106 19583 14109
rect 19742 14106 19748 14108
rect 19517 14104 19748 14106
rect 19517 14048 19522 14104
rect 19578 14048 19748 14104
rect 19517 14046 19748 14048
rect 19517 14043 19583 14046
rect 19742 14044 19748 14046
rect 19812 14044 19818 14108
rect 20478 14044 20484 14108
rect 20548 14106 20554 14108
rect 23422 14106 23428 14108
rect 20548 14046 23428 14106
rect 20548 14044 20554 14046
rect 23422 14044 23428 14046
rect 23492 14044 23498 14108
rect 4337 13970 4403 13973
rect 25129 13970 25195 13973
rect 4337 13968 25195 13970
rect 4337 13912 4342 13968
rect 4398 13912 25134 13968
rect 25190 13912 25195 13968
rect 4337 13910 25195 13912
rect 4337 13907 4403 13910
rect 25129 13907 25195 13910
rect 10961 13834 11027 13837
rect 19558 13834 19564 13836
rect 10961 13832 19564 13834
rect 10961 13776 10966 13832
rect 11022 13776 19564 13832
rect 10961 13774 19564 13776
rect 10961 13771 11027 13774
rect 19558 13772 19564 13774
rect 19628 13772 19634 13836
rect 22645 13834 22711 13837
rect 26200 13834 27000 13864
rect 22645 13832 27000 13834
rect 22645 13776 22650 13832
rect 22706 13776 27000 13832
rect 22645 13774 27000 13776
rect 22645 13771 22711 13774
rect 26200 13744 27000 13774
rect 16389 13698 16455 13701
rect 20253 13698 20319 13701
rect 16389 13696 20319 13698
rect 16389 13640 16394 13696
rect 16450 13640 20258 13696
rect 20314 13640 20319 13696
rect 16389 13638 20319 13640
rect 16389 13635 16455 13638
rect 20253 13635 20319 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 22553 13426 22619 13429
rect 26200 13426 27000 13456
rect 22553 13424 27000 13426
rect 22553 13368 22558 13424
rect 22614 13368 27000 13424
rect 22553 13366 27000 13368
rect 22553 13363 22619 13366
rect 26200 13336 27000 13366
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 21817 13018 21883 13021
rect 26200 13018 27000 13048
rect 21817 13016 27000 13018
rect 21817 12960 21822 13016
rect 21878 12960 27000 13016
rect 21817 12958 27000 12960
rect 21817 12955 21883 12958
rect 26200 12928 27000 12958
rect 22185 12882 22251 12885
rect 22461 12882 22527 12885
rect 22185 12880 22527 12882
rect 22185 12824 22190 12880
rect 22246 12824 22466 12880
rect 22522 12824 22527 12880
rect 22185 12822 22527 12824
rect 22185 12819 22251 12822
rect 22461 12819 22527 12822
rect 9622 12684 9628 12748
rect 9692 12746 9698 12748
rect 9692 12686 16590 12746
rect 9692 12684 9698 12686
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 16530 12338 16590 12686
rect 24761 12610 24827 12613
rect 26200 12610 27000 12640
rect 24761 12608 27000 12610
rect 24761 12552 24766 12608
rect 24822 12552 27000 12608
rect 24761 12550 27000 12552
rect 24761 12547 24827 12550
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 18505 12474 18571 12477
rect 19149 12474 19215 12477
rect 19793 12476 19859 12477
rect 18505 12472 19215 12474
rect 18505 12416 18510 12472
rect 18566 12416 19154 12472
rect 19210 12416 19215 12472
rect 18505 12414 19215 12416
rect 18505 12411 18571 12414
rect 19149 12411 19215 12414
rect 19742 12412 19748 12476
rect 19812 12474 19859 12476
rect 19812 12472 19904 12474
rect 19854 12416 19904 12472
rect 19812 12414 19904 12416
rect 19812 12412 19859 12414
rect 19793 12411 19859 12412
rect 19885 12338 19951 12341
rect 16530 12336 19951 12338
rect 16530 12280 19890 12336
rect 19946 12280 19951 12336
rect 16530 12278 19951 12280
rect 19885 12275 19951 12278
rect 20805 12338 20871 12341
rect 21081 12338 21147 12341
rect 20805 12336 21147 12338
rect 20805 12280 20810 12336
rect 20866 12280 21086 12336
rect 21142 12280 21147 12336
rect 20805 12278 21147 12280
rect 20805 12275 20871 12278
rect 21081 12275 21147 12278
rect 21725 12338 21791 12341
rect 25037 12338 25103 12341
rect 21725 12336 25103 12338
rect 21725 12280 21730 12336
rect 21786 12280 25042 12336
rect 25098 12280 25103 12336
rect 21725 12278 25103 12280
rect 21725 12275 21791 12278
rect 25037 12275 25103 12278
rect 24669 12202 24735 12205
rect 26200 12202 27000 12232
rect 24669 12200 27000 12202
rect 24669 12144 24674 12200
rect 24730 12144 27000 12200
rect 24669 12142 27000 12144
rect 24669 12139 24735 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 21449 11930 21515 11933
rect 21582 11930 21588 11932
rect 21449 11928 21588 11930
rect 21449 11872 21454 11928
rect 21510 11872 21588 11928
rect 21449 11870 21588 11872
rect 21449 11867 21515 11870
rect 21582 11868 21588 11870
rect 21652 11868 21658 11932
rect 15101 11794 15167 11797
rect 20110 11794 20116 11796
rect 15101 11792 20116 11794
rect 15101 11736 15106 11792
rect 15162 11736 20116 11792
rect 15101 11734 20116 11736
rect 15101 11731 15167 11734
rect 20110 11732 20116 11734
rect 20180 11732 20186 11796
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 15653 11658 15719 11661
rect 25129 11658 25195 11661
rect 15653 11656 25195 11658
rect 15653 11600 15658 11656
rect 15714 11600 25134 11656
rect 25190 11600 25195 11656
rect 15653 11598 25195 11600
rect 15653 11595 15719 11598
rect 25129 11595 25195 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 16113 11386 16179 11389
rect 16246 11386 16252 11388
rect 16113 11384 16252 11386
rect 16113 11328 16118 11384
rect 16174 11328 16252 11384
rect 16113 11326 16252 11328
rect 16113 11323 16179 11326
rect 16246 11324 16252 11326
rect 16316 11324 16322 11388
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 15653 11250 15719 11253
rect 20662 11250 20668 11252
rect 15653 11248 20668 11250
rect 15653 11192 15658 11248
rect 15714 11192 20668 11248
rect 15653 11190 20668 11192
rect 15653 11187 15719 11190
rect 20662 11188 20668 11190
rect 20732 11188 20738 11252
rect 22185 11250 22251 11253
rect 22502 11250 22508 11252
rect 22185 11248 22508 11250
rect 22185 11192 22190 11248
rect 22246 11192 22508 11248
rect 22185 11190 22508 11192
rect 22185 11187 22251 11190
rect 22502 11188 22508 11190
rect 22572 11188 22578 11252
rect 19701 11114 19767 11117
rect 22188 11114 22248 11187
rect 19701 11112 22248 11114
rect 19701 11056 19706 11112
rect 19762 11056 22248 11112
rect 19701 11054 22248 11056
rect 19701 11051 19767 11054
rect 24761 10978 24827 10981
rect 26200 10978 27000 11008
rect 24761 10976 27000 10978
rect 24761 10920 24766 10976
rect 24822 10920 27000 10976
rect 24761 10918 27000 10920
rect 24761 10915 24827 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 17718 10644 17724 10708
rect 17788 10706 17794 10708
rect 18045 10706 18111 10709
rect 17788 10704 18111 10706
rect 17788 10648 18050 10704
rect 18106 10648 18111 10704
rect 17788 10646 18111 10648
rect 17788 10644 17794 10646
rect 18045 10643 18111 10646
rect 19517 10706 19583 10709
rect 25957 10706 26023 10709
rect 19517 10704 26023 10706
rect 19517 10648 19522 10704
rect 19578 10648 25962 10704
rect 26018 10648 26023 10704
rect 19517 10646 26023 10648
rect 19517 10643 19583 10646
rect 25957 10643 26023 10646
rect 17585 10570 17651 10573
rect 20478 10570 20484 10572
rect 17585 10568 20484 10570
rect 17585 10512 17590 10568
rect 17646 10512 20484 10568
rect 17585 10510 20484 10512
rect 17585 10507 17651 10510
rect 20478 10508 20484 10510
rect 20548 10508 20554 10572
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 15469 10298 15535 10301
rect 20713 10298 20779 10301
rect 15469 10296 20779 10298
rect 15469 10240 15474 10296
rect 15530 10240 20718 10296
rect 20774 10240 20779 10296
rect 15469 10238 20779 10240
rect 15469 10235 15535 10238
rect 20713 10235 20779 10238
rect 24577 10162 24643 10165
rect 26200 10162 27000 10192
rect 24577 10160 27000 10162
rect 24577 10104 24582 10160
rect 24638 10104 27000 10160
rect 24577 10102 27000 10104
rect 24577 10099 24643 10102
rect 26200 10072 27000 10102
rect 13486 9964 13492 10028
rect 13556 10026 13562 10028
rect 23841 10026 23907 10029
rect 13556 10024 23907 10026
rect 13556 9968 23846 10024
rect 23902 9968 23907 10024
rect 13556 9966 23907 9968
rect 13556 9964 13562 9966
rect 23841 9963 23907 9966
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 22645 9620 22711 9621
rect 22645 9618 22692 9620
rect 22600 9616 22692 9618
rect 22600 9560 22650 9616
rect 22600 9558 22692 9560
rect 22645 9556 22692 9558
rect 22756 9556 22762 9620
rect 22645 9555 22711 9556
rect 15878 9420 15884 9484
rect 15948 9482 15954 9484
rect 19425 9482 19491 9485
rect 15948 9480 19491 9482
rect 15948 9424 19430 9480
rect 19486 9424 19491 9480
rect 15948 9422 19491 9424
rect 15948 9420 15954 9422
rect 19425 9419 19491 9422
rect 20161 9482 20227 9485
rect 23473 9482 23539 9485
rect 20161 9480 23539 9482
rect 20161 9424 20166 9480
rect 20222 9424 23478 9480
rect 23534 9424 23539 9480
rect 20161 9422 23539 9424
rect 20161 9419 20227 9422
rect 23473 9419 23539 9422
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 24853 9283 24919 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 24669 8938 24735 8941
rect 26200 8938 27000 8968
rect 24669 8936 27000 8938
rect 24669 8880 24674 8936
rect 24730 8880 27000 8936
rect 24669 8878 27000 8880
rect 24669 8875 24735 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24853 8530 24919 8533
rect 26200 8530 27000 8560
rect 24853 8528 27000 8530
rect 24853 8472 24858 8528
rect 24914 8472 27000 8528
rect 24853 8470 27000 8472
rect 24853 8467 24919 8470
rect 26200 8440 27000 8470
rect 21449 8394 21515 8397
rect 21950 8394 21956 8396
rect 21449 8392 21956 8394
rect 21449 8336 21454 8392
rect 21510 8336 21956 8392
rect 21449 8334 21956 8336
rect 21449 8331 21515 8334
rect 21950 8332 21956 8334
rect 22020 8332 22026 8396
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 8122 25011 8125
rect 26200 8122 27000 8152
rect 24945 8120 27000 8122
rect 24945 8064 24950 8120
rect 25006 8064 27000 8120
rect 24945 8062 27000 8064
rect 24945 8059 25011 8062
rect 26200 8032 27000 8062
rect 13670 7788 13676 7852
rect 13740 7850 13746 7852
rect 21265 7850 21331 7853
rect 13740 7848 21331 7850
rect 13740 7792 21270 7848
rect 21326 7792 21331 7848
rect 13740 7790 21331 7792
rect 13740 7788 13746 7790
rect 21265 7787 21331 7790
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24853 6898 24919 6901
rect 26200 6898 27000 6928
rect 24853 6896 27000 6898
rect 24853 6840 24858 6896
rect 24914 6840 27000 6896
rect 24853 6838 27000 6840
rect 24853 6835 24919 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 22185 6354 22251 6357
rect 22318 6354 22324 6356
rect 22185 6352 22324 6354
rect 22185 6296 22190 6352
rect 22246 6296 22324 6352
rect 22185 6294 22324 6296
rect 22185 6291 22251 6294
rect 22318 6292 22324 6294
rect 22388 6292 22394 6356
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25129 4042 25195 4045
rect 26200 4042 27000 4072
rect 25129 4040 27000 4042
rect 25129 3984 25134 4040
rect 25190 3984 27000 4040
rect 25129 3982 27000 3984
rect 25129 3979 25195 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 24945 3226 25011 3229
rect 26200 3226 27000 3256
rect 24945 3224 27000 3226
rect 24945 3168 24950 3224
rect 25006 3168 27000 3224
rect 24945 3166 27000 3168
rect 24945 3163 25011 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22737 2002 22803 2005
rect 26200 2002 27000 2032
rect 22737 2000 27000 2002
rect 22737 1944 22742 2000
rect 22798 1944 27000 2000
rect 22737 1942 27000 1944
rect 22737 1939 22803 1942
rect 26200 1912 27000 1942
rect 22093 1594 22159 1597
rect 26200 1594 27000 1624
rect 22093 1592 27000 1594
rect 22093 1536 22098 1592
rect 22154 1536 27000 1592
rect 22093 1534 27000 1536
rect 22093 1531 22159 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 6684 25876 6748 25940
rect 4844 25604 4908 25668
rect 10548 25468 10612 25532
rect 19748 25332 19812 25396
rect 7604 25196 7668 25260
rect 22140 25196 22204 25260
rect 9444 25060 9508 25124
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 5396 24380 5460 24444
rect 16252 24108 16316 24172
rect 19196 23972 19260 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 14044 23836 14108 23900
rect 17540 23836 17604 23900
rect 18644 23564 18708 23628
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 13860 23292 13924 23356
rect 18828 22944 18892 22948
rect 18828 22888 18842 22944
rect 18842 22888 18892 22944
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 12756 22748 12820 22812
rect 18828 22884 18892 22888
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 21588 22476 21652 22540
rect 12756 22340 12820 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 13676 22128 13740 22132
rect 13676 22072 13690 22128
rect 13690 22072 13740 22128
rect 13676 22068 13740 22072
rect 21404 22068 21468 22132
rect 22324 21932 22388 21996
rect 9628 21796 9692 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 22508 21524 22572 21588
rect 14228 21252 14292 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 17356 20904 17420 20908
rect 17356 20848 17406 20904
rect 17406 20848 17420 20904
rect 17356 20844 17420 20848
rect 13492 20768 13556 20772
rect 13492 20712 13542 20768
rect 13542 20712 13556 20768
rect 13492 20708 13556 20712
rect 15884 20768 15948 20772
rect 15884 20712 15898 20768
rect 15898 20712 15948 20768
rect 15884 20708 15948 20712
rect 19564 20768 19628 20772
rect 19564 20712 19578 20768
rect 19578 20712 19628 20768
rect 19564 20708 19628 20712
rect 20668 20708 20732 20772
rect 22140 20708 22204 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 20116 20300 20180 20364
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12572 19892 12636 19956
rect 14044 20164 14108 20228
rect 15148 20164 15212 20228
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 17172 19892 17236 19956
rect 18460 19892 18524 19956
rect 5396 19620 5460 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 12572 19620 12636 19684
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18460 19484 18524 19548
rect 14228 19348 14292 19412
rect 17172 19348 17236 19412
rect 17356 19348 17420 19412
rect 17540 19348 17604 19412
rect 18828 19348 18892 19412
rect 19380 19348 19444 19412
rect 6684 19212 6748 19276
rect 17724 19076 17788 19140
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 15516 18396 15580 18460
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 19748 17988 19812 18052
rect 23428 17988 23492 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 4844 17716 4908 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 7604 17232 7668 17236
rect 7604 17176 7618 17232
rect 7618 17176 7668 17232
rect 7604 17172 7668 17176
rect 21956 17036 22020 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 19196 16764 19260 16828
rect 13860 16628 13924 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 15148 16084 15212 16148
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18644 15948 18708 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 21404 15676 21468 15740
rect 9444 15600 9508 15604
rect 9444 15544 9458 15600
rect 9458 15544 9508 15600
rect 9444 15540 9508 15544
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 22692 15268 22756 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 10548 15056 10612 15060
rect 10548 15000 10562 15056
rect 10562 15000 10612 15056
rect 10548 14996 10612 15000
rect 22140 15132 22204 15196
rect 19380 14860 19444 14924
rect 22324 14996 22388 15060
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 15516 14452 15580 14516
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 19748 14044 19812 14108
rect 20484 14044 20548 14108
rect 23428 14044 23492 14108
rect 19564 13772 19628 13836
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 9628 12684 9692 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 19748 12472 19812 12476
rect 19748 12416 19798 12472
rect 19798 12416 19812 12472
rect 19748 12412 19812 12416
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 21588 11868 21652 11932
rect 20116 11732 20180 11796
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 16252 11324 16316 11388
rect 20668 11188 20732 11252
rect 22508 11188 22572 11252
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 17724 10644 17788 10708
rect 20484 10508 20548 10572
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 13492 9964 13556 10028
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 22692 9616 22756 9620
rect 22692 9560 22706 9616
rect 22706 9560 22756 9616
rect 22692 9556 22756 9560
rect 15884 9420 15948 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 21956 8332 22020 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 13676 7788 13740 7852
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 22324 6292 22388 6356
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 6683 25940 6749 25941
rect 6683 25876 6684 25940
rect 6748 25876 6749 25940
rect 6683 25875 6749 25876
rect 4843 25668 4909 25669
rect 4843 25604 4844 25668
rect 4908 25604 4909 25668
rect 4843 25603 4909 25604
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 4846 17781 4906 25603
rect 5395 24444 5461 24445
rect 5395 24380 5396 24444
rect 5460 24380 5461 24444
rect 5395 24379 5461 24380
rect 5398 19685 5458 24379
rect 5395 19684 5461 19685
rect 5395 19620 5396 19684
rect 5460 19620 5461 19684
rect 5395 19619 5461 19620
rect 6686 19277 6746 25875
rect 10547 25532 10613 25533
rect 10547 25468 10548 25532
rect 10612 25468 10613 25532
rect 10547 25467 10613 25468
rect 7603 25260 7669 25261
rect 7603 25196 7604 25260
rect 7668 25196 7669 25260
rect 7603 25195 7669 25196
rect 6683 19276 6749 19277
rect 6683 19212 6684 19276
rect 6748 19212 6749 19276
rect 6683 19211 6749 19212
rect 4843 17780 4909 17781
rect 4843 17716 4844 17780
rect 4908 17716 4909 17780
rect 4843 17715 4909 17716
rect 7606 17237 7666 25195
rect 9443 25124 9509 25125
rect 9443 25060 9444 25124
rect 9508 25060 9509 25124
rect 9443 25059 9509 25060
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7603 17236 7669 17237
rect 7603 17172 7604 17236
rect 7668 17172 7669 17236
rect 7603 17171 7669 17172
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 9446 15605 9506 25059
rect 9627 21860 9693 21861
rect 9627 21796 9628 21860
rect 9692 21796 9693 21860
rect 9627 21795 9693 21796
rect 9443 15604 9509 15605
rect 9443 15540 9444 15604
rect 9508 15540 9509 15604
rect 9443 15539 9509 15540
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 9630 12749 9690 21795
rect 10550 15061 10610 25467
rect 19747 25396 19813 25397
rect 19747 25332 19748 25396
rect 19812 25332 19813 25396
rect 19747 25331 19813 25332
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 16251 24172 16317 24173
rect 16251 24108 16252 24172
rect 16316 24108 16317 24172
rect 16251 24107 16317 24108
rect 14043 23900 14109 23901
rect 14043 23836 14044 23900
rect 14108 23836 14109 23900
rect 14043 23835 14109 23836
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12755 22812 12821 22813
rect 12755 22748 12756 22812
rect 12820 22748 12821 22812
rect 12755 22747 12821 22748
rect 12758 22405 12818 22747
rect 12755 22404 12821 22405
rect 12755 22340 12756 22404
rect 12820 22340 12821 22404
rect 12755 22339 12821 22340
rect 12944 22336 13264 23360
rect 13859 23356 13925 23357
rect 13859 23292 13860 23356
rect 13924 23292 13925 23356
rect 13859 23291 13925 23292
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 13675 22132 13741 22133
rect 13675 22068 13676 22132
rect 13740 22068 13741 22132
rect 13675 22067 13741 22068
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 13491 20772 13557 20773
rect 13491 20708 13492 20772
rect 13556 20708 13557 20772
rect 13491 20707 13557 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12571 19956 12637 19957
rect 12571 19892 12572 19956
rect 12636 19892 12637 19956
rect 12571 19891 12637 19892
rect 12574 19685 12634 19891
rect 12571 19684 12637 19685
rect 12571 19620 12572 19684
rect 12636 19620 12637 19684
rect 12571 19619 12637 19620
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 10547 15060 10613 15061
rect 10547 14996 10548 15060
rect 10612 14996 10613 15060
rect 10547 14995 10613 14996
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 9627 12748 9693 12749
rect 9627 12684 9628 12748
rect 9692 12684 9693 12748
rect 9627 12683 9693 12684
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 13494 10029 13554 20707
rect 13491 10028 13557 10029
rect 13491 9964 13492 10028
rect 13556 9964 13557 10028
rect 13491 9963 13557 9964
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 13678 7853 13738 22067
rect 13862 16693 13922 23291
rect 14046 20229 14106 23835
rect 14227 21316 14293 21317
rect 14227 21252 14228 21316
rect 14292 21252 14293 21316
rect 14227 21251 14293 21252
rect 14043 20228 14109 20229
rect 14043 20164 14044 20228
rect 14108 20164 14109 20228
rect 14043 20163 14109 20164
rect 14230 19413 14290 21251
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 15147 20228 15213 20229
rect 15147 20164 15148 20228
rect 15212 20164 15213 20228
rect 15147 20163 15213 20164
rect 14227 19412 14293 19413
rect 14227 19348 14228 19412
rect 14292 19348 14293 19412
rect 14227 19347 14293 19348
rect 13859 16692 13925 16693
rect 13859 16628 13860 16692
rect 13924 16628 13925 16692
rect 13859 16627 13925 16628
rect 15150 16149 15210 20163
rect 15515 18460 15581 18461
rect 15515 18396 15516 18460
rect 15580 18396 15581 18460
rect 15515 18395 15581 18396
rect 15147 16148 15213 16149
rect 15147 16084 15148 16148
rect 15212 16084 15213 16148
rect 15147 16083 15213 16084
rect 15518 14517 15578 18395
rect 15515 14516 15581 14517
rect 15515 14452 15516 14516
rect 15580 14452 15581 14516
rect 15515 14451 15581 14452
rect 15886 9485 15946 20707
rect 16254 11389 16314 24107
rect 17944 23968 18264 24528
rect 19195 24036 19261 24037
rect 19195 23972 19196 24036
rect 19260 23972 19261 24036
rect 19195 23971 19261 23972
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17539 23900 17605 23901
rect 17539 23836 17540 23900
rect 17604 23836 17605 23900
rect 17539 23835 17605 23836
rect 17355 20908 17421 20909
rect 17355 20844 17356 20908
rect 17420 20844 17421 20908
rect 17355 20843 17421 20844
rect 17171 19956 17237 19957
rect 17171 19892 17172 19956
rect 17236 19892 17237 19956
rect 17171 19891 17237 19892
rect 17174 19413 17234 19891
rect 17358 19413 17418 20843
rect 17542 19413 17602 23835
rect 17944 22880 18264 23904
rect 18643 23628 18709 23629
rect 18643 23564 18644 23628
rect 18708 23564 18709 23628
rect 18643 23563 18709 23564
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 18459 19956 18525 19957
rect 18459 19892 18460 19956
rect 18524 19892 18525 19956
rect 18459 19891 18525 19892
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17171 19412 17237 19413
rect 17171 19348 17172 19412
rect 17236 19348 17237 19412
rect 17171 19347 17237 19348
rect 17355 19412 17421 19413
rect 17355 19348 17356 19412
rect 17420 19348 17421 19412
rect 17355 19347 17421 19348
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17723 19140 17789 19141
rect 17723 19076 17724 19140
rect 17788 19076 17789 19140
rect 17723 19075 17789 19076
rect 16251 11388 16317 11389
rect 16251 11324 16252 11388
rect 16316 11324 16317 11388
rect 16251 11323 16317 11324
rect 17726 10709 17786 19075
rect 17944 18528 18264 19552
rect 18462 19549 18522 19891
rect 18459 19548 18525 19549
rect 18459 19484 18460 19548
rect 18524 19484 18525 19548
rect 18459 19483 18525 19484
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 18646 16013 18706 23563
rect 18827 22948 18893 22949
rect 18827 22884 18828 22948
rect 18892 22884 18893 22948
rect 18827 22883 18893 22884
rect 18830 19413 18890 22883
rect 18827 19412 18893 19413
rect 18827 19348 18828 19412
rect 18892 19348 18893 19412
rect 18827 19347 18893 19348
rect 19198 16829 19258 23971
rect 19563 20772 19629 20773
rect 19563 20708 19564 20772
rect 19628 20708 19629 20772
rect 19563 20707 19629 20708
rect 19379 19412 19445 19413
rect 19379 19348 19380 19412
rect 19444 19348 19445 19412
rect 19379 19347 19445 19348
rect 19195 16828 19261 16829
rect 19195 16764 19196 16828
rect 19260 16764 19261 16828
rect 19195 16763 19261 16764
rect 18643 16012 18709 16013
rect 18643 15948 18644 16012
rect 18708 15948 18709 16012
rect 18643 15947 18709 15948
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 19382 14925 19442 19347
rect 19379 14924 19445 14925
rect 19379 14860 19380 14924
rect 19444 14860 19445 14924
rect 19379 14859 19445 14860
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 19566 13837 19626 20707
rect 19750 18053 19810 25331
rect 22139 25260 22205 25261
rect 22139 25196 22140 25260
rect 22204 25196 22205 25260
rect 22139 25195 22205 25196
rect 21587 22540 21653 22541
rect 21587 22476 21588 22540
rect 21652 22476 21653 22540
rect 21587 22475 21653 22476
rect 21403 22132 21469 22133
rect 21403 22068 21404 22132
rect 21468 22068 21469 22132
rect 21403 22067 21469 22068
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 20115 20364 20181 20365
rect 20115 20300 20116 20364
rect 20180 20300 20181 20364
rect 20115 20299 20181 20300
rect 19747 18052 19813 18053
rect 19747 17988 19748 18052
rect 19812 17988 19813 18052
rect 19747 17987 19813 17988
rect 19747 14108 19813 14109
rect 19747 14044 19748 14108
rect 19812 14044 19813 14108
rect 19747 14043 19813 14044
rect 19563 13836 19629 13837
rect 19563 13772 19564 13836
rect 19628 13772 19629 13836
rect 19563 13771 19629 13772
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 19750 12477 19810 14043
rect 19747 12476 19813 12477
rect 19747 12412 19748 12476
rect 19812 12412 19813 12476
rect 19747 12411 19813 12412
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 20118 11797 20178 20299
rect 20483 14108 20549 14109
rect 20483 14044 20484 14108
rect 20548 14044 20549 14108
rect 20483 14043 20549 14044
rect 20115 11796 20181 11797
rect 20115 11732 20116 11796
rect 20180 11732 20181 11796
rect 20115 11731 20181 11732
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17723 10708 17789 10709
rect 17723 10644 17724 10708
rect 17788 10644 17789 10708
rect 17723 10643 17789 10644
rect 17944 9824 18264 10848
rect 20486 10573 20546 14043
rect 20670 11253 20730 20707
rect 21406 15741 21466 22067
rect 21403 15740 21469 15741
rect 21403 15676 21404 15740
rect 21468 15676 21469 15740
rect 21403 15675 21469 15676
rect 21590 11933 21650 22475
rect 22142 20773 22202 25195
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22323 21996 22389 21997
rect 22323 21932 22324 21996
rect 22388 21932 22389 21996
rect 22323 21931 22389 21932
rect 22139 20772 22205 20773
rect 22139 20708 22140 20772
rect 22204 20708 22205 20772
rect 22139 20707 22205 20708
rect 21955 17100 22021 17101
rect 21955 17036 21956 17100
rect 22020 17036 22021 17100
rect 21955 17035 22021 17036
rect 21587 11932 21653 11933
rect 21587 11868 21588 11932
rect 21652 11868 21653 11932
rect 21587 11867 21653 11868
rect 20667 11252 20733 11253
rect 20667 11188 20668 11252
rect 20732 11188 20733 11252
rect 20667 11187 20733 11188
rect 20483 10572 20549 10573
rect 20483 10508 20484 10572
rect 20548 10508 20549 10572
rect 20483 10507 20549 10508
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 15883 9484 15949 9485
rect 15883 9420 15884 9484
rect 15948 9420 15949 9484
rect 15883 9419 15949 9420
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 13675 7852 13741 7853
rect 13675 7788 13676 7852
rect 13740 7788 13741 7852
rect 13675 7787 13741 7788
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 7648 18264 8672
rect 21958 8397 22018 17035
rect 22326 15330 22386 21931
rect 22507 21588 22573 21589
rect 22507 21524 22508 21588
rect 22572 21524 22573 21588
rect 22507 21523 22573 21524
rect 22142 15270 22386 15330
rect 22142 15197 22202 15270
rect 22139 15196 22205 15197
rect 22139 15132 22140 15196
rect 22204 15132 22205 15196
rect 22139 15131 22205 15132
rect 22323 15060 22389 15061
rect 22323 14996 22324 15060
rect 22388 14996 22389 15060
rect 22323 14995 22389 14996
rect 21955 8396 22021 8397
rect 21955 8332 21956 8396
rect 22020 8332 22021 8396
rect 21955 8331 22021 8332
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 22326 6357 22386 14995
rect 22510 11253 22570 21523
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 23427 18052 23493 18053
rect 23427 17988 23428 18052
rect 23492 17988 23493 18052
rect 23427 17987 23493 17988
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22691 15332 22757 15333
rect 22691 15268 22692 15332
rect 22756 15268 22757 15332
rect 22691 15267 22757 15268
rect 22507 11252 22573 11253
rect 22507 11188 22508 11252
rect 22572 11188 22573 11252
rect 22507 11187 22573 11188
rect 22694 9621 22754 15267
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 23430 14109 23490 17987
rect 23427 14108 23493 14109
rect 23427 14044 23428 14108
rect 23492 14044 23493 14108
rect 23427 14043 23493 14044
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22691 9620 22757 9621
rect 22691 9556 22692 9620
rect 22756 9556 22757 9620
rect 22691 9555 22757 9556
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22323 6356 22389 6357
rect 22323 6292 22324 6356
rect 22388 6292 22389 6356
rect 22323 6291 22389 6292
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1676037725
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1676037725
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1676037725
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1676037725
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1676037725
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1676037725
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1676037725
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 5152 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1676037725
transform 1 0 5152 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 15364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1676037725
transform 1 0 20516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1676037725
transform 1 0 25300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1676037725
transform 1 0 16192 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform 1 0 20240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1676037725
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 25300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold8_A
timestamp 1676037725
transform 1 0 6440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 22080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 21344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2024 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 2668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 6440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 1472 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 8556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 25392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 1656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1676037725
transform 1 0 1472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 2208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 25208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 6716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14996 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 4140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1676037725
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1676037725
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1676037725
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1676037725
transform 1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1676037725
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_70
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1676037725
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_70
timestamp 1676037725
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1676037725
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1676037725
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_225
timestamp 1676037725
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1676037725
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1676037725
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1676037725
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1676037725
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_221
timestamp 1676037725
transform 1 0 21436 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1676037725
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1676037725
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_226
timestamp 1676037725
transform 1 0 21896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1676037725
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1676037725
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1676037725
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_213
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1676037725
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_222
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1676037725
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1676037725
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1676037725
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1676037725
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1676037725
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_241
timestamp 1676037725
transform 1 0 23276 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1676037725
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1676037725
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1676037725
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1676037725
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1676037725
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_214
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1676037725
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1676037725
transform 1 0 21896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_232
timestamp 1676037725
transform 1 0 22448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_258
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_171
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_257
timestamp 1676037725
transform 1 0 24748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_126
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1676037725
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1676037725
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_199
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1676037725
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1676037725
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1676037725
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1676037725
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1676037725
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_249
timestamp 1676037725
transform 1 0 24012 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1676037725
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_90
timestamp 1676037725
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1676037725
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_263
timestamp 1676037725
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1676037725
transform 1 0 4324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1676037725
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_49
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1676037725
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1676037725
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1676037725
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_8
timestamp 1676037725
transform 1 0 1840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1676037725
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1676037725
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1676037725
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1676037725
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1676037725
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1676037725
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_187
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1676037725
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1676037725
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1676037725
transform 1 0 1840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_14
timestamp 1676037725
transform 1 0 2392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1676037725
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1676037725
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1676037725
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_247
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_12
timestamp 1676037725
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_19
timestamp 1676037725
transform 1 0 2852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1676037725
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1676037725
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1676037725
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1676037725
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_206
timestamp 1676037725
transform 1 0 20056 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1676037725
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_219
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1676037725
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_40
timestamp 1676037725
transform 1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1676037725
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1676037725
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1676037725
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_171
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_214
timestamp 1676037725
transform 1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1676037725
transform 1 0 1932 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_13
timestamp 1676037725
transform 1 0 2300 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_63
timestamp 1676037725
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1676037725
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1676037725
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_241
timestamp 1676037725
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1676037725
transform 1 0 6532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1676037725
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1676037725
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1676037725
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1676037725
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1676037725
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1676037725
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_8
timestamp 1676037725
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1676037725
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_96
timestamp 1676037725
transform 1 0 9936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_124
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1676037725
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_8
timestamp 1676037725
transform 1 0 1840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1676037725
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_68
timestamp 1676037725
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1676037725
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1676037725
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1676037725
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1676037725
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_203
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_8
timestamp 1676037725
transform 1 0 1840 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1676037725
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1676037725
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1676037725
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_139
timestamp 1676037725
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_150
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1676037725
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_227
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1676037725
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_143
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1676037725
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_162
timestamp 1676037725
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1676037725
transform 1 0 17664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1676037725
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1676037725
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_227
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold5
timestamp 1676037725
transform 1 0 14444 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 5152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 6624 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 23184 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 2024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__165
timestamp 1676037725
transform 1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__134
timestamp 1676037725
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__139
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__140
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 5336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__162
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__164
timestamp 1676037725
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__166
timestamp 1676037725
transform 1 0 25024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__167
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__132
timestamp 1676037725
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__133
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__135
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__136
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__137
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__138
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__141
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__147
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15732 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__157
timestamp 1676037725
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 20608 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__142
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__143
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__144
timestamp 1676037725
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__145
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__146
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__148
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__149
timestamp 1676037725
transform 1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__150
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal1 6670 2822 6670 2822 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal1 21620 8466 21620 8466 0 chanx_right_in[0]
rlabel metal2 21482 7871 21482 7871 0 chanx_right_in[10]
rlabel metal2 16882 17391 16882 17391 0 chanx_right_in[11]
rlabel metal1 13984 15674 13984 15674 0 chanx_right_in[12]
rlabel metal1 13478 18836 13478 18836 0 chanx_right_in[13]
rlabel metal3 17204 17476 17204 17476 0 chanx_right_in[14]
rlabel metal2 14766 17561 14766 17561 0 chanx_right_in[15]
rlabel metal1 13478 13906 13478 13906 0 chanx_right_in[16]
rlabel metal2 13846 14858 13846 14858 0 chanx_right_in[17]
rlabel metal3 12604 16048 12604 16048 0 chanx_right_in[18]
rlabel viali 7406 17172 7406 17172 0 chanx_right_in[19]
rlabel metal1 17894 12954 17894 12954 0 chanx_right_in[1]
rlabel metal1 22678 9112 22678 9112 0 chanx_right_in[20]
rlabel metal1 18906 10710 18906 10710 0 chanx_right_in[21]
rlabel metal3 18860 12444 18860 12444 0 chanx_right_in[22]
rlabel metal2 21482 11356 21482 11356 0 chanx_right_in[23]
rlabel via2 25162 11645 25162 11645 0 chanx_right_in[24]
rlabel metal3 21229 20740 21229 20740 0 chanx_right_in[25]
rlabel metal2 14490 16490 14490 16490 0 chanx_right_in[26]
rlabel metal1 11270 14042 11270 14042 0 chanx_right_in[27]
rlabel via2 10534 15011 10534 15011 0 chanx_right_in[28]
rlabel metal3 17250 25024 17250 25024 0 chanx_right_in[29]
rlabel metal1 22333 10778 22333 10778 0 chanx_right_in[2]
rlabel metal1 22264 4590 22264 4590 0 chanx_right_in[3]
rlabel metal1 19228 13294 19228 13294 0 chanx_right_in[4]
rlabel metal1 18446 12614 18446 12614 0 chanx_right_in[5]
rlabel metal2 22586 9401 22586 9401 0 chanx_right_in[6]
rlabel metal1 24656 9146 24656 9146 0 chanx_right_in[7]
rlabel metal2 22126 12036 22126 12036 0 chanx_right_in[8]
rlabel metal1 19596 13430 19596 13430 0 chanx_right_in[9]
rlabel metal2 25070 1853 25070 1853 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24380 6834 24380 6834 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal3 25584 7684 25584 7684 0 chanx_right_out[17]
rlabel metal1 24426 7922 24426 7922 0 chanx_right_out[18]
rlabel metal1 24104 8534 24104 8534 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 24702 8109 24702 8109 0 chanx_right_out[20]
rlabel metal1 24380 9010 24380 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal2 24610 9265 24610 9265 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 24794 10217 24794 10217 0 chanx_right_out[25]
rlabel metal1 24380 11186 24380 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24702 11373 24702 11373 0 chanx_right_out[28]
rlabel metal3 25584 12580 25584 12580 0 chanx_right_out[29]
rlabel metal2 22126 2805 22126 2805 0 chanx_right_out[2]
rlabel metal1 21160 2482 21160 2482 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25676 3196 25676 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 25162 3553 25162 3553 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel metal1 2346 18258 2346 18258 0 chany_top_in[0]
rlabel metal2 16422 25629 16422 25629 0 chany_top_in[10]
rlabel metal1 16652 21318 16652 21318 0 chany_top_in[11]
rlabel metal1 18032 19958 18032 19958 0 chany_top_in[12]
rlabel metal1 1656 17646 1656 17646 0 chany_top_in[13]
rlabel metal2 16698 16116 16698 16116 0 chany_top_in[14]
rlabel metal2 17572 19482 17572 19482 0 chany_top_in[15]
rlabel metal2 18446 25585 18446 25585 0 chany_top_in[16]
rlabel metal2 18998 26105 18998 26105 0 chany_top_in[17]
rlabel metal1 7866 18292 7866 18292 0 chany_top_in[18]
rlabel metal2 19734 26173 19734 26173 0 chany_top_in[19]
rlabel metal1 4738 18938 4738 18938 0 chany_top_in[1]
rlabel metal2 20102 25969 20102 25969 0 chany_top_in[20]
rlabel metal2 20194 26248 20194 26248 0 chany_top_in[21]
rlabel metal3 12604 22848 12604 22848 0 chany_top_in[22]
rlabel metal3 17549 23324 17549 23324 0 chany_top_in[23]
rlabel metal2 15042 20417 15042 20417 0 chany_top_in[24]
rlabel metal2 12650 23409 12650 23409 0 chany_top_in[25]
rlabel metal2 2162 20298 2162 20298 0 chany_top_in[26]
rlabel metal1 10166 15470 10166 15470 0 chany_top_in[27]
rlabel metal2 22901 26316 22901 26316 0 chany_top_in[28]
rlabel metal3 18354 13668 18354 13668 0 chany_top_in[29]
rlabel metal2 13478 24252 13478 24252 0 chany_top_in[2]
rlabel metal1 9016 16694 9016 16694 0 chany_top_in[3]
rlabel metal2 13938 24667 13938 24667 0 chany_top_in[4]
rlabel metal2 9338 24004 9338 24004 0 chany_top_in[5]
rlabel metal2 14950 24728 14950 24728 0 chany_top_in[6]
rlabel metal1 20470 20230 20470 20230 0 chany_top_in[7]
rlabel metal1 14030 23256 14030 23256 0 chany_top_in[8]
rlabel metal2 13294 23018 13294 23018 0 chany_top_in[9]
rlabel metal1 2070 19278 2070 19278 0 chany_top_out[0]
rlabel metal1 4692 23766 4692 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 6992 20978 6992 20978 0 chany_top_out[14]
rlabel metal2 7268 21454 7268 21454 0 chany_top_out[15]
rlabel metal2 5842 24242 5842 24242 0 chany_top_out[16]
rlabel metal1 7130 23154 7130 23154 0 chany_top_out[17]
rlabel metal1 8188 22066 8188 22066 0 chany_top_out[18]
rlabel metal1 7268 24106 7268 24106 0 chany_top_out[19]
rlabel metal1 2300 19890 2300 19890 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8234 23188 8234 23188 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9660 23766 9660 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal1 11132 24242 11132 24242 0 chany_top_out[26]
rlabel metal1 11914 23154 11914 23154 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel metal1 12650 24276 12650 24276 0 chany_top_out[29]
rlabel metal2 2714 24888 2714 24888 0 chany_top_out[2]
rlabel metal1 3220 26418 3220 26418 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4324 20978 4324 20978 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3956 23154 3956 23154 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal1 21758 18326 21758 18326 0 clknet_0_prog_clk
rlabel metal1 10488 13158 10488 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15640 15538 15640 15538 0 clknet_3_1__leaf_prog_clk
rlabel metal2 9062 20978 9062 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 14076 18394 14076 18394 0 clknet_3_3__leaf_prog_clk
rlabel metal1 16928 14926 16928 14926 0 clknet_3_4__leaf_prog_clk
rlabel metal1 20838 13362 20838 13362 0 clknet_3_5__leaf_prog_clk
rlabel metal1 20378 18700 20378 18700 0 clknet_3_6__leaf_prog_clk
rlabel metal1 23368 21522 23368 21522 0 clknet_3_7__leaf_prog_clk
rlabel metal2 8694 4454 8694 4454 0 net1
rlabel metal4 19596 17272 19596 17272 0 net10
rlabel metal1 24794 3026 24794 3026 0 net100
rlabel via3 22701 9588 22701 9588 0 net101
rlabel metal1 1978 19380 1978 19380 0 net102
rlabel metal2 19274 22967 19274 22967 0 net103
rlabel metal2 13386 21437 13386 21437 0 net104
rlabel metal2 6486 19924 6486 19924 0 net105
rlabel metal1 3082 24174 3082 24174 0 net106
rlabel metal1 7498 17850 7498 17850 0 net107
rlabel metal1 7728 17034 7728 17034 0 net108
rlabel metal2 12742 23154 12742 23154 0 net109
rlabel metal3 17756 18428 17756 18428 0 net11
rlabel metal1 14996 19958 14996 19958 0 net110
rlabel metal1 19550 22202 19550 22202 0 net111
rlabel metal2 18722 24072 18722 24072 0 net112
rlabel metal2 2254 19601 2254 19601 0 net113
rlabel metal1 2691 18870 2691 18870 0 net114
rlabel metal1 6072 19482 6072 19482 0 net115
rlabel metal1 6394 17306 6394 17306 0 net116
rlabel metal1 5152 19346 5152 19346 0 net117
rlabel metal1 7498 18802 7498 18802 0 net118
rlabel metal2 6210 21675 6210 21675 0 net119
rlabel metal2 15318 19601 15318 19601 0 net12
rlabel metal1 7452 19890 7452 19890 0 net120
rlabel metal1 10856 23086 10856 23086 0 net121
rlabel metal1 5750 17714 5750 17714 0 net122
rlabel metal2 12558 24293 12558 24293 0 net123
rlabel metal1 2254 20944 2254 20944 0 net124
rlabel metal2 15962 20281 15962 20281 0 net125
rlabel metal2 2714 20026 2714 20026 0 net126
rlabel metal1 2990 21590 2990 21590 0 net127
rlabel metal2 5842 19652 5842 19652 0 net128
rlabel metal1 3772 22610 3772 22610 0 net129
rlabel metal1 14628 20910 14628 20910 0 net13
rlabel metal2 13662 21267 13662 21267 0 net130
rlabel metal2 15134 21886 15134 21886 0 net131
rlabel metal1 20792 15402 20792 15402 0 net132
rlabel metal1 19274 14314 19274 14314 0 net133
rlabel metal1 4738 18190 4738 18190 0 net134
rlabel metal1 17710 12274 17710 12274 0 net135
rlabel metal1 18952 12818 18952 12818 0 net136
rlabel metal1 21160 12818 21160 12818 0 net137
rlabel metal1 23966 9962 23966 9962 0 net138
rlabel metal2 20194 13481 20194 13481 0 net139
rlabel via3 15893 20740 15893 20740 0 net14
rlabel metal2 13570 14654 13570 14654 0 net140
rlabel metal1 20240 19822 20240 19822 0 net141
rlabel metal2 14306 20706 14306 20706 0 net142
rlabel metal1 12512 21658 12512 21658 0 net143
rlabel metal2 4738 16286 4738 16286 0 net144
rlabel metal2 10074 20774 10074 20774 0 net145
rlabel metal1 9614 19754 9614 19754 0 net146
rlabel metal1 18354 20910 18354 20910 0 net147
rlabel metal1 9384 18734 9384 18734 0 net148
rlabel metal2 12466 20672 12466 20672 0 net149
rlabel metal1 18262 10506 18262 10506 0 net15
rlabel metal1 12144 18394 12144 18394 0 net150
rlabel metal2 11178 18122 11178 18122 0 net151
rlabel metal2 15410 15861 15410 15861 0 net152
rlabel metal1 10488 16218 10488 16218 0 net153
rlabel metal1 13478 15470 13478 15470 0 net154
rlabel metal2 13938 15606 13938 15606 0 net155
rlabel metal1 14030 17714 14030 17714 0 net156
rlabel metal2 15410 23953 15410 23953 0 net157
rlabel metal1 17572 23834 17572 23834 0 net158
rlabel metal1 22218 19414 22218 19414 0 net159
rlabel metal3 17503 19108 17503 19108 0 net16
rlabel metal2 21298 14994 21298 14994 0 net160
rlabel metal2 12558 15623 12558 15623 0 net161
rlabel metal1 22908 6834 22908 6834 0 net162
rlabel metal1 22862 9010 22862 9010 0 net163
rlabel metal1 22494 7854 22494 7854 0 net164
rlabel via2 2254 17731 2254 17731 0 net165
rlabel via2 25070 12291 25070 12291 0 net166
rlabel metal1 21344 15470 21344 15470 0 net167
rlabel metal1 23782 16762 23782 16762 0 net168
rlabel metal2 2346 24242 2346 24242 0 net169
rlabel metal2 17020 17306 17020 17306 0 net17
rlabel metal2 25254 16388 25254 16388 0 net170
rlabel metal1 21528 17238 21528 17238 0 net171
rlabel metal1 20102 22644 20102 22644 0 net172
rlabel metal2 7222 2890 7222 2890 0 net173
rlabel metal1 9844 8874 9844 8874 0 net174
rlabel metal2 7498 3332 7498 3332 0 net175
rlabel metal1 6831 2414 6831 2414 0 net176
rlabel metal2 15134 11645 15134 11645 0 net18
rlabel metal1 16100 23766 16100 23766 0 net19
rlabel metal1 16082 19754 16082 19754 0 net2
rlabel via2 13386 20757 13386 20757 0 net20
rlabel metal1 11868 14042 11868 14042 0 net21
rlabel metal4 19412 17136 19412 17136 0 net22
rlabel metal2 13938 18904 13938 18904 0 net23
rlabel metal1 15686 20434 15686 20434 0 net24
rlabel metal1 18170 17578 18170 17578 0 net25
rlabel metal1 19228 13498 19228 13498 0 net26
rlabel metal1 17112 17170 17112 17170 0 net27
rlabel metal1 17342 9350 17342 9350 0 net28
rlabel metal2 23874 9945 23874 9945 0 net29
rlabel metal1 13248 21930 13248 21930 0 net3
rlabel metal2 15962 19924 15962 19924 0 net30
rlabel metal1 17480 22542 17480 22542 0 net31
rlabel metal2 2806 18955 2806 18955 0 net32
rlabel metal2 4462 18717 4462 18717 0 net33
rlabel metal2 21574 15878 21574 15878 0 net34
rlabel metal2 18630 16490 18630 16490 0 net35
rlabel metal1 19642 18190 19642 18190 0 net36
rlabel metal1 17434 16422 17434 16422 0 net37
rlabel metal1 15640 14790 15640 14790 0 net38
rlabel metal1 7222 19482 7222 19482 0 net39
rlabel metal2 8418 17408 8418 17408 0 net4
rlabel metal3 12420 15096 12420 15096 0 net40
rlabel metal2 16514 17663 16514 17663 0 net41
rlabel metal3 17204 18904 17204 18904 0 net42
rlabel metal1 3680 18394 3680 18394 0 net43
rlabel metal2 8510 17051 8510 17051 0 net44
rlabel metal2 8234 18649 8234 18649 0 net45
rlabel metal3 14812 17748 14812 17748 0 net46
rlabel metal3 17204 16252 17204 16252 0 net47
rlabel metal1 13294 21386 13294 21386 0 net48
rlabel metal1 25852 9146 25852 9146 0 net49
rlabel metal1 12926 14280 12926 14280 0 net5
rlabel metal1 2208 18938 2208 18938 0 net50
rlabel metal2 17342 24038 17342 24038 0 net51
rlabel metal1 19504 9894 19504 9894 0 net52
rlabel via2 1610 24123 1610 24123 0 net53
rlabel metal1 19964 11118 19964 11118 0 net54
rlabel metal2 6578 15657 6578 15657 0 net55
rlabel metal1 25530 11254 25530 11254 0 net56
rlabel metal1 20976 16082 20976 16082 0 net57
rlabel metal2 4002 24871 4002 24871 0 net58
rlabel metal1 18998 18598 18998 18598 0 net59
rlabel metal1 13386 16184 13386 16184 0 net6
rlabel metal4 15548 16456 15548 16456 0 net60
rlabel metal4 18676 19788 18676 19788 0 net61
rlabel metal1 15870 24242 15870 24242 0 net62
rlabel metal1 17940 18258 17940 18258 0 net63
rlabel metal1 18676 18734 18676 18734 0 net64
rlabel metal1 20930 17544 20930 17544 0 net65
rlabel metal1 20976 19482 20976 19482 0 net66
rlabel metal1 13064 19142 13064 19142 0 net67
rlabel metal1 18722 17850 18722 17850 0 net68
rlabel metal2 2254 22304 2254 22304 0 net69
rlabel metal2 8602 17816 8602 17816 0 net7
rlabel metal1 17664 17510 17664 17510 0 net70
rlabel metal1 21482 2414 21482 2414 0 net71
rlabel metal1 20102 3060 20102 3060 0 net72
rlabel metal1 22862 5202 22862 5202 0 net73
rlabel metal1 23966 4148 23966 4148 0 net74
rlabel metal1 23184 5678 23184 5678 0 net75
rlabel metal1 22310 6358 22310 6358 0 net76
rlabel metal1 23920 5202 23920 5202 0 net77
rlabel metal1 22678 6732 22678 6732 0 net78
rlabel metal1 22310 7344 22310 7344 0 net79
rlabel metal1 3312 17510 3312 17510 0 net8
rlabel metal1 24840 6290 24840 6290 0 net80
rlabel metal1 23506 7854 23506 7854 0 net81
rlabel metal1 22126 8432 22126 8432 0 net82
rlabel metal1 20700 3502 20700 3502 0 net83
rlabel metal1 23184 7378 23184 7378 0 net84
rlabel metal1 21482 6630 21482 6630 0 net85
rlabel metal1 22126 9588 22126 9588 0 net86
rlabel metal1 23092 8466 23092 8466 0 net87
rlabel metal1 22126 10608 22126 10608 0 net88
rlabel metal1 21988 10506 21988 10506 0 net89
rlabel metal1 13570 14042 13570 14042 0 net9
rlabel metal1 22678 11186 22678 11186 0 net90
rlabel metal1 22126 11696 22126 11696 0 net91
rlabel metal2 23966 11356 23966 11356 0 net92
rlabel metal2 23598 9860 23598 9860 0 net93
rlabel metal1 20608 13838 20608 13838 0 net94
rlabel metal1 19136 3026 19136 3026 0 net95
rlabel metal1 23736 2414 23736 2414 0 net96
rlabel metal2 22310 3740 22310 3740 0 net97
rlabel metal1 23184 3502 23184 3502 0 net98
rlabel metal1 22862 4114 22862 4114 0 net99
rlabel metal2 18998 15606 18998 15606 0 prog_clk
rlabel metal1 24334 16082 24334 16082 0 prog_reset
rlabel metal1 1886 23222 1886 23222 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 20654 23681 20654 23681 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 24886 11050 24886 11050 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 20654 22083 20654 22083 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 15226 16626 15226 16626 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal2 19918 19822 19918 19822 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal2 19734 19193 19734 19193 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25254 19516 25254 19516 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal2 23966 18870 23966 18870 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal1 25116 19482 25116 19482 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 22218 16932 22218 16932 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal2 21666 19278 21666 19278 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 23966 15572 23966 15572 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22586 17850 22586 17850 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 23598 12274 23598 12274 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24518 15130 24518 15130 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal1 23000 12954 23000 12954 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 23230 12410 23230 12410 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal2 21942 22474 21942 22474 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 21160 20570 21160 20570 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 21298 13872 21298 13872 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 20509 13498 20509 13498 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 20194 16422 20194 16422 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 20739 16762 20739 16762 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal2 18906 15980 18906 15980 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal2 20102 19482 20102 19482 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal2 18630 14620 18630 14620 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal1 19274 15674 19274 15674 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal1 25392 18190 25392 18190 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal1 18722 24276 18722 24276 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17296 13158 17296 13158 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18492 14518 18492 14518 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 19136 12682 19136 12682 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 17756 12750 17756 12750 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20654 12682 20654 12682 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal1 20240 17714 20240 17714 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal2 21206 12155 21206 12155 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 24380 22406 24380 22406 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 17664 23630 17664 23630 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 17526 21556 17526 21556 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15916 18666 15916 18666 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal1 20424 19890 20424 19890 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 15088 22746 15088 22746 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 15226 20298 15226 20298 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal1 15318 21862 15318 21862 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal2 12834 21216 12834 21216 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal1 14582 19482 14582 19482 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal2 12466 22304 12466 22304 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal2 12742 21454 12742 21454 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 10534 20672 10534 20672 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal1 12282 22474 12282 22474 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 10810 18768 10810 18768 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 10810 19754 10810 19754 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 19136 20978 19136 20978 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal2 20930 20264 20930 20264 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 10074 17340 10074 17340 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal1 11224 18122 11224 18122 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12650 18207 12650 18207 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel metal1 14306 17034 14306 17034 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12374 17306 12374 17306 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 15134 17510 15134 17510 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 12282 14892 12282 14892 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal2 13478 16728 13478 16728 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20424 24242 20424 24242 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal1 20470 23154 20470 23154 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 11086 15402 11086 15402 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal1 15134 14960 15134 14960 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14398 13226 14398 13226 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 13984 13430 13984 13430 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14582 15232 14582 15232 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 16928 13498 16928 13498 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16422 14246 16422 14246 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 16560 23154 16560 23154 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal1 17112 22678 17112 22678 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 16790 22984 16790 22984 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 21574 8058 21574 8058 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 17503 21318 17503 21318 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 19482 20056 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24886 12818 24886 12818 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18630 5882 18630 5882 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 24564 21862 24564 21862 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 22287 6324 22287 6324 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 11254 24058 11254 0 sb_0__0_.mux_right_track_12.out
rlabel metal1 22218 16218 22218 16218 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23782 11118 23782 11118 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 10098 19688 10098 0 sb_0__0_.mux_right_track_14.out
rlabel metal2 23874 18224 23874 18224 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21758 10642 21758 10642 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21482 6800 21482 6800 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 23644 14450 23644 14450 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19826 10642 19826 10642 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 7854 19826 7854 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 24978 13362 24978 13362 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18906 13192 18906 13192 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13892 12206 13892 12206 0 sb_0__0_.mux_right_track_2.out
rlabel metal2 24978 24038 24978 24038 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 14812 19244 14812 19244 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20838 8602 20838 8602 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 20930 14042 20930 14042 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 10642 20792 10642 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 9044 19458 9044 0 sb_0__0_.mux_right_track_30.out
rlabel metal2 21206 17510 21206 17510 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21298 8942 21298 8942 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22126 8466 22126 8466 0 sb_0__0_.mux_right_track_32.out
rlabel metal2 20010 18326 20010 18326 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22218 7888 22218 7888 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 7854 24702 7854 0 sb_0__0_.mux_right_track_34.out
rlabel metal1 19688 14382 19688 14382 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19780 14518 19780 14518 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15226 15300 15226 15300 0 sb_0__0_.mux_right_track_4.out
rlabel metal1 18538 24038 18538 24038 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15042 17459 15042 17459 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 6766 23782 6766 0 sb_0__0_.mux_right_track_44.out
rlabel metal2 17526 16048 17526 16048 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 14042 17112 14042 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24886 5712 24886 5712 0 sb_0__0_.mux_right_track_46.out
rlabel metal1 19320 12954 19320 12954 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19182 12614 19182 12614 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24104 4590 24104 4590 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20194 12954 20194 12954 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 7378 20562 7378 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 3502 24702 3502 0 sb_0__0_.mux_right_track_50.out
rlabel metal1 25438 10030 25438 10030 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21850 7956 21850 7956 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13386 9554 13386 9554 0 sb_0__0_.mux_right_track_6.out
rlabel metal2 16882 23392 16882 23392 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24748 17850 24748 17850 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12466 16065 12466 16065 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19734 10336 19734 10336 0 sb_0__0_.mux_right_track_8.out
rlabel metal4 17572 21624 17572 21624 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 19067 10540 19067 10540 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4646 17102 4646 17102 0 sb_0__0_.mux_top_track_0.out
rlabel metal2 14306 19176 14306 19176 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15456 19482 15456 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 19618 14950 19618 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7176 18802 7176 18802 0 sb_0__0_.mux_top_track_10.out
rlabel metal1 17710 21896 17710 21896 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8602 20876 8602 20876 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2898 18836 2898 18836 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 15226 21114 15226 21114 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3082 18258 3082 18258 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6026 17204 6026 17204 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 16422 22134 16422 22134 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11500 22406 11500 22406 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8326 18904 8326 18904 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 14536 21046 14536 21046 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8510 19652 8510 19652 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2806 18700 2806 18700 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 11178 19754 11178 19754 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8740 20026 8740 20026 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13570 22797 13570 22797 0 sb_0__0_.mux_top_track_2.out
rlabel metal1 18354 21046 18354 21046 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17848 21114 17848 21114 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel viali 8050 17172 8050 17172 0 sb_0__0_.mux_top_track_28.out
rlabel metal1 14996 18394 14996 18394 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3450 18802 3450 18802 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7176 17714 7176 17714 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 16790 20026 16790 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8510 24344 8510 24344 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7176 18938 7176 18938 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 15778 18122 15778 18122 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11822 18156 11822 18156 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6670 19482 6670 19482 0 sb_0__0_.mux_top_track_34.out
rlabel metal2 15042 16864 15042 16864 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10810 16150 10810 16150 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12558 24072 12558 24072 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 22678 21114 22678 21114 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17710 24174 17710 24174 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4738 18292 4738 18292 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 13386 15912 13386 15912 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10028 15946 10028 15946 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6486 18258 6486 18258 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13846 15402 13846 15402 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12374 15317 12374 15317 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7544 22678 7544 22678 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 19366 16184 19366 16184 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13570 15742 13570 15742 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5382 18972 5382 18972 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 15318 17850 15318 17850 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9430 18836 9430 18836 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5290 17034 5290 17034 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 16192 21658 16192 21658 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 23086 17158 23086 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal4 12788 22576 12788 22576 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 5198 20468 5198 20468 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 19780 21658 19780 21658 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 23800 14122 23800 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1702 22882 1702 22882 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1932 20502 1932 20502 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 1610 22746 1610 22746 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 1564 21590 1564 21590 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
