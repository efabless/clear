VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 86.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 82.000 37.170 86.000 ;
    END
  END IO_ISOL_N
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 82.000 30.730 86.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 82.000 33.950 86.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END bottom_grid_pin_16_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END bottom_grid_pin_8_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 64.640 100.000 65.240 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.680 100.000 67.280 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.720 100.000 69.320 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.760 100.000 71.360 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 73.480 100.000 74.080 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 75.520 100.000 76.120 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.560 100.000 78.160 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 79.600 100.000 80.200 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 81.640 100.000 82.240 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 83.680 100.000 84.280 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 45.600 100.000 46.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 49.680 100.000 50.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.720 100.000 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 53.760 100.000 54.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 58.520 100.000 59.120 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 60.560 100.000 61.160 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 62.600 100.000 63.200 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 0.720 100.000 1.320 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 21.800 100.000 22.400 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 23.840 100.000 24.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.880 100.000 26.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.920 100.000 28.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 30.640 100.000 31.240 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 32.680 100.000 33.280 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 34.720 100.000 35.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.760 100.000 37.360 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 38.800 100.000 39.400 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.760 100.000 3.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 4.800 100.000 5.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 8.880 100.000 9.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 12.960 100.000 13.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.680 100.000 16.280 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 17.720 100.000 18.320 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.760 100.000 20.360 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 82.000 40.390 86.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END prog_clk_0_W_out
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 82.000 43.610 86.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 82.000 59.710 86.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 82.000 72.590 86.000 ;
    END
  END top_width_0_height_0__pin_11_lower
  PIN top_width_0_height_0__pin_11_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 82.000 17.850 86.000 ;
    END
  END top_width_0_height_0__pin_11_upper
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 82.000 62.930 86.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 82.000 75.810 86.000 ;
    END
  END top_width_0_height_0__pin_13_lower
  PIN top_width_0_height_0__pin_13_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 82.000 21.070 86.000 ;
    END
  END top_width_0_height_0__pin_13_upper
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 82.000 66.150 86.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 82.000 79.030 86.000 ;
    END
  END top_width_0_height_0__pin_15_lower
  PIN top_width_0_height_0__pin_15_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 82.000 24.290 86.000 ;
    END
  END top_width_0_height_0__pin_15_upper
  PIN top_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 82.000 69.370 86.000 ;
    END
  END top_width_0_height_0__pin_16_
  PIN top_width_0_height_0__pin_17_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 82.000 82.250 86.000 ;
    END
  END top_width_0_height_0__pin_17_lower
  PIN top_width_0_height_0__pin_17_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 82.000 27.510 86.000 ;
    END
  END top_width_0_height_0__pin_17_upper
  PIN top_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 82.000 85.470 86.000 ;
    END
  END top_width_0_height_0__pin_1_lower
  PIN top_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 82.000 1.750 86.000 ;
    END
  END top_width_0_height_0__pin_1_upper
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 82.000 46.830 86.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_3_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 82.000 88.690 86.000 ;
    END
  END top_width_0_height_0__pin_3_lower
  PIN top_width_0_height_0__pin_3_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 82.000 4.970 86.000 ;
    END
  END top_width_0_height_0__pin_3_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 82.000 50.050 86.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 82.000 91.910 86.000 ;
    END
  END top_width_0_height_0__pin_5_lower
  PIN top_width_0_height_0__pin_5_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 82.000 8.190 86.000 ;
    END
  END top_width_0_height_0__pin_5_upper
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 82.000 53.270 86.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 82.000 95.130 86.000 ;
    END
  END top_width_0_height_0__pin_7_lower
  PIN top_width_0_height_0__pin_7_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 82.000 11.410 86.000 ;
    END
  END top_width_0_height_0__pin_7_upper
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 82.000 56.490 86.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 82.000 98.350 86.000 ;
    END
  END top_width_0_height_0__pin_9_lower
  PIN top_width_0_height_0__pin_9_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 82.000 14.630 86.000 ;
    END
  END top_width_0_height_0__pin_9_upper
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 73.680 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 73.680 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 73.680 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.375 10.640 35.975 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.075 75.735 ;
      LAYER met1 ;
        RECT 0.990 5.480 98.370 75.780 ;
      LAYER met2 ;
        RECT 1.020 81.720 1.190 84.165 ;
        RECT 2.030 81.720 4.410 84.165 ;
        RECT 5.250 81.720 7.630 84.165 ;
        RECT 8.470 81.720 10.850 84.165 ;
        RECT 11.690 81.720 14.070 84.165 ;
        RECT 14.910 81.720 17.290 84.165 ;
        RECT 18.130 81.720 20.510 84.165 ;
        RECT 21.350 81.720 23.730 84.165 ;
        RECT 24.570 81.720 26.950 84.165 ;
        RECT 27.790 81.720 30.170 84.165 ;
        RECT 31.010 81.720 33.390 84.165 ;
        RECT 34.230 81.720 36.610 84.165 ;
        RECT 37.450 81.720 39.830 84.165 ;
        RECT 40.670 81.720 43.050 84.165 ;
        RECT 43.890 81.720 46.270 84.165 ;
        RECT 47.110 81.720 49.490 84.165 ;
        RECT 50.330 81.720 52.710 84.165 ;
        RECT 53.550 81.720 55.930 84.165 ;
        RECT 56.770 81.720 59.150 84.165 ;
        RECT 59.990 81.720 62.370 84.165 ;
        RECT 63.210 81.720 65.590 84.165 ;
        RECT 66.430 81.720 68.810 84.165 ;
        RECT 69.650 81.720 72.030 84.165 ;
        RECT 72.870 81.720 75.250 84.165 ;
        RECT 76.090 81.720 78.470 84.165 ;
        RECT 79.310 81.720 81.690 84.165 ;
        RECT 82.530 81.720 84.910 84.165 ;
        RECT 85.750 81.720 88.130 84.165 ;
        RECT 88.970 81.720 91.350 84.165 ;
        RECT 92.190 81.720 94.570 84.165 ;
        RECT 95.410 81.720 97.790 84.165 ;
        RECT 1.020 4.280 98.340 81.720 ;
        RECT 1.570 0.835 3.030 4.280 ;
        RECT 3.870 0.835 5.330 4.280 ;
        RECT 6.170 0.835 8.090 4.280 ;
        RECT 8.930 0.835 10.390 4.280 ;
        RECT 11.230 0.835 13.150 4.280 ;
        RECT 13.990 0.835 15.450 4.280 ;
        RECT 16.290 0.835 17.750 4.280 ;
        RECT 18.590 0.835 20.510 4.280 ;
        RECT 21.350 0.835 22.810 4.280 ;
        RECT 23.650 0.835 25.570 4.280 ;
        RECT 26.410 0.835 27.870 4.280 ;
        RECT 28.710 0.835 30.630 4.280 ;
        RECT 31.470 0.835 32.930 4.280 ;
        RECT 33.770 0.835 35.230 4.280 ;
        RECT 36.070 0.835 37.990 4.280 ;
        RECT 38.830 0.835 40.290 4.280 ;
        RECT 41.130 0.835 43.050 4.280 ;
        RECT 43.890 0.835 45.350 4.280 ;
        RECT 46.190 0.835 48.110 4.280 ;
        RECT 48.950 0.835 50.410 4.280 ;
        RECT 51.250 0.835 52.710 4.280 ;
        RECT 53.550 0.835 55.470 4.280 ;
        RECT 56.310 0.835 57.770 4.280 ;
        RECT 58.610 0.835 60.530 4.280 ;
        RECT 61.370 0.835 62.830 4.280 ;
        RECT 63.670 0.835 65.590 4.280 ;
        RECT 66.430 0.835 67.890 4.280 ;
        RECT 68.730 0.835 70.190 4.280 ;
        RECT 71.030 0.835 72.950 4.280 ;
        RECT 73.790 0.835 75.250 4.280 ;
        RECT 76.090 0.835 78.010 4.280 ;
        RECT 78.850 0.835 80.310 4.280 ;
        RECT 81.150 0.835 83.070 4.280 ;
        RECT 83.910 0.835 85.370 4.280 ;
        RECT 86.210 0.835 87.670 4.280 ;
        RECT 88.510 0.835 90.430 4.280 ;
        RECT 91.270 0.835 92.730 4.280 ;
        RECT 93.570 0.835 95.490 4.280 ;
        RECT 96.330 0.835 97.790 4.280 ;
      LAYER met3 ;
        RECT 4.400 83.280 95.600 84.145 ;
        RECT 4.000 82.640 96.000 83.280 ;
        RECT 4.400 81.240 95.600 82.640 ;
        RECT 4.000 80.600 96.000 81.240 ;
        RECT 4.400 79.200 95.600 80.600 ;
        RECT 4.000 78.560 96.000 79.200 ;
        RECT 4.400 77.160 95.600 78.560 ;
        RECT 4.000 76.520 96.000 77.160 ;
        RECT 4.400 75.120 95.600 76.520 ;
        RECT 4.000 74.480 96.000 75.120 ;
        RECT 4.400 73.080 95.600 74.480 ;
        RECT 4.000 72.440 96.000 73.080 ;
        RECT 4.400 71.760 96.000 72.440 ;
        RECT 4.400 71.040 95.600 71.760 ;
        RECT 4.000 70.400 95.600 71.040 ;
        RECT 4.400 70.360 95.600 70.400 ;
        RECT 4.400 69.720 96.000 70.360 ;
        RECT 4.400 69.000 95.600 69.720 ;
        RECT 4.000 68.360 95.600 69.000 ;
        RECT 4.400 68.320 95.600 68.360 ;
        RECT 4.400 67.680 96.000 68.320 ;
        RECT 4.400 66.960 95.600 67.680 ;
        RECT 4.000 66.320 95.600 66.960 ;
        RECT 4.400 66.280 95.600 66.320 ;
        RECT 4.400 65.640 96.000 66.280 ;
        RECT 4.400 64.920 95.600 65.640 ;
        RECT 4.000 64.280 95.600 64.920 ;
        RECT 4.400 64.240 95.600 64.280 ;
        RECT 4.400 63.600 96.000 64.240 ;
        RECT 4.400 62.880 95.600 63.600 ;
        RECT 4.000 62.240 95.600 62.880 ;
        RECT 4.400 62.200 95.600 62.240 ;
        RECT 4.400 61.560 96.000 62.200 ;
        RECT 4.400 60.840 95.600 61.560 ;
        RECT 4.000 60.200 95.600 60.840 ;
        RECT 4.400 60.160 95.600 60.200 ;
        RECT 4.400 59.520 96.000 60.160 ;
        RECT 4.400 58.800 95.600 59.520 ;
        RECT 4.000 58.120 95.600 58.800 ;
        RECT 4.000 57.480 96.000 58.120 ;
        RECT 4.400 56.800 96.000 57.480 ;
        RECT 4.400 56.080 95.600 56.800 ;
        RECT 4.000 55.440 95.600 56.080 ;
        RECT 4.400 55.400 95.600 55.440 ;
        RECT 4.400 54.760 96.000 55.400 ;
        RECT 4.400 54.040 95.600 54.760 ;
        RECT 4.000 53.400 95.600 54.040 ;
        RECT 4.400 53.360 95.600 53.400 ;
        RECT 4.400 52.720 96.000 53.360 ;
        RECT 4.400 52.000 95.600 52.720 ;
        RECT 4.000 51.360 95.600 52.000 ;
        RECT 4.400 51.320 95.600 51.360 ;
        RECT 4.400 50.680 96.000 51.320 ;
        RECT 4.400 49.960 95.600 50.680 ;
        RECT 4.000 49.320 95.600 49.960 ;
        RECT 4.400 49.280 95.600 49.320 ;
        RECT 4.400 48.640 96.000 49.280 ;
        RECT 4.400 47.920 95.600 48.640 ;
        RECT 4.000 47.280 95.600 47.920 ;
        RECT 4.400 47.240 95.600 47.280 ;
        RECT 4.400 46.600 96.000 47.240 ;
        RECT 4.400 45.880 95.600 46.600 ;
        RECT 4.000 45.240 95.600 45.880 ;
        RECT 4.400 45.200 95.600 45.240 ;
        RECT 4.400 44.560 96.000 45.200 ;
        RECT 4.400 43.840 95.600 44.560 ;
        RECT 4.000 43.200 95.600 43.840 ;
        RECT 4.400 43.160 95.600 43.200 ;
        RECT 4.400 41.840 96.000 43.160 ;
        RECT 4.400 41.800 95.600 41.840 ;
        RECT 4.000 41.160 95.600 41.800 ;
        RECT 4.400 40.440 95.600 41.160 ;
        RECT 4.400 39.800 96.000 40.440 ;
        RECT 4.400 39.760 95.600 39.800 ;
        RECT 4.000 39.120 95.600 39.760 ;
        RECT 4.400 38.400 95.600 39.120 ;
        RECT 4.400 37.760 96.000 38.400 ;
        RECT 4.400 37.720 95.600 37.760 ;
        RECT 4.000 37.080 95.600 37.720 ;
        RECT 4.400 36.360 95.600 37.080 ;
        RECT 4.400 35.720 96.000 36.360 ;
        RECT 4.400 35.680 95.600 35.720 ;
        RECT 4.000 35.040 95.600 35.680 ;
        RECT 4.400 34.320 95.600 35.040 ;
        RECT 4.400 33.680 96.000 34.320 ;
        RECT 4.400 33.640 95.600 33.680 ;
        RECT 4.000 33.000 95.600 33.640 ;
        RECT 4.400 32.280 95.600 33.000 ;
        RECT 4.400 31.640 96.000 32.280 ;
        RECT 4.400 31.600 95.600 31.640 ;
        RECT 4.000 30.960 95.600 31.600 ;
        RECT 4.400 30.240 95.600 30.960 ;
        RECT 4.400 29.560 96.000 30.240 ;
        RECT 4.000 28.920 96.000 29.560 ;
        RECT 4.000 28.240 95.600 28.920 ;
        RECT 4.400 27.520 95.600 28.240 ;
        RECT 4.400 26.880 96.000 27.520 ;
        RECT 4.400 26.840 95.600 26.880 ;
        RECT 4.000 26.200 95.600 26.840 ;
        RECT 4.400 25.480 95.600 26.200 ;
        RECT 4.400 24.840 96.000 25.480 ;
        RECT 4.400 24.800 95.600 24.840 ;
        RECT 4.000 24.160 95.600 24.800 ;
        RECT 4.400 23.440 95.600 24.160 ;
        RECT 4.400 22.800 96.000 23.440 ;
        RECT 4.400 22.760 95.600 22.800 ;
        RECT 4.000 22.120 95.600 22.760 ;
        RECT 4.400 21.400 95.600 22.120 ;
        RECT 4.400 20.760 96.000 21.400 ;
        RECT 4.400 20.720 95.600 20.760 ;
        RECT 4.000 20.080 95.600 20.720 ;
        RECT 4.400 19.360 95.600 20.080 ;
        RECT 4.400 18.720 96.000 19.360 ;
        RECT 4.400 18.680 95.600 18.720 ;
        RECT 4.000 18.040 95.600 18.680 ;
        RECT 4.400 17.320 95.600 18.040 ;
        RECT 4.400 16.680 96.000 17.320 ;
        RECT 4.400 16.640 95.600 16.680 ;
        RECT 4.000 16.000 95.600 16.640 ;
        RECT 4.400 15.280 95.600 16.000 ;
        RECT 4.400 14.600 96.000 15.280 ;
        RECT 4.000 13.960 96.000 14.600 ;
        RECT 4.400 12.560 95.600 13.960 ;
        RECT 4.000 11.920 96.000 12.560 ;
        RECT 4.400 10.520 95.600 11.920 ;
        RECT 4.000 9.880 96.000 10.520 ;
        RECT 4.400 8.480 95.600 9.880 ;
        RECT 4.000 7.840 96.000 8.480 ;
        RECT 4.400 6.440 95.600 7.840 ;
        RECT 4.000 5.800 96.000 6.440 ;
        RECT 4.400 4.400 95.600 5.800 ;
        RECT 4.000 3.760 96.000 4.400 ;
        RECT 4.400 2.360 95.600 3.760 ;
        RECT 4.000 1.720 96.000 2.360 ;
        RECT 4.400 0.855 95.600 1.720 ;
      LAYER met4 ;
        RECT 36.375 10.640 48.800 73.680 ;
        RECT 51.200 10.640 63.625 73.680 ;
        RECT 66.025 10.640 78.455 73.680 ;
  END
END cbx_1__0_
END LIBRARY

