magic
tech sky130A
magscale 1 2
timestamp 1679348813
<< viali >>
rect 23397 54281 23431 54315
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9597 54145 9631 54179
rect 12173 54145 12207 54179
rect 14473 54145 14507 54179
rect 15117 54145 15151 54179
rect 17049 54145 17083 54179
rect 17877 54145 17911 54179
rect 19441 54145 19475 54179
rect 19717 54145 19751 54179
rect 20729 54145 20763 54179
rect 22017 54145 22051 54179
rect 23213 54145 23247 54179
rect 24593 54145 24627 54179
rect 2513 54077 2547 54111
rect 5181 54077 5215 54111
rect 7849 54077 7883 54111
rect 9873 54077 9907 54111
rect 12633 54077 12667 54111
rect 22201 54009 22235 54043
rect 14289 53941 14323 53975
rect 14933 53941 14967 53975
rect 16865 53941 16899 53975
rect 17693 53941 17727 53975
rect 20913 53941 20947 53975
rect 24777 53941 24811 53975
rect 2053 53601 2087 53635
rect 4445 53601 4479 53635
rect 7113 53601 7147 53635
rect 11253 53601 11287 53635
rect 1777 53533 1811 53567
rect 4169 53533 4203 53567
rect 6837 53533 6871 53567
rect 10793 53533 10827 53567
rect 23121 53533 23155 53567
rect 23765 53533 23799 53567
rect 25053 53533 25087 53567
rect 23213 53397 23247 53431
rect 23949 53397 23983 53431
rect 25237 53397 25271 53431
rect 5181 53193 5215 53227
rect 5365 53057 5399 53091
rect 24317 53057 24351 53091
rect 25053 53057 25087 53091
rect 24501 52853 24535 52887
rect 25237 52853 25271 52887
rect 25329 52445 25363 52479
rect 24961 52377 24995 52411
rect 6653 52105 6687 52139
rect 6837 51969 6871 52003
rect 25329 51969 25363 52003
rect 25145 51765 25179 51799
rect 8309 51561 8343 51595
rect 9229 51493 9263 51527
rect 7849 51357 7883 51391
rect 8493 51357 8527 51391
rect 9413 51357 9447 51391
rect 7665 51289 7699 51323
rect 24961 51289 24995 51323
rect 25053 51221 25087 51255
rect 24961 50881 24995 50915
rect 25053 50677 25087 50711
rect 7849 50473 7883 50507
rect 9597 50473 9631 50507
rect 8033 50405 8067 50439
rect 7573 50269 7607 50303
rect 9505 50269 9539 50303
rect 24501 49793 24535 49827
rect 24777 49725 24811 49759
rect 10701 49317 10735 49351
rect 11713 49317 11747 49351
rect 10517 49113 10551 49147
rect 11529 49113 11563 49147
rect 25145 49113 25179 49147
rect 25237 49045 25271 49079
rect 8401 48841 8435 48875
rect 6653 48637 6687 48671
rect 6929 48637 6963 48671
rect 10368 48093 10402 48127
rect 25145 48025 25179 48059
rect 10471 47957 10505 47991
rect 25237 47957 25271 47991
rect 9873 47753 9907 47787
rect 9413 47617 9447 47651
rect 25329 47617 25363 47651
rect 9505 47413 9539 47447
rect 25145 47413 25179 47447
rect 14289 47073 14323 47107
rect 11656 47005 11690 47039
rect 11759 46937 11793 46971
rect 14473 46937 14507 46971
rect 16129 46937 16163 46971
rect 10701 46665 10735 46699
rect 12357 46597 12391 46631
rect 8309 46529 8343 46563
rect 10241 46529 10275 46563
rect 14473 46529 14507 46563
rect 25329 46529 25363 46563
rect 8125 46461 8159 46495
rect 12173 46461 12207 46495
rect 13737 46461 13771 46495
rect 14657 46461 14691 46495
rect 16313 46461 16347 46495
rect 8493 46393 8527 46427
rect 10425 46325 10459 46359
rect 25145 46325 25179 46359
rect 12679 46121 12713 46155
rect 15669 45985 15703 46019
rect 12576 45917 12610 45951
rect 13312 45917 13346 45951
rect 25329 45917 25363 45951
rect 13415 45849 13449 45883
rect 15853 45849 15887 45883
rect 17509 45849 17543 45883
rect 25145 45781 25179 45815
rect 10885 45033 10919 45067
rect 9137 44897 9171 44931
rect 25329 44829 25363 44863
rect 9413 44761 9447 44795
rect 25145 44693 25179 44727
rect 9597 44489 9631 44523
rect 9137 44353 9171 44387
rect 10609 44353 10643 44387
rect 25145 44353 25179 44387
rect 8953 44285 8987 44319
rect 25329 44217 25363 44251
rect 10701 44149 10735 44183
rect 11069 44149 11103 44183
rect 20729 43809 20763 43843
rect 20453 43741 20487 43775
rect 22201 43605 22235 43639
rect 25145 43265 25179 43299
rect 25237 43061 25271 43095
rect 9781 42721 9815 42755
rect 10241 42721 10275 42755
rect 9597 42653 9631 42687
rect 25145 42585 25179 42619
rect 25329 42585 25363 42619
rect 11161 42313 11195 42347
rect 9413 42109 9447 42143
rect 9689 42109 9723 42143
rect 10793 41769 10827 41803
rect 10333 41633 10367 41667
rect 10149 41565 10183 41599
rect 25145 41497 25179 41531
rect 25237 41429 25271 41463
rect 25329 41089 25363 41123
rect 25145 40885 25179 40919
rect 25145 40137 25179 40171
rect 25329 40001 25363 40035
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25329 38301 25363 38335
rect 25145 38165 25179 38199
rect 8677 37961 8711 37995
rect 8861 37825 8895 37859
rect 25145 37825 25179 37859
rect 25329 37689 25363 37723
rect 25145 36737 25179 36771
rect 25237 36533 25271 36567
rect 25329 36125 25363 36159
rect 25145 35989 25179 36023
rect 11161 35785 11195 35819
rect 22017 35785 22051 35819
rect 22477 35785 22511 35819
rect 21097 35717 21131 35751
rect 21189 35717 21223 35751
rect 22385 35649 22419 35683
rect 9413 35581 9447 35615
rect 9689 35581 9723 35615
rect 21281 35581 21315 35615
rect 22661 35581 22695 35615
rect 20729 35445 20763 35479
rect 23305 35105 23339 35139
rect 23121 35037 23155 35071
rect 23213 35037 23247 35071
rect 25329 35037 25363 35071
rect 22753 34901 22787 34935
rect 25145 34901 25179 34935
rect 25145 34697 25179 34731
rect 25329 34561 25363 34595
rect 9137 34153 9171 34187
rect 25145 34153 25179 34187
rect 15393 34017 15427 34051
rect 21649 34017 21683 34051
rect 9321 33949 9355 33983
rect 19441 33949 19475 33983
rect 25329 33949 25363 33983
rect 14657 33881 14691 33915
rect 19717 33881 19751 33915
rect 21925 33881 21959 33915
rect 21189 33813 21223 33847
rect 23397 33813 23431 33847
rect 19809 33541 19843 33575
rect 19533 33473 19567 33507
rect 22017 33473 22051 33507
rect 25329 33473 25363 33507
rect 22293 33405 22327 33439
rect 23765 33405 23799 33439
rect 21281 33269 21315 33303
rect 25145 33269 25179 33303
rect 24041 33065 24075 33099
rect 24593 32997 24627 33031
rect 22293 32929 22327 32963
rect 22569 32929 22603 32963
rect 25053 32929 25087 32963
rect 25145 32929 25179 32963
rect 20729 32861 20763 32895
rect 19993 32793 20027 32827
rect 24961 32793 24995 32827
rect 25237 32521 25271 32555
rect 15393 32453 15427 32487
rect 19809 32453 19843 32487
rect 22845 32453 22879 32487
rect 19533 32385 19567 32419
rect 22109 32385 22143 32419
rect 23489 32385 23523 32419
rect 16129 32317 16163 32351
rect 17325 32317 17359 32351
rect 17601 32317 17635 32351
rect 23765 32317 23799 32351
rect 19073 32181 19107 32215
rect 21281 32181 21315 32215
rect 18521 31977 18555 32011
rect 21649 31977 21683 32011
rect 15577 31909 15611 31943
rect 23029 31909 23063 31943
rect 25145 31909 25179 31943
rect 16129 31841 16163 31875
rect 16773 31841 16807 31875
rect 17049 31841 17083 31875
rect 19441 31841 19475 31875
rect 19717 31841 19751 31875
rect 22201 31841 22235 31875
rect 23581 31841 23615 31875
rect 16037 31773 16071 31807
rect 22109 31773 22143 31807
rect 23489 31773 23523 31807
rect 25329 31773 25363 31807
rect 22017 31705 22051 31739
rect 15945 31637 15979 31671
rect 21189 31637 21223 31671
rect 23397 31637 23431 31671
rect 20637 31433 20671 31467
rect 13553 31365 13587 31399
rect 20545 31365 20579 31399
rect 22661 31365 22695 31399
rect 15945 31297 15979 31331
rect 16037 31297 16071 31331
rect 17233 31297 17267 31331
rect 22385 31297 22419 31331
rect 25329 31297 25363 31331
rect 13277 31229 13311 31263
rect 16221 31229 16255 31263
rect 17325 31229 17359 31263
rect 17509 31229 17543 31263
rect 20729 31229 20763 31263
rect 16865 31161 16899 31195
rect 15025 31093 15059 31127
rect 15577 31093 15611 31127
rect 20177 31093 20211 31127
rect 24133 31093 24167 31127
rect 25145 31093 25179 31127
rect 9137 30889 9171 30923
rect 18521 30889 18555 30923
rect 22385 30889 22419 30923
rect 16773 30753 16807 30787
rect 20637 30753 20671 30787
rect 9321 30685 9355 30719
rect 14289 30685 14323 30719
rect 20177 30685 20211 30719
rect 25329 30685 25363 30719
rect 15025 30617 15059 30651
rect 17049 30617 17083 30651
rect 20913 30617 20947 30651
rect 25145 30549 25179 30583
rect 14289 30277 14323 30311
rect 20177 30277 20211 30311
rect 20269 30277 20303 30311
rect 22477 30277 22511 30311
rect 9045 30209 9079 30243
rect 11713 30209 11747 30243
rect 21465 30209 21499 30243
rect 22385 30209 22419 30243
rect 11989 30141 12023 30175
rect 15117 30141 15151 30175
rect 20453 30141 20487 30175
rect 22661 30141 22695 30175
rect 23305 30141 23339 30175
rect 23581 30141 23615 30175
rect 25053 30141 25087 30175
rect 8861 30073 8895 30107
rect 13461 30005 13495 30039
rect 19809 30005 19843 30039
rect 22017 30005 22051 30039
rect 18797 29801 18831 29835
rect 12909 29733 12943 29767
rect 20637 29733 20671 29767
rect 11161 29665 11195 29699
rect 15853 29665 15887 29699
rect 17049 29665 17083 29699
rect 19901 29665 19935 29699
rect 20085 29665 20119 29699
rect 21189 29665 21223 29699
rect 15577 29597 15611 29631
rect 25329 29597 25363 29631
rect 11437 29529 11471 29563
rect 17325 29529 17359 29563
rect 21005 29529 21039 29563
rect 21097 29529 21131 29563
rect 15209 29461 15243 29495
rect 15669 29461 15703 29495
rect 19441 29461 19475 29495
rect 19809 29461 19843 29495
rect 25145 29461 25179 29495
rect 9505 29257 9539 29291
rect 16037 29257 16071 29291
rect 19717 29257 19751 29291
rect 24041 29257 24075 29291
rect 9873 29189 9907 29223
rect 15945 29189 15979 29223
rect 23949 29189 23983 29223
rect 9965 29121 9999 29155
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 18797 29121 18831 29155
rect 19625 29121 19659 29155
rect 22201 29121 22235 29155
rect 24961 29121 24995 29155
rect 10057 29053 10091 29087
rect 15117 29053 15151 29087
rect 16129 29053 16163 29087
rect 17325 29053 17359 29087
rect 17417 29053 17451 29087
rect 19901 29053 19935 29087
rect 22937 29053 22971 29087
rect 24133 29053 24167 29087
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 19257 28985 19291 29019
rect 23581 28985 23615 29019
rect 24777 28985 24811 29019
rect 13632 28917 13666 28951
rect 10885 28713 10919 28747
rect 18889 28713 18923 28747
rect 19901 28713 19935 28747
rect 23121 28713 23155 28747
rect 15945 28645 15979 28679
rect 9137 28577 9171 28611
rect 11437 28577 11471 28611
rect 15393 28577 15427 28611
rect 16497 28577 16531 28611
rect 17417 28577 17451 28611
rect 20545 28577 20579 28611
rect 20821 28577 20855 28611
rect 23581 28577 23615 28611
rect 23765 28577 23799 28611
rect 17141 28509 17175 28543
rect 23489 28509 23523 28543
rect 24777 28509 24811 28543
rect 9413 28441 9447 28475
rect 11713 28441 11747 28475
rect 13185 28373 13219 28407
rect 14749 28373 14783 28407
rect 15117 28373 15151 28407
rect 15209 28373 15243 28407
rect 16313 28373 16347 28407
rect 16405 28373 16439 28407
rect 22293 28373 22327 28407
rect 14105 28169 14139 28203
rect 18521 28169 18555 28203
rect 24685 28169 24719 28203
rect 14013 28101 14047 28135
rect 20361 28101 20395 28135
rect 21097 28101 21131 28135
rect 17233 28033 17267 28067
rect 18429 28033 18463 28067
rect 22017 28033 22051 28067
rect 24593 28033 24627 28067
rect 14289 27965 14323 27999
rect 17325 27965 17359 27999
rect 17417 27965 17451 27999
rect 18613 27965 18647 27999
rect 22293 27965 22327 27999
rect 24777 27965 24811 27999
rect 13645 27829 13679 27863
rect 16865 27829 16899 27863
rect 18061 27829 18095 27863
rect 23765 27829 23799 27863
rect 24225 27829 24259 27863
rect 18153 27625 18187 27659
rect 20256 27625 20290 27659
rect 23581 27625 23615 27659
rect 10517 27489 10551 27523
rect 13553 27489 13587 27523
rect 15761 27489 15795 27523
rect 19993 27489 20027 27523
rect 22845 27489 22879 27523
rect 25053 27489 25087 27523
rect 25237 27489 25271 27523
rect 13461 27421 13495 27455
rect 24961 27421 24995 27455
rect 10793 27353 10827 27387
rect 13369 27353 13403 27387
rect 15577 27353 15611 27387
rect 22661 27353 22695 27387
rect 12265 27285 12299 27319
rect 13001 27285 13035 27319
rect 15209 27285 15243 27319
rect 15669 27285 15703 27319
rect 21741 27285 21775 27319
rect 22201 27285 22235 27319
rect 22569 27285 22603 27319
rect 24593 27285 24627 27319
rect 10977 27081 11011 27115
rect 15669 27081 15703 27115
rect 19717 27081 19751 27115
rect 21189 27081 21223 27115
rect 13369 27013 13403 27047
rect 15761 27013 15795 27047
rect 9229 26945 9263 26979
rect 13093 26945 13127 26979
rect 17969 26945 18003 26979
rect 21097 26945 21131 26979
rect 9505 26877 9539 26911
rect 15853 26877 15887 26911
rect 18245 26877 18279 26911
rect 21281 26877 21315 26911
rect 23305 26877 23339 26911
rect 23581 26877 23615 26911
rect 20729 26809 20763 26843
rect 14841 26741 14875 26775
rect 15301 26741 15335 26775
rect 25053 26741 25087 26775
rect 12173 26537 12207 26571
rect 21189 26537 21223 26571
rect 24593 26537 24627 26571
rect 14289 26469 14323 26503
rect 22017 26469 22051 26503
rect 22661 26469 22695 26503
rect 23857 26469 23891 26503
rect 10425 26401 10459 26435
rect 10701 26401 10735 26435
rect 14841 26401 14875 26435
rect 16037 26401 16071 26435
rect 16129 26401 16163 26435
rect 19441 26401 19475 26435
rect 19717 26401 19751 26435
rect 23213 26401 23247 26435
rect 25053 26401 25087 26435
rect 25145 26401 25179 26435
rect 18429 26333 18463 26367
rect 22201 26333 22235 26367
rect 24041 26333 24075 26367
rect 14657 26265 14691 26299
rect 23029 26265 23063 26299
rect 23121 26265 23155 26299
rect 14749 26197 14783 26231
rect 15577 26197 15611 26231
rect 15945 26197 15979 26231
rect 24961 26197 24995 26231
rect 10885 25993 10919 26027
rect 12081 25993 12115 26027
rect 12541 25993 12575 26027
rect 14013 25993 14047 26027
rect 15301 25993 15335 26027
rect 18245 25993 18279 26027
rect 22385 25993 22419 26027
rect 22477 25993 22511 26027
rect 25329 25993 25363 26027
rect 9413 25925 9447 25959
rect 18337 25925 18371 25959
rect 9137 25857 9171 25891
rect 12449 25857 12483 25891
rect 13921 25857 13955 25891
rect 15209 25857 15243 25891
rect 16221 25857 16255 25891
rect 17049 25857 17083 25891
rect 12633 25789 12667 25823
rect 14197 25789 14231 25823
rect 15393 25789 15427 25823
rect 18521 25789 18555 25823
rect 22661 25789 22695 25823
rect 23581 25789 23615 25823
rect 23857 25789 23891 25823
rect 14841 25721 14875 25755
rect 16865 25721 16899 25755
rect 13553 25653 13587 25687
rect 17877 25653 17911 25687
rect 19901 25653 19935 25687
rect 22017 25653 22051 25687
rect 10609 25449 10643 25483
rect 13737 25381 13771 25415
rect 16957 25381 16991 25415
rect 11161 25313 11195 25347
rect 11989 25313 12023 25347
rect 14841 25313 14875 25347
rect 16313 25313 16347 25347
rect 21097 25313 21131 25347
rect 10977 25245 11011 25279
rect 17141 25245 17175 25279
rect 17785 25245 17819 25279
rect 18889 25245 18923 25279
rect 19809 25245 19843 25279
rect 20913 25245 20947 25279
rect 21741 25245 21775 25279
rect 22661 25245 22695 25279
rect 25329 25245 25363 25279
rect 11069 25177 11103 25211
rect 12265 25177 12299 25211
rect 14657 25177 14691 25211
rect 16129 25177 16163 25211
rect 19993 25177 20027 25211
rect 23857 25177 23891 25211
rect 14289 25109 14323 25143
rect 14749 25109 14783 25143
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 17601 25109 17635 25143
rect 21557 25109 21591 25143
rect 25145 25109 25179 25143
rect 12081 24905 12115 24939
rect 17233 24905 17267 24939
rect 18429 24837 18463 24871
rect 22477 24837 22511 24871
rect 12173 24769 12207 24803
rect 13001 24769 13035 24803
rect 17325 24769 17359 24803
rect 18521 24769 18555 24803
rect 19717 24769 19751 24803
rect 22569 24769 22603 24803
rect 9321 24701 9355 24735
rect 9597 24701 9631 24735
rect 12265 24701 12299 24735
rect 13277 24701 13311 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19993 24701 20027 24735
rect 21465 24701 21499 24735
rect 22661 24701 22695 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 25329 24701 25363 24735
rect 11069 24565 11103 24599
rect 11713 24565 11747 24599
rect 14749 24565 14783 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 22109 24565 22143 24599
rect 11148 24361 11182 24395
rect 24777 24361 24811 24395
rect 10885 24225 10919 24259
rect 18613 24225 18647 24259
rect 18797 24225 18831 24259
rect 19441 24225 19475 24259
rect 21189 24225 21223 24259
rect 21925 24225 21959 24259
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 15945 24089 15979 24123
rect 19717 24089 19751 24123
rect 22201 24089 22235 24123
rect 12633 24021 12667 24055
rect 18153 24021 18187 24055
rect 23673 24021 23707 24055
rect 13645 23817 13679 23851
rect 14933 23817 14967 23851
rect 17233 23817 17267 23851
rect 19717 23817 19751 23851
rect 20913 23817 20947 23851
rect 21005 23817 21039 23851
rect 24961 23817 24995 23851
rect 9045 23749 9079 23783
rect 14841 23681 14875 23715
rect 18245 23681 18279 23715
rect 22385 23681 22419 23715
rect 8769 23613 8803 23647
rect 13737 23613 13771 23647
rect 13829 23613 13863 23647
rect 15025 23613 15059 23647
rect 17325 23613 17359 23647
rect 17417 23613 17451 23647
rect 19809 23613 19843 23647
rect 19993 23613 20027 23647
rect 21097 23613 21131 23647
rect 23213 23613 23247 23647
rect 23489 23613 23523 23647
rect 14473 23545 14507 23579
rect 10517 23477 10551 23511
rect 13277 23477 13311 23511
rect 15853 23477 15887 23511
rect 16865 23477 16899 23511
rect 18061 23477 18095 23511
rect 19349 23477 19383 23511
rect 20545 23477 20579 23511
rect 22201 23477 22235 23511
rect 9137 23273 9171 23307
rect 14749 23273 14783 23307
rect 20913 23273 20947 23307
rect 16037 23205 16071 23239
rect 9689 23137 9723 23171
rect 11805 23137 11839 23171
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18245 23137 18279 23171
rect 18429 23137 18463 23171
rect 20177 23137 20211 23171
rect 23489 23137 23523 23171
rect 25053 23137 25087 23171
rect 25237 23137 25271 23171
rect 11713 23069 11747 23103
rect 15117 23069 15151 23103
rect 18153 23069 18187 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 21833 23069 21867 23103
rect 22661 23069 22695 23103
rect 24961 23069 24995 23103
rect 9597 23001 9631 23035
rect 11621 23001 11655 23035
rect 9505 22933 9539 22967
rect 11253 22933 11287 22967
rect 13001 22933 13035 22967
rect 13369 22933 13403 22967
rect 13461 22933 13495 22967
rect 15209 22933 15243 22967
rect 17785 22933 17819 22967
rect 19533 22933 19567 22967
rect 21649 22933 21683 22967
rect 24593 22933 24627 22967
rect 16865 22729 16899 22763
rect 12633 22661 12667 22695
rect 21189 22661 21223 22695
rect 23305 22661 23339 22695
rect 8033 22593 8067 22627
rect 12357 22593 12391 22627
rect 17049 22593 17083 22627
rect 21097 22593 21131 22627
rect 22293 22593 22327 22627
rect 23949 22593 23983 22627
rect 8309 22525 8343 22559
rect 9781 22525 9815 22559
rect 21281 22525 21315 22559
rect 24777 22525 24811 22559
rect 14105 22389 14139 22423
rect 20177 22389 20211 22423
rect 20729 22389 20763 22423
rect 21097 22185 21131 22219
rect 23765 22185 23799 22219
rect 23305 22117 23339 22151
rect 11161 22049 11195 22083
rect 11345 22049 11379 22083
rect 12357 22049 12391 22083
rect 12449 22049 12483 22083
rect 15301 22049 15335 22083
rect 15393 22049 15427 22083
rect 16313 22049 16347 22083
rect 20177 22049 20211 22083
rect 20361 22049 20395 22083
rect 21557 22049 21591 22083
rect 25053 22049 25087 22083
rect 25145 22049 25179 22083
rect 10057 21981 10091 22015
rect 16037 21981 16071 22015
rect 20085 21981 20119 22015
rect 23949 21981 23983 22015
rect 24961 21981 24995 22015
rect 21833 21913 21867 21947
rect 10701 21845 10735 21879
rect 11069 21845 11103 21879
rect 11897 21845 11931 21879
rect 12265 21845 12299 21879
rect 14841 21845 14875 21879
rect 15209 21845 15243 21879
rect 17785 21845 17819 21879
rect 19717 21845 19751 21879
rect 24593 21845 24627 21879
rect 9781 21641 9815 21675
rect 10425 21641 10459 21675
rect 18245 21641 18279 21675
rect 19257 21641 19291 21675
rect 25053 21641 25087 21675
rect 10793 21573 10827 21607
rect 8033 21505 8067 21539
rect 11897 21505 11931 21539
rect 13093 21505 13127 21539
rect 15577 21505 15611 21539
rect 18429 21505 18463 21539
rect 19349 21505 19383 21539
rect 20269 21505 20303 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 10885 21437 10919 21471
rect 10977 21437 11011 21471
rect 13369 21437 13403 21471
rect 14841 21437 14875 21471
rect 19533 21437 19567 21471
rect 21281 21437 21315 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 23581 21437 23615 21471
rect 15761 21369 15795 21403
rect 8296 21301 8330 21335
rect 18889 21301 18923 21335
rect 22017 21301 22051 21335
rect 8585 21097 8619 21131
rect 9505 21097 9539 21131
rect 16957 21097 16991 21131
rect 20637 21029 20671 21063
rect 22201 21029 22235 21063
rect 7113 20961 7147 20995
rect 10057 20961 10091 20995
rect 12449 20961 12483 20995
rect 15209 20961 15243 20995
rect 19993 20961 20027 20995
rect 21097 20961 21131 20995
rect 21189 20961 21223 20995
rect 25145 20961 25179 20995
rect 6837 20893 6871 20927
rect 9873 20893 9907 20927
rect 10701 20893 10735 20927
rect 19809 20893 19843 20927
rect 19901 20893 19935 20927
rect 21005 20893 21039 20927
rect 22661 20893 22695 20927
rect 25053 20893 25087 20927
rect 10977 20825 11011 20859
rect 15485 20825 15519 20859
rect 23857 20825 23891 20859
rect 9965 20757 9999 20791
rect 19441 20757 19475 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 15485 20553 15519 20587
rect 22109 20553 22143 20587
rect 25329 20553 25363 20587
rect 10885 20485 10919 20519
rect 17141 20485 17175 20519
rect 7757 20417 7791 20451
rect 12725 20417 12759 20451
rect 15393 20417 15427 20451
rect 16865 20417 16899 20451
rect 19257 20417 19291 20451
rect 20085 20417 20119 20451
rect 22293 20417 22327 20451
rect 22937 20417 22971 20451
rect 8033 20349 8067 20383
rect 9781 20349 9815 20383
rect 10977 20349 11011 20383
rect 13001 20349 13035 20383
rect 15577 20349 15611 20383
rect 18613 20349 18647 20383
rect 21281 20349 21315 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 14473 20213 14507 20247
rect 15025 20213 15059 20247
rect 19073 20213 19107 20247
rect 22753 20213 22787 20247
rect 9394 20009 9428 20043
rect 11345 20009 11379 20043
rect 16037 20009 16071 20043
rect 16497 20009 16531 20043
rect 23857 20009 23891 20043
rect 9137 19873 9171 19907
rect 11989 19873 12023 19907
rect 14289 19873 14323 19907
rect 18061 19873 18095 19907
rect 19901 19873 19935 19907
rect 22109 19873 22143 19907
rect 16681 19805 16715 19839
rect 17969 19805 18003 19839
rect 18889 19805 18923 19839
rect 14565 19737 14599 19771
rect 20177 19737 20211 19771
rect 22385 19737 22419 19771
rect 10885 19669 10919 19703
rect 11713 19669 11747 19703
rect 11805 19669 11839 19703
rect 17509 19669 17543 19703
rect 17877 19669 17911 19703
rect 18705 19669 18739 19703
rect 21649 19669 21683 19703
rect 8769 19465 8803 19499
rect 14197 19465 14231 19499
rect 14933 19465 14967 19499
rect 15577 19465 15611 19499
rect 17049 19465 17083 19499
rect 17509 19465 17543 19499
rect 18981 19465 19015 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22201 19465 22235 19499
rect 22661 19465 22695 19499
rect 25145 19465 25179 19499
rect 15945 19397 15979 19431
rect 16037 19397 16071 19431
rect 17417 19397 17451 19431
rect 23673 19397 23707 19431
rect 9137 19329 9171 19363
rect 9229 19329 9263 19363
rect 11897 19329 11931 19363
rect 12449 19329 12483 19363
rect 15117 19329 15151 19363
rect 19165 19329 19199 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 12725 19261 12759 19295
rect 16129 19261 16163 19295
rect 17601 19261 17635 19295
rect 20637 19261 20671 19295
rect 21465 19261 21499 19295
rect 22753 19261 22787 19295
rect 8309 19125 8343 19159
rect 20085 19125 20119 19159
rect 8401 18921 8435 18955
rect 10057 18921 10091 18955
rect 11529 18921 11563 18955
rect 21649 18921 21683 18955
rect 20269 18853 20303 18887
rect 6929 18785 6963 18819
rect 10609 18785 10643 18819
rect 12081 18785 12115 18819
rect 17233 18785 17267 18819
rect 17417 18785 17451 18819
rect 23857 18785 23891 18819
rect 6653 18717 6687 18751
rect 10425 18717 10459 18751
rect 12909 18717 12943 18751
rect 16221 18717 16255 18751
rect 17141 18717 17175 18751
rect 19625 18717 19659 18751
rect 20453 18717 20487 18751
rect 21097 18717 21131 18751
rect 21833 18717 21867 18751
rect 22661 18717 22695 18751
rect 24777 18717 24811 18751
rect 11897 18649 11931 18683
rect 11989 18649 12023 18683
rect 10517 18581 10551 18615
rect 16037 18581 16071 18615
rect 16773 18581 16807 18615
rect 19441 18581 19475 18615
rect 20913 18581 20947 18615
rect 24593 18581 24627 18615
rect 9413 18377 9447 18411
rect 10333 18377 10367 18411
rect 13737 18377 13771 18411
rect 14105 18377 14139 18411
rect 13277 18309 13311 18343
rect 22661 18309 22695 18343
rect 23581 18309 23615 18343
rect 10241 18241 10275 18275
rect 16865 18241 16899 18275
rect 20545 18241 20579 18275
rect 21189 18241 21223 18275
rect 23305 18241 23339 18275
rect 7665 18173 7699 18207
rect 7941 18173 7975 18207
rect 10425 18173 10459 18207
rect 14197 18173 14231 18207
rect 14289 18173 14323 18207
rect 17141 18173 17175 18207
rect 25329 18173 25363 18207
rect 9873 18105 9907 18139
rect 20361 18105 20395 18139
rect 18613 18037 18647 18071
rect 21005 18037 21039 18071
rect 22753 18037 22787 18071
rect 7849 17833 7883 17867
rect 21189 17833 21223 17867
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 11805 17697 11839 17731
rect 13093 17697 13127 17731
rect 18429 17697 18463 17731
rect 18613 17697 18647 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 7389 17629 7423 17663
rect 9321 17629 9355 17663
rect 9781 17629 9815 17663
rect 12357 17629 12391 17663
rect 13645 17629 13679 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 19441 17629 19475 17663
rect 22017 17629 22051 17663
rect 22661 17629 22695 17663
rect 8217 17561 8251 17595
rect 18337 17561 18371 17595
rect 19717 17561 19751 17595
rect 8309 17493 8343 17527
rect 16681 17493 16715 17527
rect 17969 17493 18003 17527
rect 22109 17493 22143 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 12357 17289 12391 17323
rect 13185 17289 13219 17323
rect 18889 17289 18923 17323
rect 21189 17289 21223 17323
rect 10977 17221 11011 17255
rect 16957 17221 16991 17255
rect 18245 17221 18279 17255
rect 23305 17221 23339 17255
rect 10241 17153 10275 17187
rect 12449 17153 12483 17187
rect 13277 17153 13311 17187
rect 14473 17153 14507 17187
rect 19073 17153 19107 17187
rect 19993 17153 20027 17187
rect 21097 17153 21131 17187
rect 22201 17153 22235 17187
rect 24133 17153 24167 17187
rect 8125 17085 8159 17119
rect 8309 17085 8343 17119
rect 9505 17085 9539 17119
rect 9597 17085 9631 17119
rect 12541 17085 12575 17119
rect 13369 17085 13403 17119
rect 14749 17085 14783 17119
rect 21373 17085 21407 17119
rect 24777 17085 24811 17119
rect 7665 17017 7699 17051
rect 11989 17017 12023 17051
rect 16221 17017 16255 17051
rect 17141 17017 17175 17051
rect 19809 17017 19843 17051
rect 12817 16949 12851 16983
rect 18337 16949 18371 16983
rect 20729 16949 20763 16983
rect 24777 16745 24811 16779
rect 10977 16609 11011 16643
rect 11805 16609 11839 16643
rect 12081 16609 12115 16643
rect 15117 16609 15151 16643
rect 16221 16609 16255 16643
rect 16313 16609 16347 16643
rect 18337 16609 18371 16643
rect 20269 16609 20303 16643
rect 16129 16541 16163 16575
rect 21005 16541 21039 16575
rect 21649 16541 21683 16575
rect 22661 16541 22695 16575
rect 10793 16473 10827 16507
rect 15025 16473 15059 16507
rect 17509 16473 17543 16507
rect 19441 16473 19475 16507
rect 23857 16473 23891 16507
rect 10425 16405 10459 16439
rect 10885 16405 10919 16439
rect 13553 16405 13587 16439
rect 14565 16405 14599 16439
rect 14933 16405 14967 16439
rect 15761 16405 15795 16439
rect 20821 16405 20855 16439
rect 21465 16405 21499 16439
rect 10241 16201 10275 16235
rect 12173 16201 12207 16235
rect 12541 16201 12575 16235
rect 14565 16201 14599 16235
rect 15025 16201 15059 16235
rect 10701 16133 10735 16167
rect 17233 16133 17267 16167
rect 6561 16065 6595 16099
rect 10609 16065 10643 16099
rect 12633 16065 12667 16099
rect 13737 16065 13771 16099
rect 14933 16065 14967 16099
rect 15945 16065 15979 16099
rect 18061 16065 18095 16099
rect 18705 16065 18739 16099
rect 19717 16065 19751 16099
rect 24409 16065 24443 16099
rect 25053 16065 25087 16099
rect 6837 15997 6871 16031
rect 10793 15997 10827 16031
rect 12725 15997 12759 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 15117 15997 15151 16031
rect 19993 15997 20027 16031
rect 22017 15997 22051 16031
rect 22293 15997 22327 16031
rect 13369 15929 13403 15963
rect 8309 15861 8343 15895
rect 17325 15861 17359 15895
rect 17877 15861 17911 15895
rect 18521 15861 18555 15895
rect 21465 15861 21499 15895
rect 23765 15861 23799 15895
rect 24869 15861 24903 15895
rect 9137 15657 9171 15691
rect 11713 15657 11747 15691
rect 16576 15657 16610 15691
rect 9689 15521 9723 15555
rect 12265 15521 12299 15555
rect 16313 15521 16347 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 24041 15521 24075 15555
rect 14473 15453 14507 15487
rect 15853 15453 15887 15487
rect 21833 15453 21867 15487
rect 24777 15453 24811 15487
rect 12081 15385 12115 15419
rect 19717 15385 19751 15419
rect 9505 15317 9539 15351
rect 9597 15317 9631 15351
rect 12173 15317 12207 15351
rect 18061 15317 18095 15351
rect 21189 15317 21223 15351
rect 21649 15317 21683 15351
rect 24593 15317 24627 15351
rect 10149 15113 10183 15147
rect 13645 15113 13679 15147
rect 14013 15113 14047 15147
rect 15945 15113 15979 15147
rect 19993 15113 20027 15147
rect 21189 15113 21223 15147
rect 22293 15113 22327 15147
rect 10517 15045 10551 15079
rect 18705 15045 18739 15079
rect 10609 14977 10643 15011
rect 19901 14977 19935 15011
rect 21097 14977 21131 15011
rect 22477 14977 22511 15011
rect 23949 14977 23983 15011
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9689 14909 9723 14943
rect 10701 14909 10735 14943
rect 14105 14909 14139 14943
rect 14289 14909 14323 14943
rect 16037 14909 16071 14943
rect 16221 14909 16255 14943
rect 20085 14909 20119 14943
rect 21373 14909 21407 14943
rect 24777 14909 24811 14943
rect 15577 14841 15611 14875
rect 19533 14841 19567 14875
rect 18797 14773 18831 14807
rect 20729 14773 20763 14807
rect 8125 14569 8159 14603
rect 6377 14433 6411 14467
rect 6653 14433 6687 14467
rect 11989 14433 12023 14467
rect 13645 14433 13679 14467
rect 16957 14433 16991 14467
rect 22293 14433 22327 14467
rect 9965 14365 9999 14399
rect 12541 14365 12575 14399
rect 13369 14365 13403 14399
rect 16773 14365 16807 14399
rect 17785 14365 17819 14399
rect 20453 14365 20487 14399
rect 24777 14365 24811 14399
rect 10241 14297 10275 14331
rect 22569 14297 22603 14331
rect 13001 14229 13035 14263
rect 13461 14229 13495 14263
rect 16405 14229 16439 14263
rect 16865 14229 16899 14263
rect 20269 14229 20303 14263
rect 24041 14229 24075 14263
rect 24593 14229 24627 14263
rect 13001 14025 13035 14059
rect 18613 14025 18647 14059
rect 20177 14025 20211 14059
rect 8033 13957 8067 13991
rect 9781 13957 9815 13991
rect 10977 13957 11011 13991
rect 19533 13957 19567 13991
rect 25145 13957 25179 13991
rect 10241 13889 10275 13923
rect 20361 13889 20395 13923
rect 21097 13889 21131 13923
rect 22293 13889 22327 13923
rect 24133 13889 24167 13923
rect 7757 13821 7791 13855
rect 13093 13821 13127 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 15577 13821 15611 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 19717 13821 19751 13855
rect 23305 13821 23339 13855
rect 20913 13753 20947 13787
rect 11897 13685 11931 13719
rect 12633 13685 12667 13719
rect 14092 13685 14126 13719
rect 8217 13481 8251 13515
rect 9229 13481 9263 13515
rect 13001 13481 13035 13515
rect 6469 13345 6503 13379
rect 9689 13345 9723 13379
rect 9781 13345 9815 13379
rect 10425 13345 10459 13379
rect 13553 13345 13587 13379
rect 15761 13345 15795 13379
rect 21281 13345 21315 13379
rect 21465 13345 21499 13379
rect 15577 13277 15611 13311
rect 19441 13277 19475 13311
rect 21189 13277 21223 13311
rect 22201 13277 22235 13311
rect 22845 13277 22879 13311
rect 24777 13277 24811 13311
rect 6745 13209 6779 13243
rect 9597 13209 9631 13243
rect 10701 13209 10735 13243
rect 13369 13209 13403 13243
rect 17877 13209 17911 13243
rect 18061 13209 18095 13243
rect 18613 13209 18647 13243
rect 20269 13209 20303 13243
rect 23857 13209 23891 13243
rect 12173 13141 12207 13175
rect 13461 13141 13495 13175
rect 15209 13141 15243 13175
rect 15669 13141 15703 13175
rect 18705 13141 18739 13175
rect 20821 13141 20855 13175
rect 24593 13141 24627 13175
rect 6653 12937 6687 12971
rect 7849 12937 7883 12971
rect 9045 12937 9079 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 13737 12937 13771 12971
rect 15301 12937 15335 12971
rect 17325 12937 17359 12971
rect 18061 12937 18095 12971
rect 18705 12937 18739 12971
rect 19073 12937 19107 12971
rect 21189 12937 21223 12971
rect 22017 12937 22051 12971
rect 8217 12869 8251 12903
rect 10885 12869 10919 12903
rect 11897 12869 11931 12903
rect 12725 12869 12759 12903
rect 15393 12869 15427 12903
rect 23305 12869 23339 12903
rect 7021 12801 7055 12835
rect 9413 12801 9447 12835
rect 14105 12801 14139 12835
rect 17233 12801 17267 12835
rect 18245 12801 18279 12835
rect 20085 12801 20119 12835
rect 21097 12801 21131 12835
rect 22201 12801 22235 12835
rect 7113 12733 7147 12767
rect 7205 12733 7239 12767
rect 8309 12733 8343 12767
rect 8401 12733 8435 12767
rect 9505 12733 9539 12767
rect 9689 12733 9723 12767
rect 10977 12733 11011 12767
rect 14197 12733 14231 12767
rect 14289 12733 14323 12767
rect 15485 12733 15519 12767
rect 17509 12733 17543 12767
rect 19165 12733 19199 12767
rect 19349 12733 19383 12767
rect 21373 12733 21407 12767
rect 23029 12733 23063 12767
rect 19901 12665 19935 12699
rect 20729 12665 20763 12699
rect 14933 12597 14967 12631
rect 16865 12597 16899 12631
rect 24777 12597 24811 12631
rect 7573 12393 7607 12427
rect 8401 12393 8435 12427
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 14381 12393 14415 12427
rect 10793 12257 10827 12291
rect 12081 12257 12115 12291
rect 13277 12257 13311 12291
rect 14933 12257 14967 12291
rect 20361 12257 20395 12291
rect 13001 12189 13035 12223
rect 17233 12189 17267 12223
rect 18705 12189 18739 12223
rect 19533 12189 19567 12223
rect 22845 12189 22879 12223
rect 24777 12189 24811 12223
rect 11805 12121 11839 12155
rect 13093 12121 13127 12155
rect 14841 12121 14875 12155
rect 17969 12121 18003 12155
rect 18889 12121 18923 12155
rect 20637 12121 20671 12155
rect 23857 12121 23891 12155
rect 10609 12053 10643 12087
rect 10701 12053 10735 12087
rect 11897 12053 11931 12087
rect 14749 12053 14783 12087
rect 19625 12053 19659 12087
rect 22109 12053 22143 12087
rect 24593 12053 24627 12087
rect 9045 11849 9079 11883
rect 9781 11849 9815 11883
rect 11989 11849 12023 11883
rect 12357 11849 12391 11883
rect 13185 11849 13219 11883
rect 13645 11849 13679 11883
rect 14381 11849 14415 11883
rect 14749 11849 14783 11883
rect 17325 11849 17359 11883
rect 18061 11849 18095 11883
rect 19625 11849 19659 11883
rect 10241 11781 10275 11815
rect 20913 11781 20947 11815
rect 22385 11781 22419 11815
rect 23397 11781 23431 11815
rect 10149 11713 10183 11747
rect 12449 11713 12483 11747
rect 13553 11713 13587 11747
rect 17233 11713 17267 11747
rect 18429 11713 18463 11747
rect 19993 11713 20027 11747
rect 22201 11713 22235 11747
rect 23121 11713 23155 11747
rect 7297 11645 7331 11679
rect 7573 11645 7607 11679
rect 10333 11645 10367 11679
rect 12541 11645 12575 11679
rect 13737 11645 13771 11679
rect 14841 11645 14875 11679
rect 14933 11645 14967 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 20085 11645 20119 11679
rect 20269 11645 20303 11679
rect 16865 11577 16899 11611
rect 21005 11509 21039 11543
rect 24869 11509 24903 11543
rect 12633 11305 12667 11339
rect 17233 11305 17267 11339
rect 19625 11305 19659 11339
rect 21649 11305 21683 11339
rect 22109 11305 22143 11339
rect 24593 11305 24627 11339
rect 16497 11237 16531 11271
rect 17877 11237 17911 11271
rect 20821 11237 20855 11271
rect 9413 11169 9447 11203
rect 11989 11169 12023 11203
rect 13277 11169 13311 11203
rect 14749 11169 14783 11203
rect 18337 11169 18371 11203
rect 18521 11169 18555 11203
rect 23581 11169 23615 11203
rect 9137 11101 9171 11135
rect 13001 11101 13035 11135
rect 17417 11101 17451 11135
rect 20177 11101 20211 11135
rect 21005 11101 21039 11135
rect 22293 11101 22327 11135
rect 22937 11101 22971 11135
rect 24777 11101 24811 11135
rect 11805 11033 11839 11067
rect 11897 11033 11931 11067
rect 13093 11033 13127 11067
rect 15025 11033 15059 11067
rect 18245 11033 18279 11067
rect 20361 11033 20395 11067
rect 10885 10965 10919 10999
rect 11437 10965 11471 10999
rect 22753 10965 22787 10999
rect 9965 10761 9999 10795
rect 12541 10761 12575 10795
rect 13737 10761 13771 10795
rect 15577 10761 15611 10795
rect 8493 10693 8527 10727
rect 13001 10693 13035 10727
rect 14105 10693 14139 10727
rect 15945 10693 15979 10727
rect 19993 10693 20027 10727
rect 23213 10693 23247 10727
rect 12909 10625 12943 10659
rect 17509 10625 17543 10659
rect 18705 10625 18739 10659
rect 22201 10625 22235 10659
rect 23121 10625 23155 10659
rect 24133 10625 24167 10659
rect 8217 10557 8251 10591
rect 13185 10557 13219 10591
rect 14197 10557 14231 10591
rect 14381 10557 14415 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 18429 10557 18463 10591
rect 19717 10557 19751 10591
rect 21465 10557 21499 10591
rect 23397 10557 23431 10591
rect 24777 10557 24811 10591
rect 11161 10421 11195 10455
rect 12081 10421 12115 10455
rect 17601 10421 17635 10455
rect 22017 10421 22051 10455
rect 22753 10421 22787 10455
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 14565 10217 14599 10251
rect 24593 10217 24627 10251
rect 12817 10149 12851 10183
rect 18153 10149 18187 10183
rect 9321 10081 9355 10115
rect 12081 10081 12115 10115
rect 12173 10081 12207 10115
rect 13277 10081 13311 10115
rect 13461 10081 13495 10115
rect 15117 10081 15151 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 21373 10081 21407 10115
rect 21465 10081 21499 10115
rect 22293 10081 22327 10115
rect 22569 10081 22603 10115
rect 11989 10013 12023 10047
rect 17693 10013 17727 10047
rect 20269 10013 20303 10047
rect 21281 10013 21315 10047
rect 24777 10013 24811 10047
rect 9597 9945 9631 9979
rect 13185 9945 13219 9979
rect 15025 9945 15059 9979
rect 16865 9945 16899 9979
rect 19533 9945 19567 9979
rect 14933 9877 14967 9911
rect 16957 9877 16991 9911
rect 17509 9877 17543 9911
rect 18521 9877 18555 9911
rect 19625 9877 19659 9911
rect 20361 9877 20395 9911
rect 20913 9877 20947 9911
rect 24041 9877 24075 9911
rect 14381 9605 14415 9639
rect 15669 9605 15703 9639
rect 15577 9537 15611 9571
rect 17233 9537 17267 9571
rect 20269 9537 20303 9571
rect 22293 9537 22327 9571
rect 24133 9537 24167 9571
rect 11713 9469 11747 9503
rect 11989 9469 12023 9503
rect 13461 9469 13495 9503
rect 14473 9469 14507 9503
rect 14657 9469 14691 9503
rect 15761 9469 15795 9503
rect 17693 9469 17727 9503
rect 17969 9469 18003 9503
rect 20361 9469 20395 9503
rect 20545 9469 20579 9503
rect 23305 9469 23339 9503
rect 24685 9469 24719 9503
rect 15209 9401 15243 9435
rect 14013 9333 14047 9367
rect 19441 9333 19475 9367
rect 19901 9333 19935 9367
rect 21281 9333 21315 9367
rect 11621 9129 11655 9163
rect 13001 9061 13035 9095
rect 17141 9061 17175 9095
rect 18705 9061 18739 9095
rect 9137 8993 9171 9027
rect 12173 8993 12207 9027
rect 13461 8993 13495 9027
rect 13553 8993 13587 9027
rect 14933 8993 14967 9027
rect 16497 8993 16531 9027
rect 17601 8993 17635 9027
rect 17693 8993 17727 9027
rect 20085 8993 20119 9027
rect 20177 8993 20211 9027
rect 11989 8925 12023 8959
rect 16313 8925 16347 8959
rect 18889 8921 18923 8955
rect 19993 8925 20027 8959
rect 20821 8925 20855 8959
rect 22661 8925 22695 8959
rect 24777 8925 24811 8959
rect 9413 8857 9447 8891
rect 12081 8857 12115 8891
rect 14749 8857 14783 8891
rect 21833 8857 21867 8891
rect 23857 8857 23891 8891
rect 10885 8789 10919 8823
rect 13369 8789 13403 8823
rect 14289 8789 14323 8823
rect 14657 8789 14691 8823
rect 15945 8789 15979 8823
rect 16405 8789 16439 8823
rect 17509 8789 17543 8823
rect 19625 8789 19659 8823
rect 24593 8789 24627 8823
rect 11713 8585 11747 8619
rect 16865 8585 16899 8619
rect 18889 8585 18923 8619
rect 21465 8585 21499 8619
rect 13921 8517 13955 8551
rect 11161 8449 11195 8483
rect 12081 8449 12115 8483
rect 14841 8449 14875 8483
rect 15117 8449 15151 8483
rect 17233 8449 17267 8483
rect 18797 8449 18831 8483
rect 19717 8449 19751 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 12173 8381 12207 8415
rect 12357 8381 12391 8415
rect 17325 8381 17359 8415
rect 17417 8381 17451 8415
rect 18981 8381 19015 8415
rect 22569 8381 22603 8415
rect 24777 8381 24811 8415
rect 14105 8313 14139 8347
rect 16313 8313 16347 8347
rect 13369 8245 13403 8279
rect 18429 8245 18463 8279
rect 19980 8245 20014 8279
rect 11805 8041 11839 8075
rect 14289 8041 14323 8075
rect 16773 8041 16807 8075
rect 24685 8041 24719 8075
rect 10333 7973 10367 8007
rect 18153 7973 18187 8007
rect 10885 7905 10919 7939
rect 12357 7905 12391 7939
rect 13645 7905 13679 7939
rect 14841 7905 14875 7939
rect 15485 7905 15519 7939
rect 17325 7905 17359 7939
rect 18797 7905 18831 7939
rect 22293 7905 22327 7939
rect 22569 7905 22603 7939
rect 10793 7837 10827 7871
rect 13369 7837 13403 7871
rect 14657 7837 14691 7871
rect 15761 7837 15795 7871
rect 17141 7837 17175 7871
rect 20637 7837 20671 7871
rect 24869 7837 24903 7871
rect 12173 7769 12207 7803
rect 13461 7769 13495 7803
rect 18521 7769 18555 7803
rect 19533 7769 19567 7803
rect 19717 7769 19751 7803
rect 21649 7769 21683 7803
rect 10701 7701 10735 7735
rect 12265 7701 12299 7735
rect 13001 7701 13035 7735
rect 14749 7701 14783 7735
rect 17233 7701 17267 7735
rect 18613 7701 18647 7735
rect 24041 7701 24075 7735
rect 10701 7497 10735 7531
rect 11713 7497 11747 7531
rect 12081 7429 12115 7463
rect 12173 7429 12207 7463
rect 16129 7429 16163 7463
rect 17049 7429 17083 7463
rect 25145 7429 25179 7463
rect 13277 7361 13311 7395
rect 20085 7361 20119 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 8953 7293 8987 7327
rect 9229 7293 9263 7327
rect 12265 7293 12299 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 17693 7293 17727 7327
rect 17969 7293 18003 7327
rect 19441 7293 19475 7327
rect 21281 7293 21315 7327
rect 23305 7293 23339 7327
rect 17233 7225 17267 7259
rect 15485 7157 15519 7191
rect 16221 7157 16255 7191
rect 20164 6953 20198 6987
rect 22372 6953 22406 6987
rect 11069 6817 11103 6851
rect 12541 6817 12575 6851
rect 13645 6817 13679 6851
rect 15577 6817 15611 6851
rect 16957 6817 16991 6851
rect 19901 6817 19935 6851
rect 22098 6817 22132 6851
rect 25145 6817 25179 6851
rect 10793 6749 10827 6783
rect 13461 6749 13495 6783
rect 14565 6749 14599 6783
rect 17693 6749 17727 6783
rect 13369 6681 13403 6715
rect 16773 6681 16807 6715
rect 18705 6681 18739 6715
rect 25053 6681 25087 6715
rect 13001 6613 13035 6647
rect 14381 6613 14415 6647
rect 15025 6613 15059 6647
rect 15393 6613 15427 6647
rect 15485 6613 15519 6647
rect 16313 6613 16347 6647
rect 16681 6613 16715 6647
rect 21649 6613 21683 6647
rect 23857 6613 23891 6647
rect 24593 6613 24627 6647
rect 24961 6613 24995 6647
rect 15301 6409 15335 6443
rect 18613 6409 18647 6443
rect 15761 6341 15795 6375
rect 21281 6341 21315 6375
rect 25145 6341 25179 6375
rect 13001 6273 13035 6307
rect 13737 6273 13771 6307
rect 15669 6273 15703 6307
rect 19257 6273 19291 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 24133 6273 24167 6307
rect 13461 6205 13495 6239
rect 15853 6205 15887 6239
rect 16865 6205 16899 6239
rect 17141 6205 17175 6239
rect 22477 6205 22511 6239
rect 19073 6069 19107 6103
rect 11713 5865 11747 5899
rect 24685 5865 24719 5899
rect 10241 5729 10275 5763
rect 16773 5729 16807 5763
rect 22661 5729 22695 5763
rect 9965 5661 9999 5695
rect 13737 5661 13771 5695
rect 14473 5661 14507 5695
rect 15025 5661 15059 5695
rect 15853 5661 15887 5695
rect 17693 5661 17727 5695
rect 18705 5661 18739 5695
rect 20361 5661 20395 5695
rect 22201 5661 22235 5695
rect 24869 5661 24903 5695
rect 15209 5593 15243 5627
rect 19533 5593 19567 5627
rect 19717 5593 19751 5627
rect 21281 5593 21315 5627
rect 13553 5525 13587 5559
rect 14289 5525 14323 5559
rect 14841 5321 14875 5355
rect 13369 5253 13403 5287
rect 17141 5253 17175 5287
rect 15485 5185 15519 5219
rect 19257 5185 19291 5219
rect 19717 5185 19751 5219
rect 22109 5185 22143 5219
rect 24133 5185 24167 5219
rect 13093 5117 13127 5151
rect 15761 5117 15795 5151
rect 16865 5117 16899 5151
rect 18613 5117 18647 5151
rect 19993 5117 20027 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 21465 5049 21499 5083
rect 14749 4777 14783 4811
rect 16957 4777 16991 4811
rect 23305 4777 23339 4811
rect 23857 4709 23891 4743
rect 24869 4709 24903 4743
rect 5089 4641 5123 4675
rect 13185 4641 13219 4675
rect 15209 4641 15243 4675
rect 17877 4641 17911 4675
rect 19901 4641 19935 4675
rect 7113 4573 7147 4607
rect 12449 4573 12483 4607
rect 12909 4573 12943 4607
rect 17601 4573 17635 4607
rect 19625 4573 19659 4607
rect 21465 4573 21499 4607
rect 23213 4573 23247 4607
rect 24041 4573 24075 4607
rect 24685 4573 24719 4607
rect 5365 4505 5399 4539
rect 15485 4505 15519 4539
rect 22201 4505 22235 4539
rect 15669 4233 15703 4267
rect 20913 4165 20947 4199
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 4353 4097 4387 4131
rect 6745 4097 6779 4131
rect 12265 4097 12299 4131
rect 13921 4097 13955 4131
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 18705 4097 18739 4131
rect 21005 4097 21039 4131
rect 22109 4097 22143 4131
rect 23857 4097 23891 4131
rect 13277 4029 13311 4063
rect 14197 4029 14231 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 21189 4029 21223 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 2237 3961 2271 3995
rect 4169 3961 4203 3995
rect 6561 3961 6595 3995
rect 16129 3961 16163 3995
rect 1593 3893 1627 3927
rect 20545 3893 20579 3927
rect 2881 3689 2915 3723
rect 4261 3689 4295 3723
rect 6745 3689 6779 3723
rect 8217 3689 8251 3723
rect 9689 3689 9723 3723
rect 17969 3689 18003 3723
rect 10425 3621 10459 3655
rect 1869 3553 1903 3587
rect 5181 3553 5215 3587
rect 11069 3553 11103 3587
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 19993 3553 20027 3587
rect 21741 3553 21775 3587
rect 23489 3553 23523 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 6929 3485 6963 3519
rect 8401 3485 8435 3519
rect 9873 3485 9907 3519
rect 10609 3485 10643 3519
rect 11345 3485 11379 3519
rect 12449 3485 12483 3519
rect 14473 3485 14507 3519
rect 16313 3485 16347 3519
rect 18153 3485 18187 3519
rect 18889 3485 18923 3519
rect 19625 3485 19659 3519
rect 21281 3485 21315 3519
rect 23213 3485 23247 3519
rect 24685 3485 24719 3519
rect 18705 3417 18739 3451
rect 24869 3417 24903 3451
rect 7113 3145 7147 3179
rect 8401 3145 8435 3179
rect 10977 3145 11011 3179
rect 20637 3145 20671 3179
rect 21281 3145 21315 3179
rect 24869 3145 24903 3179
rect 22109 3077 22143 3111
rect 22293 3077 22327 3111
rect 2145 3009 2179 3043
rect 3709 3009 3743 3043
rect 7297 3009 7331 3043
rect 7941 3009 7975 3043
rect 8585 3009 8619 3043
rect 9229 3009 9263 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 11161 3009 11195 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 14841 3009 14875 3043
rect 17049 3009 17083 3043
rect 18705 3009 18739 3043
rect 20821 3009 20855 3043
rect 21465 3009 21499 3043
rect 22937 3009 22971 3043
rect 23581 3009 23615 3043
rect 2421 2941 2455 2975
rect 3433 2941 3467 2975
rect 5181 2941 5215 2975
rect 5457 2941 5491 2975
rect 11713 2941 11747 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 7757 2873 7791 2907
rect 10333 2873 10367 2907
rect 22753 2873 22787 2907
rect 9045 2805 9079 2839
rect 9689 2805 9723 2839
rect 2835 2601 2869 2635
rect 7113 2601 7147 2635
rect 9137 2601 9171 2635
rect 11713 2601 11747 2635
rect 18705 2601 18739 2635
rect 21465 2601 21499 2635
rect 24777 2601 24811 2635
rect 2605 2465 2639 2499
rect 5181 2465 5215 2499
rect 8033 2465 8067 2499
rect 14933 2465 14967 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 4721 2397 4755 2431
rect 5457 2397 5491 2431
rect 7297 2397 7331 2431
rect 7757 2397 7791 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14473 2397 14507 2431
rect 16865 2397 16899 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 24041 2397 24075 2431
rect 10977 2329 11011 2363
rect 13277 2329 13311 2363
rect 4537 2261 4571 2295
rect 23857 2261 23891 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 18598 54272 18604 54324
rect 18656 54312 18662 54324
rect 23385 54315 23443 54321
rect 23385 54312 23397 54315
rect 18656 54284 23397 54312
rect 18656 54272 18662 54284
rect 23385 54281 23397 54284
rect 23431 54281 23443 54315
rect 23385 54275 23443 54281
rect 8570 54204 8576 54256
rect 8628 54244 8634 54256
rect 8628 54216 19748 54244
rect 8628 54204 8634 54216
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4062 54176 4068 54188
rect 2271 54148 4068 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4062 54136 4068 54148
rect 4120 54136 4126 54188
rect 4798 54136 4804 54188
rect 4856 54136 4862 54188
rect 7374 54136 7380 54188
rect 7432 54136 7438 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 11698 54136 11704 54188
rect 11756 54176 11762 54188
rect 12161 54179 12219 54185
rect 12161 54176 12173 54179
rect 11756 54148 12173 54176
rect 11756 54136 11762 54148
rect 12161 54145 12173 54148
rect 12207 54145 12219 54179
rect 12161 54139 12219 54145
rect 13722 54136 13728 54188
rect 13780 54176 13786 54188
rect 14461 54179 14519 54185
rect 14461 54176 14473 54179
rect 13780 54148 14473 54176
rect 13780 54136 13786 54148
rect 14461 54145 14473 54148
rect 14507 54145 14519 54179
rect 14461 54139 14519 54145
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54145 15163 54179
rect 15105 54139 15163 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54145 17095 54179
rect 17037 54139 17095 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54145 17923 54179
rect 17865 54139 17923 54145
rect 18966 54136 18972 54188
rect 19024 54176 19030 54188
rect 19720 54185 19748 54216
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 19024 54148 19441 54176
rect 19024 54136 19030 54148
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 19705 54179 19763 54185
rect 19705 54145 19717 54179
rect 19751 54145 19763 54179
rect 19705 54139 19763 54145
rect 20622 54136 20628 54188
rect 20680 54176 20686 54188
rect 20717 54179 20775 54185
rect 20717 54176 20729 54179
rect 20680 54148 20729 54176
rect 20680 54136 20686 54148
rect 20717 54145 20729 54148
rect 20763 54145 20775 54179
rect 20717 54139 20775 54145
rect 21726 54136 21732 54188
rect 21784 54176 21790 54188
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21784 54148 22017 54176
rect 21784 54136 21790 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 23106 54136 23112 54188
rect 23164 54176 23170 54188
rect 23201 54179 23259 54185
rect 23201 54176 23213 54179
rect 23164 54148 23213 54176
rect 23164 54136 23170 54148
rect 23201 54145 23213 54148
rect 23247 54145 23259 54179
rect 23201 54139 23259 54145
rect 24486 54136 24492 54188
rect 24544 54176 24550 54188
rect 24581 54179 24639 54185
rect 24581 54176 24593 54179
rect 24544 54148 24593 54176
rect 24544 54136 24550 54148
rect 24581 54145 24593 54148
rect 24627 54145 24639 54179
rect 24581 54139 24639 54145
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 5166 54068 5172 54120
rect 5224 54068 5230 54120
rect 7834 54068 7840 54120
rect 7892 54068 7898 54120
rect 9306 54068 9312 54120
rect 9364 54108 9370 54120
rect 9861 54111 9919 54117
rect 9861 54108 9873 54111
rect 9364 54080 9873 54108
rect 9364 54068 9370 54080
rect 9861 54077 9873 54080
rect 9907 54077 9919 54111
rect 9861 54071 9919 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 12621 54071 12679 54077
rect 15838 54000 15844 54052
rect 15896 54040 15902 54052
rect 22189 54043 22247 54049
rect 22189 54040 22201 54043
rect 15896 54012 22201 54040
rect 15896 54000 15902 54012
rect 22189 54009 22201 54012
rect 22235 54009 22247 54043
rect 22189 54003 22247 54009
rect 12434 53932 12440 53984
rect 12492 53972 12498 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 12492 53944 14289 53972
rect 12492 53932 12498 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 14277 53935 14335 53941
rect 14918 53932 14924 53984
rect 14976 53932 14982 53984
rect 16114 53932 16120 53984
rect 16172 53972 16178 53984
rect 16853 53975 16911 53981
rect 16853 53972 16865 53975
rect 16172 53944 16865 53972
rect 16172 53932 16178 53944
rect 16853 53941 16865 53944
rect 16899 53941 16911 53975
rect 16853 53935 16911 53941
rect 17678 53932 17684 53984
rect 17736 53932 17742 53984
rect 20898 53932 20904 53984
rect 20956 53932 20962 53984
rect 24670 53932 24676 53984
rect 24728 53972 24734 53984
rect 24765 53975 24823 53981
rect 24765 53972 24777 53975
rect 24728 53944 24777 53972
rect 24728 53932 24734 53944
rect 24765 53941 24777 53944
rect 24811 53941 24823 53975
rect 24765 53935 24823 53941
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 10686 53660 10692 53712
rect 10744 53660 10750 53712
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 3786 53592 3792 53644
rect 3844 53632 3850 53644
rect 4433 53635 4491 53641
rect 4433 53632 4445 53635
rect 3844 53604 4445 53632
rect 3844 53592 3850 53604
rect 4433 53601 4445 53604
rect 4479 53601 4491 53635
rect 4433 53595 4491 53601
rect 6546 53592 6552 53644
rect 6604 53632 6610 53644
rect 7101 53635 7159 53641
rect 7101 53632 7113 53635
rect 6604 53604 7113 53632
rect 6604 53592 6610 53604
rect 7101 53601 7113 53604
rect 7147 53601 7159 53635
rect 10704 53632 10732 53660
rect 11241 53635 11299 53641
rect 11241 53632 11253 53635
rect 10704 53604 11253 53632
rect 7101 53595 7159 53601
rect 11241 53601 11253 53604
rect 11287 53601 11299 53635
rect 11241 53595 11299 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 4157 53567 4215 53573
rect 4157 53533 4169 53567
rect 4203 53564 4215 53567
rect 6638 53564 6644 53576
rect 4203 53536 6644 53564
rect 4203 53533 4215 53536
rect 4157 53527 4215 53533
rect 1780 53496 1808 53527
rect 6638 53524 6644 53536
rect 6696 53524 6702 53576
rect 6825 53567 6883 53573
rect 6825 53533 6837 53567
rect 6871 53564 6883 53567
rect 7834 53564 7840 53576
rect 6871 53536 7840 53564
rect 6871 53533 6883 53536
rect 6825 53527 6883 53533
rect 7834 53524 7840 53536
rect 7892 53524 7898 53576
rect 10686 53524 10692 53576
rect 10744 53564 10750 53576
rect 10781 53567 10839 53573
rect 10781 53564 10793 53567
rect 10744 53536 10793 53564
rect 10744 53524 10750 53536
rect 10781 53533 10793 53536
rect 10827 53533 10839 53567
rect 10781 53527 10839 53533
rect 23109 53567 23167 53573
rect 23109 53533 23121 53567
rect 23155 53564 23167 53567
rect 23290 53564 23296 53576
rect 23155 53536 23296 53564
rect 23155 53533 23167 53536
rect 23109 53527 23167 53533
rect 23290 53524 23296 53536
rect 23348 53524 23354 53576
rect 23750 53524 23756 53576
rect 23808 53524 23814 53576
rect 25038 53524 25044 53576
rect 25096 53524 25102 53576
rect 5534 53496 5540 53508
rect 1780 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 22094 53388 22100 53440
rect 22152 53428 22158 53440
rect 23201 53431 23259 53437
rect 23201 53428 23213 53431
rect 22152 53400 23213 53428
rect 22152 53388 22158 53400
rect 23201 53397 23213 53400
rect 23247 53397 23259 53431
rect 23201 53391 23259 53397
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 25225 53431 25283 53437
rect 25225 53397 25237 53431
rect 25271 53428 25283 53431
rect 26510 53428 26516 53440
rect 25271 53400 26516 53428
rect 25271 53397 25283 53400
rect 25225 53391 25283 53397
rect 26510 53388 26516 53400
rect 26568 53388 26574 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 4062 53184 4068 53236
rect 4120 53224 4126 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 4120 53196 5181 53224
rect 4120 53184 4126 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 5353 53091 5411 53097
rect 5353 53057 5365 53091
rect 5399 53088 5411 53091
rect 7742 53088 7748 53100
rect 5399 53060 7748 53088
rect 5399 53057 5411 53060
rect 5353 53051 5411 53057
rect 7742 53048 7748 53060
rect 7800 53048 7806 53100
rect 23382 53048 23388 53100
rect 23440 53088 23446 53100
rect 24305 53091 24363 53097
rect 24305 53088 24317 53091
rect 23440 53060 24317 53088
rect 23440 53048 23446 53060
rect 24305 53057 24317 53060
rect 24351 53057 24363 53091
rect 24305 53051 24363 53057
rect 25038 53048 25044 53100
rect 25096 53048 25102 53100
rect 19978 52844 19984 52896
rect 20036 52884 20042 52896
rect 24489 52887 24547 52893
rect 24489 52884 24501 52887
rect 20036 52856 24501 52884
rect 20036 52844 20042 52856
rect 24489 52853 24501 52856
rect 24535 52853 24547 52887
rect 24489 52847 24547 52853
rect 25225 52887 25283 52893
rect 25225 52853 25237 52887
rect 25271 52884 25283 52887
rect 25774 52884 25780 52896
rect 25271 52856 25780 52884
rect 25271 52853 25283 52856
rect 25225 52847 25283 52853
rect 25774 52844 25780 52856
rect 25832 52844 25838 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 25317 52479 25375 52485
rect 25317 52445 25329 52479
rect 25363 52476 25375 52479
rect 25958 52476 25964 52488
rect 25363 52448 25964 52476
rect 25363 52445 25375 52448
rect 25317 52439 25375 52445
rect 25958 52436 25964 52448
rect 26016 52436 26022 52488
rect 24946 52368 24952 52420
rect 25004 52368 25010 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 6638 52096 6644 52148
rect 6696 52096 6702 52148
rect 6825 52003 6883 52009
rect 6825 51969 6837 52003
rect 6871 52000 6883 52003
rect 9398 52000 9404 52012
rect 6871 51972 9404 52000
rect 6871 51969 6883 51972
rect 6825 51963 6883 51969
rect 9398 51960 9404 51972
rect 9456 51960 9462 52012
rect 25317 52003 25375 52009
rect 25317 51969 25329 52003
rect 25363 52000 25375 52003
rect 25866 52000 25872 52012
rect 25363 51972 25872 52000
rect 25363 51969 25375 51972
rect 25317 51963 25375 51969
rect 25866 51960 25872 51972
rect 25924 51960 25930 52012
rect 24118 51756 24124 51808
rect 24176 51796 24182 51808
rect 25133 51799 25191 51805
rect 25133 51796 25145 51799
rect 24176 51768 25145 51796
rect 24176 51756 24182 51768
rect 25133 51765 25145 51768
rect 25179 51765 25191 51799
rect 25133 51759 25191 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 7374 51552 7380 51604
rect 7432 51592 7438 51604
rect 8297 51595 8355 51601
rect 8297 51592 8309 51595
rect 7432 51564 8309 51592
rect 7432 51552 7438 51564
rect 8297 51561 8309 51564
rect 8343 51561 8355 51595
rect 8297 51555 8355 51561
rect 7834 51484 7840 51536
rect 7892 51524 7898 51536
rect 9217 51527 9275 51533
rect 9217 51524 9229 51527
rect 7892 51496 9229 51524
rect 7892 51484 7898 51496
rect 9217 51493 9229 51496
rect 9263 51493 9275 51527
rect 9217 51487 9275 51493
rect 4798 51348 4804 51400
rect 4856 51388 4862 51400
rect 7837 51391 7895 51397
rect 7837 51388 7849 51391
rect 4856 51360 7849 51388
rect 4856 51348 4862 51360
rect 7837 51357 7849 51360
rect 7883 51357 7895 51391
rect 7837 51351 7895 51357
rect 8478 51348 8484 51400
rect 8536 51348 8542 51400
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10502 51388 10508 51400
rect 9447 51360 10508 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10502 51348 10508 51360
rect 10560 51348 10566 51400
rect 7653 51323 7711 51329
rect 7653 51289 7665 51323
rect 7699 51320 7711 51323
rect 10594 51320 10600 51332
rect 7699 51292 10600 51320
rect 7699 51289 7711 51292
rect 7653 51283 7711 51289
rect 10594 51280 10600 51292
rect 10652 51280 10658 51332
rect 24946 51280 24952 51332
rect 25004 51280 25010 51332
rect 25038 51212 25044 51264
rect 25096 51212 25102 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24946 50872 24952 50924
rect 25004 50872 25010 50924
rect 17586 50668 17592 50720
rect 17644 50708 17650 50720
rect 25041 50711 25099 50717
rect 25041 50708 25053 50711
rect 17644 50680 25053 50708
rect 17644 50668 17650 50680
rect 25041 50677 25053 50680
rect 25087 50677 25099 50711
rect 25041 50671 25099 50677
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 7837 50507 7895 50513
rect 7837 50504 7849 50507
rect 5592 50476 7849 50504
rect 5592 50464 5598 50476
rect 7837 50473 7849 50476
rect 7883 50504 7895 50507
rect 8386 50504 8392 50516
rect 7883 50476 8392 50504
rect 7883 50473 7895 50476
rect 7837 50467 7895 50473
rect 8386 50464 8392 50476
rect 8444 50464 8450 50516
rect 9582 50464 9588 50516
rect 9640 50464 9646 50516
rect 7742 50396 7748 50448
rect 7800 50436 7806 50448
rect 8021 50439 8079 50445
rect 8021 50436 8033 50439
rect 7800 50408 8033 50436
rect 7800 50396 7806 50408
rect 8021 50405 8033 50408
rect 8067 50436 8079 50439
rect 8294 50436 8300 50448
rect 8067 50408 8300 50436
rect 8067 50405 8079 50408
rect 8021 50399 8079 50405
rect 8294 50396 8300 50408
rect 8352 50396 8358 50448
rect 7561 50303 7619 50309
rect 7561 50269 7573 50303
rect 7607 50300 7619 50303
rect 8570 50300 8576 50312
rect 7607 50272 8576 50300
rect 7607 50269 7619 50272
rect 7561 50263 7619 50269
rect 8570 50260 8576 50272
rect 8628 50260 8634 50312
rect 9493 50303 9551 50309
rect 9493 50269 9505 50303
rect 9539 50300 9551 50303
rect 9582 50300 9588 50312
rect 9539 50272 9588 50300
rect 9539 50269 9551 50272
rect 9493 50263 9551 50269
rect 9582 50260 9588 50272
rect 9640 50260 9646 50312
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 24489 49827 24547 49833
rect 24489 49793 24501 49827
rect 24535 49824 24547 49827
rect 24854 49824 24860 49836
rect 24535 49796 24860 49824
rect 24535 49793 24547 49796
rect 24489 49787 24547 49793
rect 24854 49784 24860 49796
rect 24912 49784 24918 49836
rect 19794 49716 19800 49768
rect 19852 49756 19858 49768
rect 24765 49759 24823 49765
rect 24765 49756 24777 49759
rect 19852 49728 24777 49756
rect 19852 49716 19858 49728
rect 24765 49725 24777 49728
rect 24811 49725 24823 49759
rect 24765 49719 24823 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 10686 49308 10692 49360
rect 10744 49308 10750 49360
rect 11698 49308 11704 49360
rect 11756 49308 11762 49360
rect 10134 49104 10140 49156
rect 10192 49144 10198 49156
rect 10505 49147 10563 49153
rect 10505 49144 10517 49147
rect 10192 49116 10517 49144
rect 10192 49104 10198 49116
rect 10505 49113 10517 49116
rect 10551 49113 10563 49147
rect 10505 49107 10563 49113
rect 10870 49104 10876 49156
rect 10928 49144 10934 49156
rect 11517 49147 11575 49153
rect 11517 49144 11529 49147
rect 10928 49116 11529 49144
rect 10928 49104 10934 49116
rect 11517 49113 11529 49116
rect 11563 49113 11575 49147
rect 11517 49107 11575 49113
rect 25130 49104 25136 49156
rect 25188 49104 25194 49156
rect 25222 49036 25228 49088
rect 25280 49036 25286 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 8386 48832 8392 48884
rect 8444 48832 8450 48884
rect 9950 48804 9956 48816
rect 8142 48776 9956 48804
rect 9950 48764 9956 48776
rect 10008 48764 10014 48816
rect 6641 48671 6699 48677
rect 6641 48637 6653 48671
rect 6687 48637 6699 48671
rect 6641 48631 6699 48637
rect 6917 48671 6975 48677
rect 6917 48637 6929 48671
rect 6963 48668 6975 48671
rect 9490 48668 9496 48680
rect 6963 48640 9496 48668
rect 6963 48637 6975 48640
rect 6917 48631 6975 48637
rect 6656 48532 6684 48631
rect 9490 48628 9496 48640
rect 9548 48628 9554 48680
rect 9122 48600 9128 48612
rect 8036 48572 9128 48600
rect 8036 48532 8064 48572
rect 9122 48560 9128 48572
rect 9180 48560 9186 48612
rect 6656 48504 8064 48532
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 8294 48084 8300 48136
rect 8352 48124 8358 48136
rect 10356 48127 10414 48133
rect 10356 48124 10368 48127
rect 8352 48096 10368 48124
rect 8352 48084 8358 48096
rect 10356 48093 10368 48096
rect 10402 48093 10414 48127
rect 10356 48087 10414 48093
rect 25130 48016 25136 48068
rect 25188 48016 25194 48068
rect 10459 47991 10517 47997
rect 10459 47957 10471 47991
rect 10505 47988 10517 47991
rect 12342 47988 12348 48000
rect 10505 47960 12348 47988
rect 10505 47957 10517 47960
rect 10459 47951 10517 47957
rect 12342 47948 12348 47960
rect 12400 47948 12406 48000
rect 21450 47948 21456 48000
rect 21508 47988 21514 48000
rect 25225 47991 25283 47997
rect 25225 47988 25237 47991
rect 21508 47960 25237 47988
rect 21508 47948 21514 47960
rect 25225 47957 25237 47960
rect 25271 47957 25283 47991
rect 25225 47951 25283 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9214 47744 9220 47796
rect 9272 47784 9278 47796
rect 9398 47784 9404 47796
rect 9272 47756 9404 47784
rect 9272 47744 9278 47756
rect 9398 47744 9404 47756
rect 9456 47784 9462 47796
rect 9861 47787 9919 47793
rect 9861 47784 9873 47787
rect 9456 47756 9873 47784
rect 9456 47744 9462 47756
rect 9861 47753 9873 47756
rect 9907 47753 9919 47787
rect 9861 47747 9919 47753
rect 8570 47608 8576 47660
rect 8628 47648 8634 47660
rect 9401 47651 9459 47657
rect 9401 47648 9413 47651
rect 8628 47620 9413 47648
rect 8628 47608 8634 47620
rect 9401 47617 9413 47620
rect 9447 47648 9459 47651
rect 10226 47648 10232 47660
rect 9447 47620 10232 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 10226 47608 10232 47620
rect 10284 47608 10290 47660
rect 25314 47608 25320 47660
rect 25372 47608 25378 47660
rect 15930 47540 15936 47592
rect 15988 47580 15994 47592
rect 22094 47580 22100 47592
rect 15988 47552 22100 47580
rect 15988 47540 15994 47552
rect 22094 47540 22100 47552
rect 22152 47540 22158 47592
rect 9490 47404 9496 47456
rect 9548 47404 9554 47456
rect 25133 47447 25191 47453
rect 25133 47413 25145 47447
rect 25179 47444 25191 47447
rect 25406 47444 25412 47456
rect 25179 47416 25412 47444
rect 25179 47413 25191 47416
rect 25133 47407 25191 47413
rect 25406 47404 25412 47416
rect 25464 47404 25470 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 14277 47107 14335 47113
rect 14277 47073 14289 47107
rect 14323 47104 14335 47107
rect 14918 47104 14924 47116
rect 14323 47076 14924 47104
rect 14323 47073 14335 47076
rect 14277 47067 14335 47073
rect 14918 47064 14924 47076
rect 14976 47064 14982 47116
rect 9214 46996 9220 47048
rect 9272 47036 9278 47048
rect 11644 47039 11702 47045
rect 11644 47036 11656 47039
rect 9272 47008 11656 47036
rect 9272 46996 9278 47008
rect 11644 47005 11656 47008
rect 11690 47005 11702 47039
rect 11644 46999 11702 47005
rect 11747 46971 11805 46977
rect 11747 46937 11759 46971
rect 11793 46968 11805 46971
rect 14461 46971 14519 46977
rect 14461 46968 14473 46971
rect 11793 46940 14473 46968
rect 11793 46937 11805 46940
rect 11747 46931 11805 46937
rect 14461 46937 14473 46940
rect 14507 46937 14519 46971
rect 14461 46931 14519 46937
rect 16117 46971 16175 46977
rect 16117 46937 16129 46971
rect 16163 46968 16175 46971
rect 21082 46968 21088 46980
rect 16163 46940 21088 46968
rect 16163 46937 16175 46940
rect 16117 46931 16175 46937
rect 21082 46928 21088 46940
rect 21140 46928 21146 46980
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 9766 46656 9772 46708
rect 9824 46696 9830 46708
rect 10594 46696 10600 46708
rect 9824 46668 10600 46696
rect 9824 46656 9830 46668
rect 10594 46656 10600 46668
rect 10652 46696 10658 46708
rect 10689 46699 10747 46705
rect 10689 46696 10701 46699
rect 10652 46668 10701 46696
rect 10652 46656 10658 46668
rect 10689 46665 10701 46668
rect 10735 46665 10747 46699
rect 10689 46659 10747 46665
rect 12342 46588 12348 46640
rect 12400 46588 12406 46640
rect 16114 46628 16120 46640
rect 14476 46600 16120 46628
rect 8294 46520 8300 46572
rect 8352 46520 8358 46572
rect 10226 46520 10232 46572
rect 10284 46520 10290 46572
rect 14476 46569 14504 46600
rect 16114 46588 16120 46600
rect 16172 46588 16178 46640
rect 14461 46563 14519 46569
rect 14461 46529 14473 46563
rect 14507 46529 14519 46563
rect 14461 46523 14519 46529
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 7834 46452 7840 46504
rect 7892 46492 7898 46504
rect 8113 46495 8171 46501
rect 8113 46492 8125 46495
rect 7892 46464 8125 46492
rect 7892 46452 7898 46464
rect 8113 46461 8125 46464
rect 8159 46461 8171 46495
rect 8113 46455 8171 46461
rect 12161 46495 12219 46501
rect 12161 46461 12173 46495
rect 12207 46492 12219 46495
rect 12434 46492 12440 46504
rect 12207 46464 12440 46492
rect 12207 46461 12219 46464
rect 12161 46455 12219 46461
rect 12434 46452 12440 46464
rect 12492 46452 12498 46504
rect 13722 46452 13728 46504
rect 13780 46452 13786 46504
rect 14642 46452 14648 46504
rect 14700 46452 14706 46504
rect 16301 46495 16359 46501
rect 16301 46461 16313 46495
rect 16347 46492 16359 46495
rect 16390 46492 16396 46504
rect 16347 46464 16396 46492
rect 16347 46461 16359 46464
rect 16301 46455 16359 46461
rect 16390 46452 16396 46464
rect 16448 46452 16454 46504
rect 8478 46384 8484 46436
rect 8536 46384 8542 46436
rect 10410 46316 10416 46368
rect 10468 46316 10474 46368
rect 25133 46359 25191 46365
rect 25133 46325 25145 46359
rect 25179 46356 25191 46359
rect 26050 46356 26056 46368
rect 25179 46328 26056 46356
rect 25179 46325 25191 46328
rect 25133 46319 25191 46325
rect 26050 46316 26056 46328
rect 26108 46316 26114 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 12667 46155 12725 46161
rect 12667 46121 12679 46155
rect 12713 46152 12725 46155
rect 14642 46152 14648 46164
rect 12713 46124 14648 46152
rect 12713 46121 12725 46124
rect 12667 46115 12725 46121
rect 14642 46112 14648 46124
rect 14700 46112 14706 46164
rect 15657 46019 15715 46025
rect 15657 45985 15669 46019
rect 15703 46016 15715 46019
rect 17678 46016 17684 46028
rect 15703 45988 17684 46016
rect 15703 45985 15715 45988
rect 15657 45979 15715 45985
rect 17678 45976 17684 45988
rect 17736 45976 17742 46028
rect 10594 45908 10600 45960
rect 10652 45948 10658 45960
rect 12564 45951 12622 45957
rect 12564 45948 12576 45951
rect 10652 45920 12576 45948
rect 10652 45908 10658 45920
rect 12564 45917 12576 45920
rect 12610 45917 12622 45951
rect 12564 45911 12622 45917
rect 12802 45908 12808 45960
rect 12860 45948 12866 45960
rect 13300 45951 13358 45957
rect 13300 45948 13312 45951
rect 12860 45920 13312 45948
rect 12860 45908 12866 45920
rect 13300 45917 13312 45920
rect 13346 45917 13358 45951
rect 13300 45911 13358 45917
rect 25314 45908 25320 45960
rect 25372 45908 25378 45960
rect 13403 45883 13461 45889
rect 13403 45849 13415 45883
rect 13449 45880 13461 45883
rect 15841 45883 15899 45889
rect 15841 45880 15853 45883
rect 13449 45852 15853 45880
rect 13449 45849 13461 45852
rect 13403 45843 13461 45849
rect 15841 45849 15853 45852
rect 15887 45849 15899 45883
rect 15841 45843 15899 45849
rect 17494 45840 17500 45892
rect 17552 45840 17558 45892
rect 25133 45815 25191 45821
rect 25133 45781 25145 45815
rect 25179 45812 25191 45815
rect 25774 45812 25780 45824
rect 25179 45784 25780 45812
rect 25179 45781 25191 45784
rect 25133 45775 25191 45781
rect 25774 45772 25780 45784
rect 25832 45772 25838 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10502 45500 10508 45552
rect 10560 45540 10566 45552
rect 12802 45540 12808 45552
rect 10560 45512 12808 45540
rect 10560 45500 10566 45512
rect 12802 45500 12808 45512
rect 12860 45500 12866 45552
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 9398 45024 9404 45076
rect 9456 45064 9462 45076
rect 10873 45067 10931 45073
rect 10873 45064 10885 45067
rect 9456 45036 10885 45064
rect 9456 45024 9462 45036
rect 10873 45033 10885 45036
rect 10919 45033 10931 45067
rect 10873 45027 10931 45033
rect 9122 44888 9128 44940
rect 9180 44928 9186 44940
rect 9398 44928 9404 44940
rect 9180 44900 9404 44928
rect 9180 44888 9186 44900
rect 9398 44888 9404 44900
rect 9456 44888 9462 44940
rect 9950 44888 9956 44940
rect 10008 44928 10014 44940
rect 10008 44900 10640 44928
rect 10008 44888 10014 44900
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44792 9459 44795
rect 9674 44792 9680 44804
rect 9447 44764 9680 44792
rect 9447 44761 9459 44764
rect 9401 44755 9459 44761
rect 9674 44752 9680 44764
rect 9732 44752 9738 44804
rect 10612 44792 10640 44900
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 10778 44792 10784 44804
rect 10612 44778 10784 44792
rect 10626 44764 10784 44778
rect 10778 44752 10784 44764
rect 10836 44752 10842 44804
rect 9692 44724 9720 44752
rect 10410 44724 10416 44736
rect 9692 44696 10416 44724
rect 10410 44684 10416 44696
rect 10468 44684 10474 44736
rect 24946 44684 24952 44736
rect 25004 44724 25010 44736
rect 25133 44727 25191 44733
rect 25133 44724 25145 44727
rect 25004 44696 25145 44724
rect 25004 44684 25010 44696
rect 25133 44693 25145 44696
rect 25179 44693 25191 44727
rect 25133 44687 25191 44693
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 9582 44480 9588 44532
rect 9640 44480 9646 44532
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 10226 44344 10232 44396
rect 10284 44384 10290 44396
rect 10597 44387 10655 44393
rect 10597 44384 10609 44387
rect 10284 44356 10609 44384
rect 10284 44344 10290 44356
rect 10597 44353 10609 44356
rect 10643 44353 10655 44387
rect 10597 44347 10655 44353
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25133 44387 25191 44393
rect 25133 44384 25145 44387
rect 24820 44356 25145 44384
rect 24820 44344 24826 44356
rect 25133 44353 25145 44356
rect 25179 44353 25191 44387
rect 25133 44347 25191 44353
rect 8938 44276 8944 44328
rect 8996 44276 9002 44328
rect 10502 44208 10508 44260
rect 10560 44248 10566 44260
rect 10560 44220 11008 44248
rect 10560 44208 10566 44220
rect 10980 44192 11008 44220
rect 17678 44208 17684 44260
rect 17736 44248 17742 44260
rect 25222 44248 25228 44260
rect 17736 44220 25228 44248
rect 17736 44208 17742 44220
rect 25222 44208 25228 44220
rect 25280 44208 25286 44260
rect 25317 44251 25375 44257
rect 25317 44217 25329 44251
rect 25363 44248 25375 44251
rect 25498 44248 25504 44260
rect 25363 44220 25504 44248
rect 25363 44217 25375 44220
rect 25317 44211 25375 44217
rect 25498 44208 25504 44220
rect 25556 44208 25562 44260
rect 10686 44140 10692 44192
rect 10744 44140 10750 44192
rect 10962 44140 10968 44192
rect 11020 44180 11026 44192
rect 11057 44183 11115 44189
rect 11057 44180 11069 44183
rect 11020 44152 11069 44180
rect 11020 44140 11026 44152
rect 11057 44149 11069 44152
rect 11103 44149 11115 44183
rect 11057 44143 11115 44149
rect 17218 44140 17224 44192
rect 17276 44180 17282 44192
rect 23934 44180 23940 44192
rect 17276 44152 23940 44180
rect 17276 44140 17282 44152
rect 23934 44140 23940 44152
rect 23992 44140 23998 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 20717 43843 20775 43849
rect 20717 43809 20729 43843
rect 20763 43840 20775 43843
rect 24118 43840 24124 43852
rect 20763 43812 24124 43840
rect 20763 43809 20775 43812
rect 20717 43803 20775 43809
rect 24118 43800 24124 43812
rect 24176 43800 24182 43852
rect 19518 43732 19524 43784
rect 19576 43772 19582 43784
rect 20441 43775 20499 43781
rect 20441 43772 20453 43775
rect 19576 43744 20453 43772
rect 19576 43732 19582 43744
rect 20441 43741 20453 43744
rect 20487 43741 20499 43775
rect 20441 43735 20499 43741
rect 20806 43664 20812 43716
rect 20864 43704 20870 43716
rect 20864 43676 21206 43704
rect 20864 43664 20870 43676
rect 22186 43596 22192 43648
rect 22244 43596 22250 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25130 43256 25136 43308
rect 25188 43256 25194 43308
rect 25222 43052 25228 43104
rect 25280 43052 25286 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 9766 42712 9772 42764
rect 9824 42712 9830 42764
rect 10134 42712 10140 42764
rect 10192 42752 10198 42764
rect 10229 42755 10287 42761
rect 10229 42752 10241 42755
rect 10192 42724 10241 42752
rect 10192 42712 10198 42724
rect 10229 42721 10241 42724
rect 10275 42721 10287 42755
rect 10229 42715 10287 42721
rect 8846 42644 8852 42696
rect 8904 42684 8910 42696
rect 9585 42687 9643 42693
rect 9585 42684 9597 42687
rect 8904 42656 9597 42684
rect 8904 42644 8910 42656
rect 9585 42653 9597 42656
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 25130 42576 25136 42628
rect 25188 42576 25194 42628
rect 25317 42619 25375 42625
rect 25317 42585 25329 42619
rect 25363 42616 25375 42619
rect 26694 42616 26700 42628
rect 25363 42588 26700 42616
rect 25363 42585 25375 42588
rect 25317 42579 25375 42585
rect 26694 42576 26700 42588
rect 26752 42576 26758 42628
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 9674 42304 9680 42356
rect 9732 42344 9738 42356
rect 11149 42347 11207 42353
rect 11149 42344 11161 42347
rect 9732 42316 11161 42344
rect 9732 42304 9738 42316
rect 11149 42313 11161 42316
rect 11195 42313 11207 42347
rect 11149 42307 11207 42313
rect 10778 42168 10784 42220
rect 10836 42168 10842 42220
rect 9398 42100 9404 42152
rect 9456 42100 9462 42152
rect 9674 42100 9680 42152
rect 9732 42140 9738 42152
rect 10686 42140 10692 42152
rect 9732 42112 10692 42140
rect 9732 42100 9738 42112
rect 10686 42100 10692 42112
rect 10744 42100 10750 42152
rect 16298 42032 16304 42084
rect 16356 42072 16362 42084
rect 19978 42072 19984 42084
rect 16356 42044 19984 42072
rect 16356 42032 16362 42044
rect 19978 42032 19984 42044
rect 20036 42032 20042 42084
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 10781 41803 10839 41809
rect 10781 41769 10793 41803
rect 10827 41800 10839 41803
rect 10870 41800 10876 41812
rect 10827 41772 10876 41800
rect 10827 41769 10839 41772
rect 10781 41763 10839 41769
rect 10870 41760 10876 41772
rect 10928 41760 10934 41812
rect 10321 41667 10379 41673
rect 10321 41633 10333 41667
rect 10367 41664 10379 41667
rect 10962 41664 10968 41676
rect 10367 41636 10968 41664
rect 10367 41633 10379 41636
rect 10321 41627 10379 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 9214 41556 9220 41608
rect 9272 41596 9278 41608
rect 10137 41599 10195 41605
rect 10137 41596 10149 41599
rect 9272 41568 10149 41596
rect 9272 41556 9278 41568
rect 10137 41565 10149 41568
rect 10183 41565 10195 41599
rect 10137 41559 10195 41565
rect 25130 41488 25136 41540
rect 25188 41488 25194 41540
rect 25222 41420 25228 41472
rect 25280 41420 25286 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 26418 40916 26424 40928
rect 25179 40888 26424 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 26418 40876 26424 40888
rect 26476 40876 26482 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 22830 40128 22836 40180
rect 22888 40168 22894 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 22888 40140 25145 40168
rect 22888 40128 22894 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 25314 39992 25320 40044
rect 25372 39992 25378 40044
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 25314 39380 25320 39432
rect 25372 39380 25378 39432
rect 23750 39244 23756 39296
rect 23808 39284 23814 39296
rect 25133 39287 25191 39293
rect 25133 39284 25145 39287
rect 23808 39256 25145 39284
rect 23808 39244 23814 39256
rect 25133 39253 25145 39256
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 24854 38292 24860 38344
rect 24912 38332 24918 38344
rect 25222 38332 25228 38344
rect 24912 38304 25228 38332
rect 24912 38292 24918 38304
rect 25222 38292 25228 38304
rect 25280 38292 25286 38344
rect 25314 38292 25320 38344
rect 25372 38292 25378 38344
rect 24854 38156 24860 38208
rect 24912 38196 24918 38208
rect 25133 38199 25191 38205
rect 25133 38196 25145 38199
rect 24912 38168 25145 38196
rect 24912 38156 24918 38168
rect 25133 38165 25145 38168
rect 25179 38165 25191 38199
rect 25133 38159 25191 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 7834 37952 7840 38004
rect 7892 37992 7898 38004
rect 8665 37995 8723 38001
rect 8665 37992 8677 37995
rect 7892 37964 8677 37992
rect 7892 37952 7898 37964
rect 8665 37961 8677 37964
rect 8711 37961 8723 37995
rect 8665 37955 8723 37961
rect 8849 37859 8907 37865
rect 8849 37825 8861 37859
rect 8895 37856 8907 37859
rect 9490 37856 9496 37868
rect 8895 37828 9496 37856
rect 8895 37825 8907 37828
rect 8849 37819 8907 37825
rect 9490 37816 9496 37828
rect 9548 37816 9554 37868
rect 25130 37816 25136 37868
rect 25188 37816 25194 37868
rect 25317 37723 25375 37729
rect 25317 37689 25329 37723
rect 25363 37720 25375 37723
rect 25590 37720 25596 37732
rect 25363 37692 25596 37720
rect 25363 37689 25375 37692
rect 25317 37683 25375 37689
rect 25590 37680 25596 37692
rect 25648 37680 25654 37732
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 15654 37272 15660 37324
rect 15712 37312 15718 37324
rect 18598 37312 18604 37324
rect 15712 37284 18604 37312
rect 15712 37272 15718 37284
rect 18598 37272 18604 37284
rect 18656 37272 18662 37324
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 25130 36728 25136 36780
rect 25188 36728 25194 36780
rect 25225 36567 25283 36573
rect 25225 36533 25237 36567
rect 25271 36564 25283 36567
rect 25271 36536 26096 36564
rect 25271 36533 25283 36536
rect 25225 36527 25283 36533
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 25222 36320 25228 36372
rect 25280 36360 25286 36372
rect 25280 36332 26004 36360
rect 25280 36320 25286 36332
rect 25976 36304 26004 36332
rect 26068 36304 26096 36536
rect 25958 36252 25964 36304
rect 26016 36252 26022 36304
rect 26050 36252 26056 36304
rect 26108 36252 26114 36304
rect 25314 36116 25320 36168
rect 25372 36116 25378 36168
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 36020 25191 36023
rect 25222 36020 25228 36032
rect 25179 35992 25228 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 25222 35980 25228 35992
rect 25280 35980 25286 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 9674 35776 9680 35828
rect 9732 35816 9738 35828
rect 11149 35819 11207 35825
rect 11149 35816 11161 35819
rect 9732 35788 11161 35816
rect 9732 35776 9738 35788
rect 11149 35785 11161 35788
rect 11195 35785 11207 35819
rect 11149 35779 11207 35785
rect 20254 35776 20260 35828
rect 20312 35816 20318 35828
rect 22005 35819 22063 35825
rect 22005 35816 22017 35819
rect 20312 35788 22017 35816
rect 20312 35776 20318 35788
rect 22005 35785 22017 35788
rect 22051 35785 22063 35819
rect 22005 35779 22063 35785
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 25682 35816 25688 35828
rect 22511 35788 25688 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 25682 35776 25688 35788
rect 25740 35776 25746 35828
rect 21082 35708 21088 35760
rect 21140 35708 21146 35760
rect 21177 35751 21235 35757
rect 21177 35717 21189 35751
rect 21223 35748 21235 35751
rect 26326 35748 26332 35760
rect 21223 35720 26332 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 26326 35708 26332 35720
rect 26384 35708 26390 35760
rect 10778 35640 10784 35692
rect 10836 35640 10842 35692
rect 16390 35640 16396 35692
rect 16448 35680 16454 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 16448 35652 22385 35680
rect 16448 35640 16454 35652
rect 22373 35649 22385 35652
rect 22419 35680 22431 35683
rect 22738 35680 22744 35692
rect 22419 35652 22744 35680
rect 22419 35649 22431 35652
rect 22373 35643 22431 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 9398 35572 9404 35624
rect 9456 35572 9462 35624
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 21174 35572 21180 35624
rect 21232 35612 21238 35624
rect 21269 35615 21327 35621
rect 21269 35612 21281 35615
rect 21232 35584 21281 35612
rect 21232 35572 21238 35584
rect 21269 35581 21281 35584
rect 21315 35581 21327 35615
rect 21269 35575 21327 35581
rect 22646 35572 22652 35624
rect 22704 35572 22710 35624
rect 19886 35436 19892 35488
rect 19944 35476 19950 35488
rect 20717 35479 20775 35485
rect 20717 35476 20729 35479
rect 19944 35448 20729 35476
rect 19944 35436 19950 35448
rect 20717 35445 20729 35448
rect 20763 35445 20775 35479
rect 20717 35439 20775 35445
rect 21082 35436 21088 35488
rect 21140 35476 21146 35488
rect 23382 35476 23388 35488
rect 21140 35448 23388 35476
rect 21140 35436 21146 35448
rect 23382 35436 23388 35448
rect 23440 35436 23446 35488
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 23290 35096 23296 35148
rect 23348 35096 23354 35148
rect 17494 35028 17500 35080
rect 17552 35068 17558 35080
rect 20530 35068 20536 35080
rect 17552 35040 20536 35068
rect 17552 35028 17558 35040
rect 20530 35028 20536 35040
rect 20588 35068 20594 35080
rect 23109 35071 23167 35077
rect 23109 35068 23121 35071
rect 20588 35040 23121 35068
rect 20588 35028 20594 35040
rect 23109 35037 23121 35040
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 24946 35068 24952 35080
rect 23247 35040 24952 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22520 34904 22753 34932
rect 22520 34892 22526 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 25133 34935 25191 34941
rect 25133 34901 25145 34935
rect 25179 34932 25191 34935
rect 25682 34932 25688 34944
rect 25179 34904 25688 34932
rect 25179 34901 25191 34904
rect 25133 34895 25191 34901
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 23474 34688 23480 34740
rect 23532 34728 23538 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 23532 34700 25145 34728
rect 23532 34688 23538 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 8938 34144 8944 34196
rect 8996 34184 9002 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 8996 34156 9137 34184
rect 8996 34144 9002 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 21726 34144 21732 34196
rect 21784 34184 21790 34196
rect 25133 34187 25191 34193
rect 25133 34184 25145 34187
rect 21784 34156 25145 34184
rect 21784 34144 21790 34156
rect 25133 34153 25145 34156
rect 25179 34153 25191 34187
rect 25133 34147 25191 34153
rect 9398 34008 9404 34060
rect 9456 34048 9462 34060
rect 15381 34051 15439 34057
rect 15381 34048 15393 34051
rect 9456 34020 15393 34048
rect 9456 34008 9462 34020
rect 15381 34017 15393 34020
rect 15427 34017 15439 34051
rect 15381 34011 15439 34017
rect 19702 34008 19708 34060
rect 19760 34048 19766 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 19760 34020 21649 34048
rect 19760 34008 19766 34020
rect 21637 34017 21649 34020
rect 21683 34048 21695 34051
rect 22278 34048 22284 34060
rect 21683 34020 22284 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 9030 33940 9036 33992
rect 9088 33980 9094 33992
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 9088 33952 9321 33980
rect 9088 33940 9094 33952
rect 9309 33949 9321 33952
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 20806 33940 20812 33992
rect 20864 33940 20870 33992
rect 25314 33940 25320 33992
rect 25372 33940 25378 33992
rect 14642 33872 14648 33924
rect 14700 33872 14706 33924
rect 19705 33915 19763 33921
rect 19705 33881 19717 33915
rect 19751 33912 19763 33915
rect 19978 33912 19984 33924
rect 19751 33884 19984 33912
rect 19751 33881 19763 33884
rect 19705 33875 19763 33881
rect 19978 33872 19984 33884
rect 20036 33872 20042 33924
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 21959 33884 22094 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 22066 33844 22094 33884
rect 22922 33872 22928 33924
rect 22980 33872 22986 33924
rect 22554 33844 22560 33856
rect 22066 33816 22560 33844
rect 22554 33804 22560 33816
rect 22612 33804 22618 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23256 33816 23397 33844
rect 23256 33804 23262 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 22646 33640 22652 33652
rect 19812 33612 22652 33640
rect 19812 33581 19840 33612
rect 22646 33600 22652 33612
rect 22704 33640 22710 33652
rect 23198 33640 23204 33652
rect 22704 33612 23204 33640
rect 22704 33600 22710 33612
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 19797 33575 19855 33581
rect 19797 33541 19809 33575
rect 19843 33541 19855 33575
rect 19797 33535 19855 33541
rect 20806 33532 20812 33584
rect 20864 33532 20870 33584
rect 22278 33572 22284 33584
rect 22020 33544 22284 33572
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 22922 33532 22928 33584
rect 22980 33532 22986 33584
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 25317 33507 25375 33513
rect 25317 33473 25329 33507
rect 25363 33504 25375 33507
rect 25406 33504 25412 33516
rect 25363 33476 25412 33504
rect 25363 33473 25375 33476
rect 25317 33467 25375 33473
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22370 33436 22376 33448
rect 22327 33408 22376 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 22646 33396 22652 33448
rect 22704 33436 22710 33448
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 22704 33408 23765 33436
rect 22704 33396 22710 33408
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20438 33300 20444 33312
rect 20036 33272 20444 33300
rect 20036 33260 20042 33272
rect 20438 33260 20444 33272
rect 20496 33300 20502 33312
rect 21269 33303 21327 33309
rect 21269 33300 21281 33303
rect 20496 33272 21281 33300
rect 20496 33260 20502 33272
rect 21269 33269 21281 33272
rect 21315 33269 21327 33303
rect 21269 33263 21327 33269
rect 22922 33260 22928 33312
rect 22980 33300 22986 33312
rect 23658 33300 23664 33312
rect 22980 33272 23664 33300
rect 22980 33260 22986 33272
rect 23658 33260 23664 33272
rect 23716 33260 23722 33312
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25866 33300 25872 33312
rect 25179 33272 25872 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25866 33260 25872 33272
rect 25924 33260 25930 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 20898 33096 20904 33108
rect 16724 33068 20904 33096
rect 16724 33056 16730 33068
rect 20898 33056 20904 33068
rect 20956 33056 20962 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 23290 33096 23296 33108
rect 22428 33068 23296 33096
rect 22428 33056 22434 33068
rect 23290 33056 23296 33068
rect 23348 33096 23354 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 23348 33068 24041 33096
rect 23348 33056 23354 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 25222 33056 25228 33108
rect 25280 33096 25286 33108
rect 25682 33096 25688 33108
rect 25280 33068 25688 33096
rect 25280 33056 25286 33068
rect 25682 33056 25688 33068
rect 25740 33056 25746 33108
rect 23566 32988 23572 33040
rect 23624 33028 23630 33040
rect 24581 33031 24639 33037
rect 24581 33028 24593 33031
rect 23624 33000 24593 33028
rect 23624 32988 23630 33000
rect 24581 32997 24593 33000
rect 24627 32997 24639 33031
rect 26418 33028 26424 33040
rect 24581 32991 24639 32997
rect 25056 33000 26424 33028
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 23842 32960 23848 32972
rect 22603 32932 23848 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 23842 32920 23848 32932
rect 23900 32960 23906 32972
rect 24762 32960 24768 32972
rect 23900 32932 24768 32960
rect 23900 32920 23906 32932
rect 24762 32920 24768 32932
rect 24820 32920 24826 32972
rect 25056 32969 25084 33000
rect 26418 32988 26424 33000
rect 26476 32988 26482 33040
rect 25041 32963 25099 32969
rect 25041 32929 25053 32963
rect 25087 32929 25099 32963
rect 25041 32923 25099 32929
rect 25130 32920 25136 32972
rect 25188 32920 25194 32972
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 20717 32895 20775 32901
rect 20717 32892 20729 32895
rect 19484 32864 20729 32892
rect 19484 32852 19490 32864
rect 20717 32861 20729 32864
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 23658 32852 23664 32904
rect 23716 32852 23722 32904
rect 14642 32784 14648 32836
rect 14700 32824 14706 32836
rect 19981 32827 20039 32833
rect 19981 32824 19993 32827
rect 14700 32796 19993 32824
rect 14700 32784 14706 32796
rect 19981 32793 19993 32796
rect 20027 32824 20039 32827
rect 20346 32824 20352 32836
rect 20027 32796 20352 32824
rect 20027 32793 20039 32796
rect 19981 32787 20039 32793
rect 20346 32784 20352 32796
rect 20404 32784 20410 32836
rect 24949 32827 25007 32833
rect 24949 32793 24961 32827
rect 24995 32824 25007 32827
rect 25222 32824 25228 32836
rect 24995 32796 25228 32824
rect 24995 32793 25007 32796
rect 24949 32787 25007 32793
rect 25222 32784 25228 32796
rect 25280 32784 25286 32836
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 21174 32552 21180 32564
rect 19812 32524 21180 32552
rect 14274 32444 14280 32496
rect 14332 32484 14338 32496
rect 14642 32484 14648 32496
rect 14332 32456 14648 32484
rect 14332 32444 14338 32456
rect 14642 32444 14648 32456
rect 14700 32484 14706 32496
rect 15381 32487 15439 32493
rect 15381 32484 15393 32487
rect 14700 32456 15393 32484
rect 14700 32444 14706 32456
rect 15381 32453 15393 32456
rect 15427 32453 15439 32487
rect 15381 32447 15439 32453
rect 18322 32444 18328 32496
rect 18380 32444 18386 32496
rect 19812 32493 19840 32524
rect 21174 32512 21180 32524
rect 21232 32512 21238 32564
rect 24486 32552 24492 32564
rect 24136 32524 24492 32552
rect 19797 32487 19855 32493
rect 19797 32453 19809 32487
rect 19843 32453 19855 32487
rect 19797 32447 19855 32453
rect 20806 32444 20812 32496
rect 20864 32444 20870 32496
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22833 32487 22891 32493
rect 22833 32484 22845 32487
rect 22336 32456 22845 32484
rect 22336 32444 22342 32456
rect 22833 32453 22845 32456
rect 22879 32484 22891 32487
rect 22879 32456 23520 32484
rect 22879 32453 22891 32456
rect 22833 32447 22891 32453
rect 19426 32376 19432 32428
rect 19484 32416 19490 32428
rect 23492 32425 23520 32456
rect 23658 32444 23664 32496
rect 23716 32484 23722 32496
rect 24136 32484 24164 32524
rect 24486 32512 24492 32524
rect 24544 32512 24550 32564
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 25225 32555 25283 32561
rect 25225 32552 25237 32555
rect 24820 32524 25237 32552
rect 24820 32512 24826 32524
rect 25225 32521 25237 32524
rect 25271 32521 25283 32555
rect 25225 32515 25283 32521
rect 23716 32456 24242 32484
rect 23716 32444 23722 32456
rect 19521 32419 19579 32425
rect 19521 32416 19533 32419
rect 19484 32388 19533 32416
rect 19484 32376 19490 32388
rect 19521 32385 19533 32388
rect 19567 32385 19579 32419
rect 19521 32379 19579 32385
rect 22097 32419 22155 32425
rect 22097 32385 22109 32419
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 12802 32308 12808 32360
rect 12860 32348 12866 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 12860 32320 16129 32348
rect 12860 32308 12866 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 16758 32348 16764 32360
rect 16163 32320 16764 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 16758 32308 16764 32320
rect 16816 32348 16822 32360
rect 17313 32351 17371 32357
rect 17313 32348 17325 32351
rect 16816 32320 17325 32348
rect 16816 32308 16822 32320
rect 17313 32317 17325 32320
rect 17359 32317 17371 32351
rect 17313 32311 17371 32317
rect 17589 32351 17647 32357
rect 17589 32317 17601 32351
rect 17635 32348 17647 32351
rect 18230 32348 18236 32360
rect 17635 32320 18236 32348
rect 17635 32317 17647 32320
rect 17589 32311 17647 32317
rect 18230 32308 18236 32320
rect 18288 32308 18294 32360
rect 20346 32308 20352 32360
rect 20404 32348 20410 32360
rect 22112 32348 22140 32379
rect 20404 32320 22140 32348
rect 23753 32351 23811 32357
rect 20404 32308 20410 32320
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 25130 32348 25136 32360
rect 23799 32320 25136 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 25130 32308 25136 32320
rect 25188 32308 25194 32360
rect 19058 32172 19064 32224
rect 19116 32172 19122 32224
rect 20806 32172 20812 32224
rect 20864 32212 20870 32224
rect 21269 32215 21327 32221
rect 21269 32212 21281 32215
rect 20864 32184 21281 32212
rect 20864 32172 20870 32184
rect 21269 32181 21281 32184
rect 21315 32181 21327 32215
rect 21269 32175 21327 32181
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 18230 31968 18236 32020
rect 18288 32008 18294 32020
rect 18509 32011 18567 32017
rect 18509 32008 18521 32011
rect 18288 31980 18521 32008
rect 18288 31968 18294 31980
rect 18509 31977 18521 31980
rect 18555 32008 18567 32011
rect 18598 32008 18604 32020
rect 18555 31980 18604 32008
rect 18555 31977 18567 31980
rect 18509 31971 18567 31977
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 19702 31968 19708 32020
rect 19760 32008 19766 32020
rect 21637 32011 21695 32017
rect 21637 32008 21649 32011
rect 19760 31980 21649 32008
rect 19760 31968 19766 31980
rect 21637 31977 21649 31980
rect 21683 31977 21695 32011
rect 23750 32008 23756 32020
rect 21637 31971 21695 31977
rect 22480 31980 23756 32008
rect 14090 31900 14096 31952
rect 14148 31940 14154 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 14148 31912 15577 31940
rect 14148 31900 14154 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 15565 31903 15623 31909
rect 19058 31900 19064 31952
rect 19116 31940 19122 31952
rect 19116 31912 19564 31940
rect 19116 31900 19122 31912
rect 16114 31832 16120 31884
rect 16172 31832 16178 31884
rect 16758 31832 16764 31884
rect 16816 31832 16822 31884
rect 17037 31875 17095 31881
rect 17037 31841 17049 31875
rect 17083 31872 17095 31875
rect 18414 31872 18420 31884
rect 17083 31844 18420 31872
rect 17083 31841 17095 31844
rect 17037 31835 17095 31841
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 19426 31832 19432 31884
rect 19484 31832 19490 31884
rect 19536 31872 19564 31912
rect 19705 31875 19763 31881
rect 19705 31872 19717 31875
rect 19536 31844 19717 31872
rect 19705 31841 19717 31844
rect 19751 31872 19763 31875
rect 22189 31875 22247 31881
rect 22189 31872 22201 31875
rect 19751 31844 22201 31872
rect 19751 31841 19763 31844
rect 19705 31835 19763 31841
rect 22189 31841 22201 31844
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31804 16083 31807
rect 16666 31804 16672 31816
rect 16071 31776 16672 31804
rect 16071 31773 16083 31776
rect 16025 31767 16083 31773
rect 16666 31764 16672 31776
rect 16724 31764 16730 31816
rect 22097 31807 22155 31813
rect 22097 31773 22109 31807
rect 22143 31804 22155 31807
rect 22480 31804 22508 31980
rect 23750 31968 23756 31980
rect 23808 31968 23814 32020
rect 23017 31943 23075 31949
rect 23017 31909 23029 31943
rect 23063 31940 23075 31943
rect 23382 31940 23388 31952
rect 23063 31912 23388 31940
rect 23063 31909 23075 31912
rect 23017 31903 23075 31909
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 25096 31912 25145 31940
rect 25096 31900 25102 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 22554 31832 22560 31884
rect 22612 31832 22618 31884
rect 22646 31832 22652 31884
rect 22704 31872 22710 31884
rect 23569 31875 23627 31881
rect 23569 31872 23581 31875
rect 22704 31844 23581 31872
rect 22704 31832 22710 31844
rect 23569 31841 23581 31844
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 22143 31776 22508 31804
rect 22572 31804 22600 31832
rect 22830 31804 22836 31816
rect 22572 31776 22836 31804
rect 22143 31773 22155 31776
rect 22097 31767 22155 31773
rect 22830 31764 22836 31776
rect 22888 31764 22894 31816
rect 22922 31764 22928 31816
rect 22980 31804 22986 31816
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 22980 31776 23489 31804
rect 22980 31764 22986 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 25314 31764 25320 31816
rect 25372 31764 25378 31816
rect 18322 31736 18328 31748
rect 18262 31708 18328 31736
rect 18322 31696 18328 31708
rect 18380 31696 18386 31748
rect 21082 31736 21088 31748
rect 20930 31708 21088 31736
rect 21082 31696 21088 31708
rect 21140 31736 21146 31748
rect 21266 31736 21272 31748
rect 21140 31708 21272 31736
rect 21140 31696 21146 31708
rect 21266 31696 21272 31708
rect 21324 31696 21330 31748
rect 22005 31739 22063 31745
rect 22005 31705 22017 31739
rect 22051 31736 22063 31739
rect 22738 31736 22744 31748
rect 22051 31708 22744 31736
rect 22051 31705 22063 31708
rect 22005 31699 22063 31705
rect 22738 31696 22744 31708
rect 22796 31696 22802 31748
rect 15933 31671 15991 31677
rect 15933 31637 15945 31671
rect 15979 31668 15991 31671
rect 17126 31668 17132 31680
rect 15979 31640 17132 31668
rect 15979 31637 15991 31640
rect 15933 31631 15991 31637
rect 17126 31628 17132 31640
rect 17184 31628 17190 31680
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 21177 31671 21235 31677
rect 21177 31668 21189 31671
rect 21048 31640 21189 31668
rect 21048 31628 21054 31640
rect 21177 31637 21189 31640
rect 21223 31637 21235 31671
rect 21177 31631 21235 31637
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 23290 31668 23296 31680
rect 22428 31640 23296 31668
rect 22428 31628 22434 31640
rect 23290 31628 23296 31640
rect 23348 31668 23354 31680
rect 23385 31671 23443 31677
rect 23385 31668 23397 31671
rect 23348 31640 23397 31668
rect 23348 31628 23354 31640
rect 23385 31637 23397 31640
rect 23431 31637 23443 31671
rect 23385 31631 23443 31637
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 20625 31467 20683 31473
rect 13556 31436 16160 31464
rect 13556 31405 13584 31436
rect 16132 31408 16160 31436
rect 20625 31433 20637 31467
rect 20671 31464 20683 31467
rect 24854 31464 24860 31476
rect 20671 31436 24860 31464
rect 20671 31433 20683 31436
rect 20625 31427 20683 31433
rect 24854 31424 24860 31436
rect 24912 31424 24918 31476
rect 13541 31399 13599 31405
rect 13541 31365 13553 31399
rect 13587 31365 13599 31399
rect 14918 31396 14924 31408
rect 14766 31368 14924 31396
rect 13541 31359 13599 31365
rect 14918 31356 14924 31368
rect 14976 31356 14982 31408
rect 16114 31356 16120 31408
rect 16172 31396 16178 31408
rect 16172 31368 17540 31396
rect 16172 31356 16178 31368
rect 15838 31288 15844 31340
rect 15896 31328 15902 31340
rect 15933 31331 15991 31337
rect 15933 31328 15945 31331
rect 15896 31300 15945 31328
rect 15896 31288 15902 31300
rect 15933 31297 15945 31300
rect 15979 31297 15991 31331
rect 15933 31291 15991 31297
rect 16022 31288 16028 31340
rect 16080 31288 16086 31340
rect 17218 31288 17224 31340
rect 17276 31288 17282 31340
rect 17512 31328 17540 31368
rect 20530 31356 20536 31408
rect 20588 31396 20594 31408
rect 22094 31396 22100 31408
rect 20588 31368 22100 31396
rect 20588 31356 20594 31368
rect 22094 31356 22100 31368
rect 22152 31356 22158 31408
rect 22646 31356 22652 31408
rect 22704 31356 22710 31408
rect 24486 31396 24492 31408
rect 23874 31368 24492 31396
rect 24486 31356 24492 31368
rect 24544 31356 24550 31408
rect 22186 31328 22192 31340
rect 17512 31300 22192 31328
rect 12802 31220 12808 31272
rect 12860 31260 12866 31272
rect 13265 31263 13323 31269
rect 13265 31260 13277 31263
rect 12860 31232 13277 31260
rect 12860 31220 12866 31232
rect 13265 31229 13277 31232
rect 13311 31229 13323 31263
rect 13265 31223 13323 31229
rect 16206 31220 16212 31272
rect 16264 31220 16270 31272
rect 17310 31220 17316 31272
rect 17368 31220 17374 31272
rect 17512 31269 17540 31300
rect 22186 31288 22192 31300
rect 22244 31288 22250 31340
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22373 31331 22431 31337
rect 22373 31328 22385 31331
rect 22336 31300 22385 31328
rect 22336 31288 22342 31300
rect 22373 31297 22385 31300
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 17497 31263 17555 31269
rect 17497 31229 17509 31263
rect 17543 31229 17555 31263
rect 17497 31223 17555 31229
rect 18414 31220 18420 31272
rect 18472 31260 18478 31272
rect 18690 31260 18696 31272
rect 18472 31232 18696 31260
rect 18472 31220 18478 31232
rect 18690 31220 18696 31232
rect 18748 31260 18754 31272
rect 20717 31263 20775 31269
rect 20717 31260 20729 31263
rect 18748 31232 20729 31260
rect 18748 31220 18754 31232
rect 20717 31229 20729 31232
rect 20763 31229 20775 31263
rect 24670 31260 24676 31272
rect 20717 31223 20775 31229
rect 22066 31232 24676 31260
rect 14550 31152 14556 31204
rect 14608 31192 14614 31204
rect 16853 31195 16911 31201
rect 16853 31192 16865 31195
rect 14608 31164 16865 31192
rect 14608 31152 14614 31164
rect 16853 31161 16865 31164
rect 16899 31161 16911 31195
rect 16853 31155 16911 31161
rect 17126 31152 17132 31204
rect 17184 31192 17190 31204
rect 22066 31192 22094 31232
rect 24670 31220 24676 31232
rect 24728 31220 24734 31272
rect 17184 31164 22094 31192
rect 17184 31152 17190 31164
rect 15010 31084 15016 31136
rect 15068 31084 15074 31136
rect 15565 31127 15623 31133
rect 15565 31093 15577 31127
rect 15611 31124 15623 31127
rect 15930 31124 15936 31136
rect 15611 31096 15936 31124
rect 15611 31093 15623 31096
rect 15565 31087 15623 31093
rect 15930 31084 15936 31096
rect 15988 31084 15994 31136
rect 18506 31084 18512 31136
rect 18564 31124 18570 31136
rect 20165 31127 20223 31133
rect 20165 31124 20177 31127
rect 18564 31096 20177 31124
rect 18564 31084 18570 31096
rect 20165 31093 20177 31096
rect 20211 31093 20223 31127
rect 20165 31087 20223 31093
rect 23658 31084 23664 31136
rect 23716 31124 23722 31136
rect 24121 31127 24179 31133
rect 24121 31124 24133 31127
rect 23716 31096 24133 31124
rect 23716 31084 23722 31096
rect 24121 31093 24133 31096
rect 24167 31093 24179 31127
rect 24121 31087 24179 31093
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 25133 31127 25191 31133
rect 25133 31124 25145 31127
rect 25004 31096 25145 31124
rect 25004 31084 25010 31096
rect 25133 31093 25145 31096
rect 25179 31093 25191 31127
rect 25133 31087 25191 31093
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 9125 30923 9183 30929
rect 9125 30889 9137 30923
rect 9171 30920 9183 30923
rect 9214 30920 9220 30932
rect 9171 30892 9220 30920
rect 9171 30889 9183 30892
rect 9125 30883 9183 30889
rect 9214 30880 9220 30892
rect 9272 30880 9278 30932
rect 17402 30880 17408 30932
rect 17460 30920 17466 30932
rect 18509 30923 18567 30929
rect 17460 30892 18460 30920
rect 17460 30880 17466 30892
rect 18432 30852 18460 30892
rect 18509 30889 18521 30923
rect 18555 30920 18567 30923
rect 18690 30920 18696 30932
rect 18555 30892 18696 30920
rect 18555 30889 18567 30892
rect 18509 30883 18567 30889
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 22373 30923 22431 30929
rect 20732 30892 22094 30920
rect 20732 30852 20760 30892
rect 18432 30824 20760 30852
rect 22066 30852 22094 30892
rect 22373 30889 22385 30923
rect 22419 30920 22431 30923
rect 22646 30920 22652 30932
rect 22419 30892 22652 30920
rect 22419 30889 22431 30892
rect 22373 30883 22431 30889
rect 22646 30880 22652 30892
rect 22704 30880 22710 30932
rect 26234 30852 26240 30864
rect 22066 30824 26240 30852
rect 26234 30812 26240 30824
rect 26292 30812 26298 30864
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30784 16819 30787
rect 19426 30784 19432 30796
rect 16807 30756 19432 30784
rect 16807 30753 16819 30756
rect 16761 30747 16819 30753
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 20625 30787 20683 30793
rect 20625 30784 20637 30787
rect 19484 30756 20637 30784
rect 19484 30744 19490 30756
rect 20625 30753 20637 30756
rect 20671 30753 20683 30787
rect 20625 30747 20683 30753
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 26510 30784 26516 30796
rect 21048 30756 26516 30784
rect 21048 30744 21054 30756
rect 26510 30744 26516 30756
rect 26568 30744 26574 30796
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9309 30719 9367 30725
rect 9309 30716 9321 30719
rect 8812 30688 9321 30716
rect 8812 30676 8818 30688
rect 9309 30685 9321 30688
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 14274 30676 14280 30728
rect 14332 30676 14338 30728
rect 20162 30676 20168 30728
rect 20220 30676 20226 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25406 30716 25412 30728
rect 25363 30688 25412 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 13906 30608 13912 30660
rect 13964 30648 13970 30660
rect 15013 30651 15071 30657
rect 15013 30648 15025 30651
rect 13964 30620 15025 30648
rect 13964 30608 13970 30620
rect 15013 30617 15025 30620
rect 15059 30617 15071 30651
rect 15013 30611 15071 30617
rect 17037 30651 17095 30657
rect 17037 30617 17049 30651
rect 17083 30617 17095 30651
rect 18322 30648 18328 30660
rect 18262 30620 18328 30648
rect 17037 30611 17095 30617
rect 17052 30580 17080 30611
rect 18322 30608 18328 30620
rect 18380 30648 18386 30660
rect 18690 30648 18696 30660
rect 18380 30620 18696 30648
rect 18380 30608 18386 30620
rect 18690 30608 18696 30620
rect 18748 30608 18754 30660
rect 20898 30608 20904 30660
rect 20956 30608 20962 30660
rect 21284 30620 21390 30648
rect 21284 30592 21312 30620
rect 18782 30580 18788 30592
rect 17052 30552 18788 30580
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 21266 30540 21272 30592
rect 21324 30540 21330 30592
rect 22738 30540 22744 30592
rect 22796 30580 22802 30592
rect 25133 30583 25191 30589
rect 25133 30580 25145 30583
rect 22796 30552 25145 30580
rect 22796 30540 22802 30552
rect 25133 30549 25145 30552
rect 25179 30549 25191 30583
rect 25133 30543 25191 30549
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 12802 30376 12808 30388
rect 12360 30348 12808 30376
rect 12360 30308 12388 30348
rect 12802 30336 12808 30348
rect 12860 30336 12866 30388
rect 16022 30336 16028 30388
rect 16080 30376 16086 30388
rect 20990 30376 20996 30388
rect 16080 30348 20996 30376
rect 16080 30336 16086 30348
rect 20990 30336 20996 30348
rect 21048 30336 21054 30388
rect 11716 30280 12388 30308
rect 7650 30200 7656 30252
rect 7708 30240 7714 30252
rect 11716 30249 11744 30280
rect 14274 30268 14280 30320
rect 14332 30268 14338 30320
rect 20162 30268 20168 30320
rect 20220 30268 20226 30320
rect 20254 30268 20260 30320
rect 20312 30268 20318 30320
rect 22462 30268 22468 30320
rect 22520 30268 22526 30320
rect 24578 30268 24584 30320
rect 24636 30268 24642 30320
rect 9033 30243 9091 30249
rect 9033 30240 9045 30243
rect 7708 30212 9045 30240
rect 7708 30200 7714 30212
rect 9033 30209 9045 30212
rect 9079 30209 9091 30243
rect 9033 30203 9091 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 14918 30240 14924 30252
rect 13110 30226 14924 30240
rect 11701 30203 11759 30209
rect 13096 30212 14924 30226
rect 11977 30175 12035 30181
rect 11977 30141 11989 30175
rect 12023 30172 12035 30175
rect 12710 30172 12716 30184
rect 12023 30144 12716 30172
rect 12023 30141 12035 30144
rect 11977 30135 12035 30141
rect 12710 30132 12716 30144
rect 12768 30132 12774 30184
rect 8846 30064 8852 30116
rect 8904 30064 8910 30116
rect 10778 29996 10784 30048
rect 10836 30036 10842 30048
rect 12526 30036 12532 30048
rect 10836 30008 12532 30036
rect 10836 29996 10842 30008
rect 12526 29996 12532 30008
rect 12584 30036 12590 30048
rect 13096 30036 13124 30212
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 20622 30240 20628 30252
rect 15028 30212 20628 30240
rect 13722 30132 13728 30184
rect 13780 30172 13786 30184
rect 15028 30172 15056 30212
rect 20622 30200 20628 30212
rect 20680 30200 20686 30252
rect 21453 30243 21511 30249
rect 21453 30209 21465 30243
rect 21499 30240 21511 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21499 30212 22385 30240
rect 21499 30209 21511 30212
rect 21453 30203 21511 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 13780 30144 15056 30172
rect 13780 30132 13786 30144
rect 15102 30132 15108 30184
rect 15160 30132 15166 30184
rect 20438 30132 20444 30184
rect 20496 30132 20502 30184
rect 22649 30175 22707 30181
rect 22649 30141 22661 30175
rect 22695 30172 22707 30175
rect 22830 30172 22836 30184
rect 22695 30144 22836 30172
rect 22695 30141 22707 30144
rect 22649 30135 22707 30141
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 23569 30175 23627 30181
rect 23569 30141 23581 30175
rect 23615 30172 23627 30175
rect 23658 30172 23664 30184
rect 23615 30144 23664 30172
rect 23615 30141 23627 30144
rect 23569 30135 23627 30141
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 25041 30175 25099 30181
rect 25041 30141 25053 30175
rect 25087 30172 25099 30175
rect 25130 30172 25136 30184
rect 25087 30144 25136 30172
rect 25087 30141 25099 30144
rect 25041 30135 25099 30141
rect 25130 30132 25136 30144
rect 25188 30132 25194 30184
rect 15562 30064 15568 30116
rect 15620 30104 15626 30116
rect 15620 30076 23428 30104
rect 15620 30064 15626 30076
rect 12584 30008 13124 30036
rect 12584 29996 12590 30008
rect 13446 29996 13452 30048
rect 13504 30036 13510 30048
rect 16114 30036 16120 30048
rect 13504 30008 16120 30036
rect 13504 29996 13510 30008
rect 16114 29996 16120 30008
rect 16172 29996 16178 30048
rect 19242 29996 19248 30048
rect 19300 30036 19306 30048
rect 19797 30039 19855 30045
rect 19797 30036 19809 30039
rect 19300 30008 19809 30036
rect 19300 29996 19306 30008
rect 19797 30005 19809 30008
rect 19843 30005 19855 30039
rect 19797 29999 19855 30005
rect 21910 29996 21916 30048
rect 21968 30036 21974 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21968 30008 22017 30036
rect 21968 29996 21974 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 23400 30036 23428 30076
rect 25958 30036 25964 30048
rect 23400 30008 25964 30036
rect 22005 29999 22063 30005
rect 25958 29996 25964 30008
rect 26016 29996 26022 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 11606 29792 11612 29844
rect 11664 29832 11670 29844
rect 13446 29832 13452 29844
rect 11664 29804 13452 29832
rect 11664 29792 11670 29804
rect 13446 29792 13452 29804
rect 13504 29792 13510 29844
rect 18782 29792 18788 29844
rect 18840 29792 18846 29844
rect 12710 29724 12716 29776
rect 12768 29764 12774 29776
rect 12897 29767 12955 29773
rect 12897 29764 12909 29767
rect 12768 29736 12909 29764
rect 12768 29724 12774 29736
rect 12897 29733 12909 29736
rect 12943 29764 12955 29767
rect 12943 29736 15884 29764
rect 12943 29733 12955 29736
rect 12897 29727 12955 29733
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11422 29696 11428 29708
rect 11195 29668 11428 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 13906 29696 13912 29708
rect 11480 29668 13912 29696
rect 11480 29656 11486 29668
rect 13906 29656 13912 29668
rect 13964 29656 13970 29708
rect 15856 29705 15884 29736
rect 18322 29724 18328 29776
rect 18380 29764 18386 29776
rect 20625 29767 20683 29773
rect 20625 29764 20637 29767
rect 18380 29736 20637 29764
rect 18380 29724 18386 29736
rect 20625 29733 20637 29736
rect 20671 29733 20683 29767
rect 20625 29727 20683 29733
rect 15841 29699 15899 29705
rect 15841 29665 15853 29699
rect 15887 29696 15899 29699
rect 16206 29696 16212 29708
rect 15887 29668 16212 29696
rect 15887 29665 15899 29668
rect 15841 29659 15899 29665
rect 16206 29656 16212 29668
rect 16264 29656 16270 29708
rect 17037 29699 17095 29705
rect 17037 29665 17049 29699
rect 17083 29696 17095 29699
rect 17862 29696 17868 29708
rect 17083 29668 17868 29696
rect 17083 29665 17095 29668
rect 17037 29659 17095 29665
rect 17862 29656 17868 29668
rect 17920 29656 17926 29708
rect 18690 29696 18696 29708
rect 18432 29668 18696 29696
rect 12526 29588 12532 29640
rect 12584 29588 12590 29640
rect 15562 29588 15568 29640
rect 15620 29588 15626 29640
rect 18432 29614 18460 29668
rect 18690 29656 18696 29668
rect 18748 29656 18754 29708
rect 19886 29656 19892 29708
rect 19944 29656 19950 29708
rect 20073 29699 20131 29705
rect 20073 29665 20085 29699
rect 20119 29696 20131 29699
rect 20806 29696 20812 29708
rect 20119 29668 20812 29696
rect 20119 29665 20131 29668
rect 20073 29659 20131 29665
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 21177 29699 21235 29705
rect 21177 29665 21189 29699
rect 21223 29665 21235 29699
rect 21177 29659 21235 29665
rect 18874 29628 18880 29640
rect 18616 29600 18880 29628
rect 11054 29520 11060 29572
rect 11112 29560 11118 29572
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11112 29532 11437 29560
rect 11112 29520 11118 29532
rect 11425 29529 11437 29532
rect 11471 29529 11483 29563
rect 11425 29523 11483 29529
rect 17313 29563 17371 29569
rect 17313 29529 17325 29563
rect 17359 29529 17371 29563
rect 17313 29523 17371 29529
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 15378 29452 15384 29504
rect 15436 29492 15442 29504
rect 15657 29495 15715 29501
rect 15657 29492 15669 29495
rect 15436 29464 15669 29492
rect 15436 29452 15442 29464
rect 15657 29461 15669 29464
rect 15703 29461 15715 29495
rect 17328 29492 17356 29523
rect 18616 29492 18644 29600
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 21192 29628 21220 29659
rect 18932 29600 21220 29628
rect 18932 29588 18938 29600
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 20622 29520 20628 29572
rect 20680 29560 20686 29572
rect 20993 29563 21051 29569
rect 20993 29560 21005 29563
rect 20680 29532 21005 29560
rect 20680 29520 20686 29532
rect 20993 29529 21005 29532
rect 21039 29529 21051 29563
rect 20993 29523 21051 29529
rect 21085 29563 21143 29569
rect 21085 29529 21097 29563
rect 21131 29560 21143 29563
rect 23474 29560 23480 29572
rect 21131 29532 23480 29560
rect 21131 29529 21143 29532
rect 21085 29523 21143 29529
rect 17328 29464 18644 29492
rect 15657 29455 15715 29461
rect 19426 29452 19432 29504
rect 19484 29452 19490 29504
rect 19518 29452 19524 29504
rect 19576 29492 19582 29504
rect 19797 29495 19855 29501
rect 19797 29492 19809 29495
rect 19576 29464 19809 29492
rect 19576 29452 19582 29464
rect 19797 29461 19809 29464
rect 19843 29461 19855 29495
rect 21008 29492 21036 29523
rect 23474 29520 23480 29532
rect 23532 29520 23538 29572
rect 23934 29492 23940 29504
rect 21008 29464 23940 29492
rect 19797 29455 19855 29461
rect 23934 29452 23940 29464
rect 23992 29452 23998 29504
rect 25130 29452 25136 29504
rect 25188 29452 25194 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 9490 29248 9496 29300
rect 9548 29248 9554 29300
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15252 29260 16037 29288
rect 15252 29248 15258 29260
rect 16025 29257 16037 29260
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 16206 29248 16212 29300
rect 16264 29288 16270 29300
rect 19426 29288 19432 29300
rect 16264 29260 19432 29288
rect 16264 29248 16270 29260
rect 19426 29248 19432 29260
rect 19484 29248 19490 29300
rect 19702 29248 19708 29300
rect 19760 29248 19766 29300
rect 24029 29291 24087 29297
rect 24029 29257 24041 29291
rect 24075 29288 24087 29291
rect 24854 29288 24860 29300
rect 24075 29260 24860 29288
rect 24075 29257 24087 29260
rect 24029 29251 24087 29257
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 9861 29223 9919 29229
rect 9861 29189 9873 29223
rect 9907 29220 9919 29223
rect 10318 29220 10324 29232
rect 9907 29192 10324 29220
rect 9907 29189 9919 29192
rect 9861 29183 9919 29189
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 13906 29220 13912 29232
rect 13372 29192 13912 29220
rect 9953 29155 10011 29161
rect 9953 29121 9965 29155
rect 9999 29152 10011 29155
rect 10226 29152 10232 29164
rect 9999 29124 10232 29152
rect 9999 29121 10011 29124
rect 9953 29115 10011 29121
rect 10226 29112 10232 29124
rect 10284 29112 10290 29164
rect 13372 29161 13400 29192
rect 13906 29180 13912 29192
rect 13964 29180 13970 29232
rect 14918 29220 14924 29232
rect 14858 29192 14924 29220
rect 14918 29180 14924 29192
rect 14976 29180 14982 29232
rect 15930 29180 15936 29232
rect 15988 29180 15994 29232
rect 17144 29192 17448 29220
rect 13357 29155 13415 29161
rect 13357 29121 13369 29155
rect 13403 29121 13415 29155
rect 17144 29152 17172 29192
rect 13357 29115 13415 29121
rect 15120 29124 17172 29152
rect 17221 29155 17279 29161
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 9732 29056 10057 29084
rect 9732 29044 9738 29056
rect 10045 29053 10057 29056
rect 10091 29084 10103 29087
rect 10870 29084 10876 29096
rect 10091 29056 10876 29084
rect 10091 29053 10103 29056
rect 10045 29047 10103 29053
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 15120 29093 15148 29124
rect 17221 29121 17233 29155
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 15105 29087 15163 29093
rect 15105 29084 15117 29087
rect 13688 29056 15117 29084
rect 13688 29044 13694 29056
rect 15105 29053 15117 29056
rect 15151 29053 15163 29087
rect 15105 29047 15163 29053
rect 16114 29044 16120 29096
rect 16172 29044 16178 29096
rect 16666 29044 16672 29096
rect 16724 29084 16730 29096
rect 16724 29056 16988 29084
rect 16724 29044 16730 29056
rect 14918 28976 14924 29028
rect 14976 29016 14982 29028
rect 14976 28988 15148 29016
rect 14976 28976 14982 28988
rect 13620 28951 13678 28957
rect 13620 28917 13632 28951
rect 13666 28948 13678 28951
rect 14182 28948 14188 28960
rect 13666 28920 14188 28948
rect 13666 28917 13678 28920
rect 13620 28911 13678 28917
rect 14182 28908 14188 28920
rect 14240 28908 14246 28960
rect 15120 28948 15148 28988
rect 15194 28976 15200 29028
rect 15252 29016 15258 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 15252 28988 15577 29016
rect 15252 28976 15258 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 15804 28988 16865 29016
rect 15804 28976 15810 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16960 29016 16988 29056
rect 17126 29044 17132 29096
rect 17184 29084 17190 29096
rect 17236 29084 17264 29115
rect 17420 29096 17448 29192
rect 23934 29180 23940 29232
rect 23992 29220 23998 29232
rect 25222 29220 25228 29232
rect 23992 29192 25228 29220
rect 23992 29180 23998 29192
rect 25222 29180 25228 29192
rect 25280 29180 25286 29232
rect 18785 29155 18843 29161
rect 18785 29121 18797 29155
rect 18831 29152 18843 29155
rect 19518 29152 19524 29164
rect 18831 29124 19524 29152
rect 18831 29121 18843 29124
rect 18785 29115 18843 29121
rect 19518 29112 19524 29124
rect 19576 29112 19582 29164
rect 19610 29112 19616 29164
rect 19668 29112 19674 29164
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 20404 29124 22201 29152
rect 20404 29112 20410 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 23474 29112 23480 29164
rect 23532 29152 23538 29164
rect 24578 29152 24584 29164
rect 23532 29124 24584 29152
rect 23532 29112 23538 29124
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 24762 29112 24768 29164
rect 24820 29152 24826 29164
rect 24949 29155 25007 29161
rect 24949 29152 24961 29155
rect 24820 29124 24961 29152
rect 24820 29112 24826 29124
rect 24949 29121 24961 29124
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 17184 29056 17264 29084
rect 17313 29087 17371 29093
rect 17184 29044 17190 29056
rect 17313 29053 17325 29087
rect 17359 29053 17371 29087
rect 17313 29047 17371 29053
rect 17328 29016 17356 29047
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 19889 29087 19947 29093
rect 19889 29053 19901 29087
rect 19935 29084 19947 29087
rect 20898 29084 20904 29096
rect 19935 29056 20904 29084
rect 19935 29053 19947 29056
rect 19889 29047 19947 29053
rect 20898 29044 20904 29056
rect 20956 29044 20962 29096
rect 22925 29087 22983 29093
rect 22925 29053 22937 29087
rect 22971 29084 22983 29087
rect 23290 29084 23296 29096
rect 22971 29056 23296 29084
rect 22971 29053 22983 29056
rect 22925 29047 22983 29053
rect 17770 29016 17776 29028
rect 16960 28988 17776 29016
rect 16853 28979 16911 28985
rect 17770 28976 17776 28988
rect 17828 28976 17834 29028
rect 19150 28976 19156 29028
rect 19208 29016 19214 29028
rect 19245 29019 19303 29025
rect 19245 29016 19257 29019
rect 19208 28988 19257 29016
rect 19208 28976 19214 28988
rect 19245 28985 19257 28988
rect 19291 28985 19303 29019
rect 19245 28979 19303 28985
rect 22186 28976 22192 29028
rect 22244 29016 22250 29028
rect 22940 29016 22968 29047
rect 23290 29044 23296 29056
rect 23348 29044 23354 29096
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 24121 29087 24179 29093
rect 24121 29084 24133 29087
rect 23808 29056 24133 29084
rect 23808 29044 23814 29056
rect 24121 29053 24133 29056
rect 24167 29053 24179 29087
rect 24121 29047 24179 29053
rect 22244 28988 22968 29016
rect 23569 29019 23627 29025
rect 22244 28976 22250 28988
rect 23569 28985 23581 29019
rect 23615 29016 23627 29019
rect 24302 29016 24308 29028
rect 23615 28988 24308 29016
rect 23615 28985 23627 28988
rect 23569 28979 23627 28985
rect 24302 28976 24308 28988
rect 24360 28976 24366 29028
rect 24765 29019 24823 29025
rect 24765 28985 24777 29019
rect 24811 29016 24823 29019
rect 24854 29016 24860 29028
rect 24811 28988 24860 29016
rect 24811 28985 24823 28988
rect 24765 28979 24823 28985
rect 24854 28976 24860 28988
rect 24912 28976 24918 29028
rect 18690 28948 18696 28960
rect 15120 28920 18696 28948
rect 18690 28908 18696 28920
rect 18748 28908 18754 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 10870 28704 10876 28756
rect 10928 28704 10934 28756
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 19610 28704 19616 28756
rect 19668 28744 19674 28756
rect 19889 28747 19947 28753
rect 19889 28744 19901 28747
rect 19668 28716 19901 28744
rect 19668 28704 19674 28716
rect 19889 28713 19901 28716
rect 19935 28713 19947 28747
rect 19889 28707 19947 28713
rect 21450 28704 21456 28756
rect 21508 28744 21514 28756
rect 23109 28747 23167 28753
rect 23109 28744 23121 28747
rect 21508 28716 23121 28744
rect 21508 28704 21514 28716
rect 23109 28713 23121 28716
rect 23155 28713 23167 28747
rect 23109 28707 23167 28713
rect 13814 28636 13820 28688
rect 13872 28676 13878 28688
rect 15933 28679 15991 28685
rect 15933 28676 15945 28679
rect 13872 28648 15945 28676
rect 13872 28636 13878 28648
rect 15933 28645 15945 28648
rect 15979 28645 15991 28679
rect 23474 28676 23480 28688
rect 15933 28639 15991 28645
rect 22066 28648 23480 28676
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 10410 28608 10416 28620
rect 9171 28580 10416 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 10410 28568 10416 28580
rect 10468 28608 10474 28620
rect 11422 28608 11428 28620
rect 10468 28580 11428 28608
rect 10468 28568 10474 28580
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 15381 28611 15439 28617
rect 15381 28608 15393 28611
rect 12492 28580 15393 28608
rect 12492 28568 12498 28580
rect 15381 28577 15393 28580
rect 15427 28608 15439 28611
rect 16485 28611 16543 28617
rect 16485 28608 16497 28611
rect 15427 28580 16497 28608
rect 15427 28577 15439 28580
rect 15381 28571 15439 28577
rect 16485 28577 16497 28580
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 19058 28608 19064 28620
rect 17451 28580 19064 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 19058 28568 19064 28580
rect 19116 28568 19122 28620
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 20530 28608 20536 28620
rect 19484 28580 20536 28608
rect 19484 28568 19490 28580
rect 20530 28568 20536 28580
rect 20588 28568 20594 28620
rect 20806 28568 20812 28620
rect 20864 28568 20870 28620
rect 21266 28568 21272 28620
rect 21324 28608 21330 28620
rect 22066 28608 22094 28648
rect 23474 28636 23480 28648
rect 23532 28636 23538 28688
rect 21324 28580 22094 28608
rect 21324 28568 21330 28580
rect 23566 28568 23572 28620
rect 23624 28568 23630 28620
rect 23753 28611 23811 28617
rect 23753 28577 23765 28611
rect 23799 28608 23811 28611
rect 23842 28608 23848 28620
rect 23799 28580 23848 28608
rect 23799 28577 23811 28580
rect 23753 28571 23811 28577
rect 23842 28568 23848 28580
rect 23900 28568 23906 28620
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 15160 28512 17141 28540
rect 15160 28500 15166 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28540 23535 28543
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 23523 28512 24777 28540
rect 23523 28509 23535 28512
rect 23477 28503 23535 28509
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 9401 28475 9459 28481
rect 9401 28441 9413 28475
rect 9447 28472 9459 28475
rect 9674 28472 9680 28484
rect 9447 28444 9680 28472
rect 9447 28441 9459 28444
rect 9401 28435 9459 28441
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 9950 28432 9956 28484
rect 10008 28432 10014 28484
rect 11606 28432 11612 28484
rect 11664 28472 11670 28484
rect 11701 28475 11759 28481
rect 11701 28472 11713 28475
rect 11664 28444 11713 28472
rect 11664 28432 11670 28444
rect 11701 28441 11713 28444
rect 11747 28441 11759 28475
rect 11701 28435 11759 28441
rect 12710 28432 12716 28484
rect 12768 28432 12774 28484
rect 18690 28472 18696 28484
rect 18630 28444 18696 28472
rect 18690 28432 18696 28444
rect 18748 28472 18754 28484
rect 18874 28472 18880 28484
rect 18748 28444 18880 28472
rect 18748 28432 18754 28444
rect 18874 28432 18880 28444
rect 18932 28432 18938 28484
rect 20806 28432 20812 28484
rect 20864 28472 20870 28484
rect 21266 28472 21272 28484
rect 20864 28444 21272 28472
rect 20864 28432 20870 28444
rect 21266 28432 21272 28444
rect 21324 28432 21330 28484
rect 26142 28472 26148 28484
rect 22204 28444 26148 28472
rect 13173 28407 13231 28413
rect 13173 28373 13185 28407
rect 13219 28404 13231 28407
rect 14182 28404 14188 28416
rect 13219 28376 14188 28404
rect 13219 28373 13231 28376
rect 13173 28367 13231 28373
rect 14182 28364 14188 28376
rect 14240 28364 14246 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 14918 28364 14924 28416
rect 14976 28404 14982 28416
rect 15105 28407 15163 28413
rect 15105 28404 15117 28407
rect 14976 28376 15117 28404
rect 14976 28364 14982 28376
rect 15105 28373 15117 28376
rect 15151 28373 15163 28407
rect 15105 28367 15163 28373
rect 15197 28407 15255 28413
rect 15197 28373 15209 28407
rect 15243 28404 15255 28407
rect 15654 28404 15660 28416
rect 15243 28376 15660 28404
rect 15243 28373 15255 28376
rect 15197 28367 15255 28373
rect 15654 28364 15660 28376
rect 15712 28404 15718 28416
rect 15930 28404 15936 28416
rect 15712 28376 15936 28404
rect 15712 28364 15718 28376
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 16298 28364 16304 28416
rect 16356 28364 16362 28416
rect 16390 28364 16396 28416
rect 16448 28404 16454 28416
rect 22204 28404 22232 28444
rect 26142 28432 26148 28444
rect 26200 28432 26206 28484
rect 16448 28376 22232 28404
rect 22281 28407 22339 28413
rect 16448 28364 16454 28376
rect 22281 28373 22293 28407
rect 22327 28404 22339 28407
rect 23750 28404 23756 28416
rect 22327 28376 23756 28404
rect 22327 28373 22339 28376
rect 22281 28367 22339 28373
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 14090 28160 14096 28212
rect 14148 28160 14154 28212
rect 18506 28160 18512 28212
rect 18564 28160 18570 28212
rect 23290 28160 23296 28212
rect 23348 28200 23354 28212
rect 24673 28203 24731 28209
rect 24673 28200 24685 28203
rect 23348 28172 24685 28200
rect 23348 28160 23354 28172
rect 24673 28169 24685 28172
rect 24719 28169 24731 28203
rect 24673 28163 24731 28169
rect 14001 28135 14059 28141
rect 14001 28101 14013 28135
rect 14047 28132 14059 28135
rect 14550 28132 14556 28144
rect 14047 28104 14556 28132
rect 14047 28101 14059 28104
rect 14001 28095 14059 28101
rect 14550 28092 14556 28104
rect 14608 28092 14614 28144
rect 17678 28092 17684 28144
rect 17736 28132 17742 28144
rect 20346 28132 20352 28144
rect 17736 28104 20352 28132
rect 17736 28092 17742 28104
rect 20346 28092 20352 28104
rect 20404 28092 20410 28144
rect 20530 28092 20536 28144
rect 20588 28132 20594 28144
rect 21085 28135 21143 28141
rect 21085 28132 21097 28135
rect 20588 28104 21097 28132
rect 20588 28092 20594 28104
rect 21085 28101 21097 28104
rect 21131 28101 21143 28135
rect 22186 28132 22192 28144
rect 21085 28095 21143 28101
rect 22020 28104 22192 28132
rect 16574 28024 16580 28076
rect 16632 28064 16638 28076
rect 17218 28064 17224 28076
rect 16632 28036 17224 28064
rect 16632 28024 16638 28036
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 22020 28073 22048 28104
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 23658 28092 23664 28144
rect 23716 28132 23722 28144
rect 23716 28104 24808 28132
rect 23716 28092 23722 28104
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 24578 28024 24584 28076
rect 24636 28024 24642 28076
rect 9398 27956 9404 28008
rect 9456 27996 9462 28008
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 9456 27968 14289 27996
rect 9456 27956 9462 27968
rect 14277 27965 14289 27968
rect 14323 27996 14335 27999
rect 15010 27996 15016 28008
rect 14323 27968 15016 27996
rect 14323 27965 14335 27968
rect 14277 27959 14335 27965
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 17310 27956 17316 28008
rect 17368 27956 17374 28008
rect 17402 27956 17408 28008
rect 17460 27956 17466 28008
rect 18598 27956 18604 28008
rect 18656 27956 18662 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 22646 27996 22652 28008
rect 22327 27968 22652 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 22646 27956 22652 27968
rect 22704 27956 22710 28008
rect 24780 28005 24808 28104
rect 24765 27999 24823 28005
rect 24765 27965 24777 27999
rect 24811 27965 24823 27999
rect 24765 27959 24823 27965
rect 12158 27820 12164 27872
rect 12216 27860 12222 27872
rect 13633 27863 13691 27869
rect 13633 27860 13645 27863
rect 12216 27832 13645 27860
rect 12216 27820 12222 27832
rect 13633 27829 13645 27832
rect 13679 27829 13691 27863
rect 13633 27823 13691 27829
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 18049 27863 18107 27869
rect 18049 27829 18061 27863
rect 18095 27860 18107 27863
rect 18782 27860 18788 27872
rect 18095 27832 18788 27860
rect 18095 27829 18107 27832
rect 18049 27823 18107 27829
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 22830 27820 22836 27872
rect 22888 27860 22894 27872
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 22888 27832 23765 27860
rect 22888 27820 22894 27832
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 24210 27820 24216 27872
rect 24268 27820 24274 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 18141 27659 18199 27665
rect 18141 27625 18153 27659
rect 18187 27656 18199 27659
rect 18414 27656 18420 27668
rect 18187 27628 18420 27656
rect 18187 27625 18199 27628
rect 18141 27619 18199 27625
rect 18414 27616 18420 27628
rect 18472 27616 18478 27668
rect 20244 27659 20302 27665
rect 20244 27625 20256 27659
rect 20290 27656 20302 27659
rect 22830 27656 22836 27668
rect 20290 27628 22836 27656
rect 20290 27625 20302 27628
rect 20244 27619 20302 27625
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 23569 27659 23627 27665
rect 23569 27625 23581 27659
rect 23615 27656 23627 27659
rect 24578 27656 24584 27668
rect 23615 27628 24584 27656
rect 23615 27625 23627 27628
rect 23569 27619 23627 27625
rect 24578 27616 24584 27628
rect 24636 27616 24642 27668
rect 22094 27548 22100 27600
rect 22152 27588 22158 27600
rect 22152 27560 23520 27588
rect 22152 27548 22158 27560
rect 9214 27480 9220 27532
rect 9272 27520 9278 27532
rect 10505 27523 10563 27529
rect 10505 27520 10517 27523
rect 9272 27492 10517 27520
rect 9272 27480 9278 27492
rect 10505 27489 10517 27492
rect 10551 27520 10563 27523
rect 13078 27520 13084 27532
rect 10551 27492 13084 27520
rect 10551 27489 10563 27492
rect 10505 27483 10563 27489
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 13538 27480 13544 27532
rect 13596 27480 13602 27532
rect 15010 27480 15016 27532
rect 15068 27520 15074 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15068 27492 15761 27520
rect 15068 27480 15074 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 15749 27483 15807 27489
rect 19981 27523 20039 27529
rect 19981 27489 19993 27523
rect 20027 27520 20039 27523
rect 20027 27492 22094 27520
rect 20027 27489 20039 27492
rect 19981 27483 20039 27489
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 14734 27452 14740 27464
rect 13495 27424 14740 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 22066 27452 22094 27492
rect 22830 27480 22836 27532
rect 22888 27480 22894 27532
rect 22186 27452 22192 27464
rect 22066 27424 22192 27452
rect 22186 27412 22192 27424
rect 22244 27452 22250 27464
rect 23290 27452 23296 27464
rect 22244 27424 23296 27452
rect 22244 27412 22250 27424
rect 23290 27412 23296 27424
rect 23348 27412 23354 27464
rect 23492 27452 23520 27560
rect 25038 27480 25044 27532
rect 25096 27480 25102 27532
rect 25222 27480 25228 27532
rect 25280 27480 25286 27532
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 23492 27424 24961 27452
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 24949 27415 25007 27421
rect 10778 27344 10784 27396
rect 10836 27344 10842 27396
rect 13357 27387 13415 27393
rect 10888 27356 11270 27384
rect 9950 27276 9956 27328
rect 10008 27316 10014 27328
rect 10888 27316 10916 27356
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 13814 27384 13820 27396
rect 13403 27356 13820 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 14274 27344 14280 27396
rect 14332 27384 14338 27396
rect 14918 27384 14924 27396
rect 14332 27356 14924 27384
rect 14332 27344 14338 27356
rect 14918 27344 14924 27356
rect 14976 27384 14982 27396
rect 15565 27387 15623 27393
rect 15565 27384 15577 27387
rect 14976 27356 15577 27384
rect 14976 27344 14982 27356
rect 15565 27353 15577 27356
rect 15611 27384 15623 27387
rect 17494 27384 17500 27396
rect 15611 27356 17500 27384
rect 15611 27353 15623 27356
rect 15565 27347 15623 27353
rect 17494 27344 17500 27356
rect 17552 27344 17558 27396
rect 20806 27344 20812 27396
rect 20864 27344 20870 27396
rect 22649 27387 22707 27393
rect 22649 27353 22661 27387
rect 22695 27384 22707 27387
rect 25866 27384 25872 27396
rect 22695 27356 25872 27384
rect 22695 27353 22707 27356
rect 22649 27347 22707 27353
rect 25866 27344 25872 27356
rect 25924 27344 25930 27396
rect 10008 27288 10916 27316
rect 12253 27319 12311 27325
rect 10008 27276 10014 27288
rect 12253 27285 12265 27319
rect 12299 27316 12311 27319
rect 12434 27316 12440 27328
rect 12299 27288 12440 27316
rect 12299 27285 12311 27288
rect 12253 27279 12311 27285
rect 12434 27276 12440 27288
rect 12492 27276 12498 27328
rect 12526 27276 12532 27328
rect 12584 27316 12590 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12584 27288 13001 27316
rect 12584 27276 12590 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 15197 27319 15255 27325
rect 15197 27285 15209 27319
rect 15243 27316 15255 27319
rect 15286 27316 15292 27328
rect 15243 27288 15292 27316
rect 15243 27285 15255 27288
rect 15197 27279 15255 27285
rect 15286 27276 15292 27288
rect 15344 27276 15350 27328
rect 15657 27319 15715 27325
rect 15657 27285 15669 27319
rect 15703 27316 15715 27319
rect 15930 27316 15936 27328
rect 15703 27288 15936 27316
rect 15703 27285 15715 27288
rect 15657 27279 15715 27285
rect 15930 27276 15936 27288
rect 15988 27276 15994 27328
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19702 27316 19708 27328
rect 19116 27288 19708 27316
rect 19116 27276 19122 27288
rect 19702 27276 19708 27288
rect 19760 27276 19766 27328
rect 20898 27276 20904 27328
rect 20956 27316 20962 27328
rect 21729 27319 21787 27325
rect 21729 27316 21741 27319
rect 20956 27288 21741 27316
rect 20956 27276 20962 27288
rect 21729 27285 21741 27288
rect 21775 27285 21787 27319
rect 21729 27279 21787 27285
rect 21818 27276 21824 27328
rect 21876 27316 21882 27328
rect 22189 27319 22247 27325
rect 22189 27316 22201 27319
rect 21876 27288 22201 27316
rect 21876 27276 21882 27288
rect 22189 27285 22201 27288
rect 22235 27285 22247 27319
rect 22189 27279 22247 27285
rect 22554 27276 22560 27328
rect 22612 27316 22618 27328
rect 22830 27316 22836 27328
rect 22612 27288 22836 27316
rect 22612 27276 22618 27288
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 24581 27319 24639 27325
rect 24581 27316 24593 27319
rect 23532 27288 24593 27316
rect 23532 27276 23538 27288
rect 24581 27285 24593 27288
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27112 11023 27115
rect 11054 27112 11060 27124
rect 11011 27084 11060 27112
rect 11011 27081 11023 27084
rect 10965 27075 11023 27081
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 13078 27072 13084 27124
rect 13136 27112 13142 27124
rect 15102 27112 15108 27124
rect 13136 27084 15108 27112
rect 13136 27072 13142 27084
rect 15102 27072 15108 27084
rect 15160 27072 15166 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16850 27112 16856 27124
rect 15703 27084 16856 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 18874 27072 18880 27124
rect 18932 27112 18938 27124
rect 18932 27084 19564 27112
rect 18932 27072 18938 27084
rect 9950 27004 9956 27056
rect 10008 27004 10014 27056
rect 9214 26936 9220 26988
rect 9272 26936 9278 26988
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 13096 26985 13124 27072
rect 13357 27047 13415 27053
rect 13357 27013 13369 27047
rect 13403 27044 13415 27047
rect 13630 27044 13636 27056
rect 13403 27016 13636 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 13814 27004 13820 27056
rect 13872 27004 13878 27056
rect 15746 27004 15752 27056
rect 15804 27004 15810 27056
rect 19536 27044 19564 27084
rect 19702 27072 19708 27124
rect 19760 27072 19766 27124
rect 21177 27115 21235 27121
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 21726 27112 21732 27124
rect 21223 27084 21732 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 21726 27072 21732 27084
rect 21784 27072 21790 27124
rect 24394 27112 24400 27124
rect 23952 27084 24400 27112
rect 20806 27044 20812 27056
rect 19458 27016 20812 27044
rect 20806 27004 20812 27016
rect 20864 27004 20870 27056
rect 23566 27004 23572 27056
rect 23624 27044 23630 27056
rect 23952 27044 23980 27084
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 23624 27016 24058 27044
rect 23624 27004 23630 27016
rect 13081 26979 13139 26985
rect 13081 26976 13093 26979
rect 12860 26948 13093 26976
rect 12860 26936 12866 26948
rect 13081 26945 13093 26948
rect 13127 26945 13139 26979
rect 13081 26939 13139 26945
rect 15102 26936 15108 26988
rect 15160 26976 15166 26988
rect 16022 26976 16028 26988
rect 15160 26948 16028 26976
rect 15160 26936 15166 26948
rect 16022 26936 16028 26948
rect 16080 26936 16086 26988
rect 17954 26936 17960 26988
rect 18012 26936 18018 26988
rect 21082 26936 21088 26988
rect 21140 26936 21146 26988
rect 9493 26911 9551 26917
rect 9493 26877 9505 26911
rect 9539 26908 9551 26911
rect 10042 26908 10048 26920
rect 9539 26880 10048 26908
rect 9539 26877 9551 26880
rect 9493 26871 9551 26877
rect 10042 26868 10048 26880
rect 10100 26868 10106 26920
rect 15841 26911 15899 26917
rect 15841 26877 15853 26911
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 21269 26911 21327 26917
rect 18279 26880 20852 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 10686 26800 10692 26852
rect 10744 26840 10750 26852
rect 12434 26840 12440 26852
rect 10744 26812 12440 26840
rect 10744 26800 10750 26812
rect 12434 26800 12440 26812
rect 12492 26800 12498 26852
rect 15856 26840 15884 26871
rect 20717 26843 20775 26849
rect 20717 26840 20729 26843
rect 14844 26812 15884 26840
rect 19352 26812 20729 26840
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 14844 26781 14872 26812
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 12032 26744 14841 26772
rect 12032 26732 12038 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 14918 26732 14924 26784
rect 14976 26772 14982 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 14976 26744 15301 26772
rect 14976 26732 14982 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 18598 26732 18604 26784
rect 18656 26772 18662 26784
rect 19352 26772 19380 26812
rect 20717 26809 20729 26812
rect 20763 26809 20775 26843
rect 20824 26840 20852 26880
rect 21269 26877 21281 26911
rect 21315 26877 21327 26911
rect 21269 26871 21327 26877
rect 21284 26840 21312 26871
rect 23290 26868 23296 26920
rect 23348 26868 23354 26920
rect 23569 26911 23627 26917
rect 23569 26877 23581 26911
rect 23615 26908 23627 26911
rect 25222 26908 25228 26920
rect 23615 26880 25228 26908
rect 23615 26877 23627 26880
rect 23569 26871 23627 26877
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 20824 26812 21312 26840
rect 20717 26803 20775 26809
rect 21192 26784 21220 26812
rect 24578 26800 24584 26852
rect 24636 26840 24642 26852
rect 25130 26840 25136 26852
rect 24636 26812 25136 26840
rect 24636 26800 24642 26812
rect 25130 26800 25136 26812
rect 25188 26800 25194 26852
rect 18656 26744 19380 26772
rect 18656 26732 18662 26744
rect 21174 26732 21180 26784
rect 21232 26732 21238 26784
rect 22646 26732 22652 26784
rect 22704 26772 22710 26784
rect 25041 26775 25099 26781
rect 25041 26772 25053 26775
rect 22704 26744 25053 26772
rect 22704 26732 22710 26744
rect 25041 26741 25053 26744
rect 25087 26741 25099 26775
rect 25041 26735 25099 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 12161 26571 12219 26577
rect 12161 26568 12173 26571
rect 10100 26540 12173 26568
rect 10100 26528 10106 26540
rect 12161 26537 12173 26540
rect 12207 26568 12219 26571
rect 13538 26568 13544 26580
rect 12207 26540 13544 26568
rect 12207 26537 12219 26540
rect 12161 26531 12219 26537
rect 13538 26528 13544 26540
rect 13596 26528 13602 26580
rect 21082 26568 21088 26580
rect 14384 26540 21088 26568
rect 11790 26460 11796 26512
rect 11848 26500 11854 26512
rect 14277 26503 14335 26509
rect 14277 26500 14289 26503
rect 11848 26472 14289 26500
rect 11848 26460 11854 26472
rect 14277 26469 14289 26472
rect 14323 26469 14335 26503
rect 14277 26463 14335 26469
rect 10410 26392 10416 26444
rect 10468 26392 10474 26444
rect 10686 26392 10692 26444
rect 10744 26392 10750 26444
rect 12066 26392 12072 26444
rect 12124 26432 12130 26444
rect 14384 26432 14412 26540
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 21174 26528 21180 26580
rect 21232 26528 21238 26580
rect 24581 26571 24639 26577
rect 24581 26537 24593 26571
rect 24627 26568 24639 26571
rect 25038 26568 25044 26580
rect 24627 26540 25044 26568
rect 24627 26537 24639 26540
rect 24581 26531 24639 26537
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 16390 26500 16396 26512
rect 16040 26472 16396 26500
rect 12124 26404 14412 26432
rect 12124 26392 12130 26404
rect 14826 26392 14832 26444
rect 14884 26392 14890 26444
rect 16040 26441 16068 26472
rect 16390 26460 16396 26472
rect 16448 26460 16454 26512
rect 16025 26435 16083 26441
rect 16025 26401 16037 26435
rect 16071 26401 16083 26435
rect 16025 26395 16083 26401
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 15010 26364 15016 26376
rect 14792 26336 15016 26364
rect 14792 26324 14798 26336
rect 15010 26324 15016 26336
rect 15068 26364 15074 26376
rect 16132 26364 16160 26395
rect 17954 26392 17960 26444
rect 18012 26432 18018 26444
rect 19426 26432 19432 26444
rect 18012 26404 19432 26432
rect 18012 26392 18018 26404
rect 19426 26392 19432 26404
rect 19484 26392 19490 26444
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26432 19763 26435
rect 20898 26432 20904 26444
rect 19751 26404 20904 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 20898 26392 20904 26404
rect 20956 26392 20962 26444
rect 15068 26336 16160 26364
rect 15068 26324 15074 26336
rect 18414 26324 18420 26376
rect 18472 26324 18478 26376
rect 20806 26324 20812 26376
rect 20864 26324 20870 26376
rect 21100 26364 21128 26528
rect 21634 26460 21640 26512
rect 21692 26500 21698 26512
rect 22005 26503 22063 26509
rect 22005 26500 22017 26503
rect 21692 26472 22017 26500
rect 21692 26460 21698 26472
rect 22005 26469 22017 26472
rect 22051 26469 22063 26503
rect 22005 26463 22063 26469
rect 22462 26460 22468 26512
rect 22520 26500 22526 26512
rect 22649 26503 22707 26509
rect 22649 26500 22661 26503
rect 22520 26472 22661 26500
rect 22520 26460 22526 26472
rect 22649 26469 22661 26472
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 23845 26503 23903 26509
rect 23845 26469 23857 26503
rect 23891 26500 23903 26503
rect 25406 26500 25412 26512
rect 23891 26472 25412 26500
rect 23891 26469 23903 26472
rect 23845 26463 23903 26469
rect 25406 26460 25412 26472
rect 25464 26460 25470 26512
rect 22278 26392 22284 26444
rect 22336 26432 22342 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 22336 26404 23213 26432
rect 22336 26392 22342 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 23201 26395 23259 26401
rect 23768 26404 24164 26432
rect 21100 26336 22094 26364
rect 9858 26256 9864 26308
rect 9916 26296 9922 26308
rect 14645 26299 14703 26305
rect 9916 26268 11178 26296
rect 9916 26256 9922 26268
rect 11072 26228 11100 26268
rect 14645 26265 14657 26299
rect 14691 26296 14703 26299
rect 15838 26296 15844 26308
rect 14691 26268 15844 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 15838 26256 15844 26268
rect 15896 26296 15902 26308
rect 16850 26296 16856 26308
rect 15896 26268 16856 26296
rect 15896 26256 15902 26268
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 22066 26296 22094 26336
rect 22186 26324 22192 26376
rect 22244 26324 22250 26376
rect 22370 26364 22376 26376
rect 22296 26336 22376 26364
rect 22296 26296 22324 26336
rect 22370 26324 22376 26336
rect 22428 26364 22434 26376
rect 23768 26364 23796 26404
rect 22428 26336 23796 26364
rect 22428 26324 22434 26336
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 24136 26364 24164 26404
rect 24946 26392 24952 26444
rect 25004 26432 25010 26444
rect 25041 26435 25099 26441
rect 25041 26432 25053 26435
rect 25004 26404 25053 26432
rect 25004 26392 25010 26404
rect 25041 26401 25053 26404
rect 25087 26401 25099 26435
rect 25041 26395 25099 26401
rect 25130 26392 25136 26444
rect 25188 26392 25194 26444
rect 24136 26336 24992 26364
rect 22066 26268 22324 26296
rect 22830 26256 22836 26308
rect 22888 26296 22894 26308
rect 23017 26299 23075 26305
rect 23017 26296 23029 26299
rect 22888 26268 23029 26296
rect 22888 26256 22894 26268
rect 23017 26265 23029 26268
rect 23063 26265 23075 26299
rect 23017 26259 23075 26265
rect 23109 26299 23167 26305
rect 23109 26265 23121 26299
rect 23155 26296 23167 26299
rect 24578 26296 24584 26308
rect 23155 26268 24584 26296
rect 23155 26265 23167 26268
rect 23109 26259 23167 26265
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 12710 26228 12716 26240
rect 11072 26200 12716 26228
rect 12710 26188 12716 26200
rect 12768 26228 12774 26240
rect 13814 26228 13820 26240
rect 12768 26200 13820 26228
rect 12768 26188 12774 26200
rect 13814 26188 13820 26200
rect 13872 26188 13878 26240
rect 14737 26231 14795 26237
rect 14737 26197 14749 26231
rect 14783 26228 14795 26231
rect 15102 26228 15108 26240
rect 14783 26200 15108 26228
rect 14783 26197 14795 26200
rect 14737 26191 14795 26197
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 15562 26188 15568 26240
rect 15620 26188 15626 26240
rect 15933 26231 15991 26237
rect 15933 26197 15945 26231
rect 15979 26228 15991 26231
rect 16298 26228 16304 26240
rect 15979 26200 16304 26228
rect 15979 26197 15991 26200
rect 15933 26191 15991 26197
rect 16298 26188 16304 26200
rect 16356 26228 16362 26240
rect 17218 26228 17224 26240
rect 16356 26200 17224 26228
rect 16356 26188 16362 26200
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 24964 26237 24992 26336
rect 25866 26296 25872 26308
rect 25608 26268 25872 26296
rect 24949 26231 25007 26237
rect 24949 26197 24961 26231
rect 24995 26228 25007 26231
rect 25608 26228 25636 26268
rect 25866 26256 25872 26268
rect 25924 26256 25930 26308
rect 24995 26200 25636 26228
rect 24995 26197 25007 26200
rect 24949 26191 25007 26197
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 10778 25984 10784 26036
rect 10836 26024 10842 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10836 25996 10885 26024
rect 10836 25984 10842 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 12069 26027 12127 26033
rect 12069 25993 12081 26027
rect 12115 26024 12127 26027
rect 12115 25996 12434 26024
rect 12115 25993 12127 25996
rect 12069 25987 12127 25993
rect 8938 25916 8944 25968
rect 8996 25956 9002 25968
rect 9398 25956 9404 25968
rect 8996 25928 9404 25956
rect 8996 25916 9002 25928
rect 9398 25916 9404 25928
rect 9456 25916 9462 25968
rect 9858 25916 9864 25968
rect 9916 25916 9922 25968
rect 12406 25956 12434 25996
rect 12526 25984 12532 26036
rect 12584 25984 12590 26036
rect 14001 26027 14059 26033
rect 14001 25993 14013 26027
rect 14047 26024 14059 26027
rect 15194 26024 15200 26036
rect 14047 25996 15200 26024
rect 14047 25993 14059 25996
rect 14001 25987 14059 25993
rect 15194 25984 15200 25996
rect 15252 25984 15258 26036
rect 15289 26027 15347 26033
rect 15289 25993 15301 26027
rect 15335 26024 15347 26027
rect 16758 26024 16764 26036
rect 15335 25996 16764 26024
rect 15335 25993 15347 25996
rect 15289 25987 15347 25993
rect 16758 25984 16764 25996
rect 16816 26024 16822 26036
rect 17586 26024 17592 26036
rect 16816 25996 17592 26024
rect 16816 25984 16822 25996
rect 17586 25984 17592 25996
rect 17644 25984 17650 26036
rect 18233 26027 18291 26033
rect 18233 25993 18245 26027
rect 18279 26024 18291 26027
rect 18414 26024 18420 26036
rect 18279 25996 18420 26024
rect 18279 25993 18291 25996
rect 18233 25987 18291 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 22370 26024 22376 26036
rect 22152 25996 22376 26024
rect 22152 25984 22158 25996
rect 22370 25984 22376 25996
rect 22428 25984 22434 26036
rect 22465 26027 22523 26033
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 22738 26024 22744 26036
rect 22511 25996 22744 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 25222 25984 25228 26036
rect 25280 26024 25286 26036
rect 25317 26027 25375 26033
rect 25317 26024 25329 26027
rect 25280 25996 25329 26024
rect 25280 25984 25286 25996
rect 25317 25993 25329 25996
rect 25363 25993 25375 26027
rect 25317 25987 25375 25993
rect 12406 25928 17080 25956
rect 9122 25848 9128 25900
rect 9180 25848 9186 25900
rect 12434 25848 12440 25900
rect 12492 25848 12498 25900
rect 13280 25860 13584 25888
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 11112 25792 12633 25820
rect 11112 25780 11118 25792
rect 12621 25789 12633 25792
rect 12667 25789 12679 25823
rect 12621 25783 12679 25789
rect 10962 25712 10968 25764
rect 11020 25752 11026 25764
rect 13280 25752 13308 25860
rect 11020 25724 13308 25752
rect 13556 25752 13584 25860
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 17052 25897 17080 25928
rect 18322 25916 18328 25968
rect 18380 25916 18386 25968
rect 24394 25916 24400 25968
rect 24452 25916 24458 25968
rect 13909 25891 13967 25897
rect 13909 25888 13921 25891
rect 13872 25860 13921 25888
rect 13872 25848 13878 25860
rect 13909 25857 13921 25860
rect 13955 25857 13967 25891
rect 15197 25891 15255 25897
rect 13909 25851 13967 25857
rect 14016 25860 14320 25888
rect 13630 25780 13636 25832
rect 13688 25820 13694 25832
rect 14016 25820 14044 25860
rect 13688 25792 14044 25820
rect 13688 25780 13694 25792
rect 14182 25780 14188 25832
rect 14240 25780 14246 25832
rect 14292 25820 14320 25860
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 16209 25891 16267 25897
rect 16209 25888 16221 25891
rect 15243 25860 16221 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 16209 25857 16221 25860
rect 16255 25857 16267 25891
rect 16209 25851 16267 25857
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 14292 25792 15393 25820
rect 15381 25789 15393 25792
rect 15427 25789 15439 25823
rect 15381 25783 15439 25789
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25820 18567 25823
rect 18690 25820 18696 25832
rect 18555 25792 18696 25820
rect 18555 25789 18567 25792
rect 18509 25783 18567 25789
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 22830 25820 22836 25832
rect 22695 25792 22836 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 22830 25780 22836 25792
rect 22888 25780 22894 25832
rect 23290 25780 23296 25832
rect 23348 25820 23354 25832
rect 23566 25820 23572 25832
rect 23348 25792 23572 25820
rect 23348 25780 23354 25792
rect 23566 25780 23572 25792
rect 23624 25780 23630 25832
rect 23845 25823 23903 25829
rect 23845 25789 23857 25823
rect 23891 25820 23903 25823
rect 25222 25820 25228 25832
rect 23891 25792 25228 25820
rect 23891 25789 23903 25792
rect 23845 25783 23903 25789
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 14829 25755 14887 25761
rect 14829 25752 14841 25755
rect 13556 25724 14841 25752
rect 11020 25712 11026 25724
rect 14829 25721 14841 25724
rect 14875 25721 14887 25755
rect 14829 25715 14887 25721
rect 16853 25755 16911 25761
rect 16853 25721 16865 25755
rect 16899 25752 16911 25755
rect 20898 25752 20904 25764
rect 16899 25724 20904 25752
rect 16899 25721 16911 25724
rect 16853 25715 16911 25721
rect 20898 25712 20904 25724
rect 20956 25712 20962 25764
rect 10410 25644 10416 25696
rect 10468 25684 10474 25696
rect 13446 25684 13452 25696
rect 10468 25656 13452 25684
rect 10468 25644 10474 25656
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 13541 25687 13599 25693
rect 13541 25653 13553 25687
rect 13587 25684 13599 25687
rect 16758 25684 16764 25696
rect 13587 25656 16764 25684
rect 13587 25653 13599 25656
rect 13541 25647 13599 25653
rect 16758 25644 16764 25656
rect 16816 25644 16822 25696
rect 16942 25644 16948 25696
rect 17000 25684 17006 25696
rect 17865 25687 17923 25693
rect 17865 25684 17877 25687
rect 17000 25656 17877 25684
rect 17000 25644 17006 25656
rect 17865 25653 17877 25656
rect 17911 25653 17923 25687
rect 17865 25647 17923 25653
rect 19886 25644 19892 25696
rect 19944 25644 19950 25696
rect 20714 25644 20720 25696
rect 20772 25684 20778 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 20772 25656 22017 25684
rect 20772 25644 20778 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 10318 25440 10324 25492
rect 10376 25480 10382 25492
rect 10597 25483 10655 25489
rect 10597 25480 10609 25483
rect 10376 25452 10609 25480
rect 10376 25440 10382 25452
rect 10597 25449 10609 25452
rect 10643 25449 10655 25483
rect 10597 25443 10655 25449
rect 11146 25440 11152 25492
rect 11204 25480 11210 25492
rect 14826 25480 14832 25492
rect 11204 25452 14832 25480
rect 11204 25440 11210 25452
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 13354 25372 13360 25424
rect 13412 25412 13418 25424
rect 13725 25415 13783 25421
rect 13725 25412 13737 25415
rect 13412 25384 13737 25412
rect 13412 25372 13418 25384
rect 13725 25381 13737 25384
rect 13771 25381 13783 25415
rect 16945 25415 17003 25421
rect 13725 25375 13783 25381
rect 13832 25384 16344 25412
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 11149 25347 11207 25353
rect 11149 25344 11161 25347
rect 9732 25316 11161 25344
rect 9732 25304 9738 25316
rect 11149 25313 11161 25316
rect 11195 25313 11207 25347
rect 11149 25307 11207 25313
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12802 25344 12808 25356
rect 12023 25316 12808 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 13832 25344 13860 25384
rect 13504 25316 13860 25344
rect 13504 25304 13510 25316
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 16316 25353 16344 25384
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 16991 25384 21036 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 16301 25347 16359 25353
rect 16301 25313 16313 25347
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 16816 25316 17816 25344
rect 16816 25304 16822 25316
rect 10962 25236 10968 25288
rect 11020 25236 11026 25288
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 17788 25285 17816 25316
rect 17129 25279 17187 25285
rect 17129 25276 17141 25279
rect 13780 25248 17141 25276
rect 13780 25236 13786 25248
rect 17129 25245 17141 25248
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 18874 25236 18880 25288
rect 18932 25236 18938 25288
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21008 25276 21036 25384
rect 21085 25347 21143 25353
rect 21085 25313 21097 25347
rect 21131 25344 21143 25347
rect 23934 25344 23940 25356
rect 21131 25316 23940 25344
rect 21131 25313 21143 25316
rect 21085 25307 21143 25313
rect 23934 25304 23940 25316
rect 23992 25304 23998 25356
rect 21729 25279 21787 25285
rect 21729 25276 21741 25279
rect 21008 25248 21741 25276
rect 21729 25245 21741 25248
rect 21775 25245 21787 25279
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 21729 25239 21787 25245
rect 22066 25248 22661 25276
rect 10778 25168 10784 25220
rect 10836 25208 10842 25220
rect 11057 25211 11115 25217
rect 11057 25208 11069 25211
rect 10836 25180 11069 25208
rect 10836 25168 10842 25180
rect 11057 25177 11069 25180
rect 11103 25177 11115 25211
rect 11057 25171 11115 25177
rect 11974 25168 11980 25220
rect 12032 25208 12038 25220
rect 12253 25211 12311 25217
rect 12253 25208 12265 25211
rect 12032 25180 12265 25208
rect 12032 25168 12038 25180
rect 12253 25177 12265 25180
rect 12299 25177 12311 25211
rect 12253 25171 12311 25177
rect 12710 25168 12716 25220
rect 12768 25168 12774 25220
rect 14645 25211 14703 25217
rect 13556 25180 14320 25208
rect 11698 25100 11704 25152
rect 11756 25140 11762 25152
rect 13556 25140 13584 25180
rect 14292 25149 14320 25180
rect 14645 25177 14657 25211
rect 14691 25208 14703 25211
rect 14826 25208 14832 25220
rect 14691 25180 14832 25208
rect 14691 25177 14703 25180
rect 14645 25171 14703 25177
rect 14826 25168 14832 25180
rect 14884 25208 14890 25220
rect 15470 25208 15476 25220
rect 14884 25180 15476 25208
rect 14884 25168 14890 25180
rect 15470 25168 15476 25180
rect 15528 25168 15534 25220
rect 16117 25211 16175 25217
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16574 25208 16580 25220
rect 16163 25180 16580 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 18506 25208 18512 25220
rect 16868 25180 18512 25208
rect 11756 25112 13584 25140
rect 14277 25143 14335 25149
rect 11756 25100 11762 25112
rect 14277 25109 14289 25143
rect 14323 25109 14335 25143
rect 14277 25103 14335 25109
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 15194 25140 15200 25152
rect 14783 25112 15200 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 15194 25100 15200 25112
rect 15252 25140 15258 25152
rect 15378 25140 15384 25152
rect 15252 25112 15384 25140
rect 15252 25100 15258 25112
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 15930 25100 15936 25152
rect 15988 25140 15994 25152
rect 16209 25143 16267 25149
rect 16209 25140 16221 25143
rect 15988 25112 16221 25140
rect 15988 25100 15994 25112
rect 16209 25109 16221 25112
rect 16255 25140 16267 25143
rect 16868 25140 16896 25180
rect 18506 25168 18512 25180
rect 18564 25168 18570 25220
rect 19978 25168 19984 25220
rect 20036 25168 20042 25220
rect 22066 25208 22094 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 21560 25180 22094 25208
rect 23845 25211 23903 25217
rect 16255 25112 16896 25140
rect 17589 25143 17647 25149
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 17589 25109 17601 25143
rect 17635 25140 17647 25143
rect 19794 25140 19800 25152
rect 17635 25112 19800 25140
rect 17635 25109 17647 25112
rect 17589 25103 17647 25109
rect 19794 25100 19800 25112
rect 19852 25100 19858 25152
rect 21560 25149 21588 25180
rect 23845 25177 23857 25211
rect 23891 25208 23903 25211
rect 24946 25208 24952 25220
rect 23891 25180 24952 25208
rect 23891 25177 23903 25180
rect 23845 25171 23903 25177
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 21545 25143 21603 25149
rect 21545 25109 21557 25143
rect 21591 25109 21603 25143
rect 21545 25103 21603 25109
rect 21726 25100 21732 25152
rect 21784 25140 21790 25152
rect 25133 25143 25191 25149
rect 25133 25140 25145 25143
rect 21784 25112 25145 25140
rect 21784 25100 21790 25112
rect 25133 25109 25145 25112
rect 25179 25109 25191 25143
rect 25133 25103 25191 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 7466 24896 7472 24948
rect 7524 24936 7530 24948
rect 12069 24939 12127 24945
rect 12069 24936 12081 24939
rect 7524 24908 12081 24936
rect 7524 24896 7530 24908
rect 12069 24905 12081 24908
rect 12115 24905 12127 24939
rect 12069 24899 12127 24905
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 18690 24936 18696 24948
rect 17276 24908 18696 24936
rect 17276 24896 17282 24908
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 9858 24828 9864 24880
rect 9916 24868 9922 24880
rect 9916 24840 10074 24868
rect 9916 24828 9922 24840
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 12768 24840 13754 24868
rect 12768 24828 12774 24840
rect 15194 24828 15200 24880
rect 15252 24868 15258 24880
rect 15252 24840 16528 24868
rect 15252 24828 15258 24840
rect 12158 24760 12164 24812
rect 12216 24760 12222 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12860 24772 13001 24800
rect 12860 24760 12866 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 16500 24800 16528 24840
rect 16574 24828 16580 24880
rect 16632 24868 16638 24880
rect 18417 24871 18475 24877
rect 18417 24868 18429 24871
rect 16632 24840 18429 24868
rect 16632 24828 16638 24840
rect 18417 24837 18429 24840
rect 18463 24868 18475 24871
rect 20254 24868 20260 24880
rect 18463 24840 20260 24868
rect 18463 24837 18475 24840
rect 18417 24831 18475 24837
rect 20254 24828 20260 24840
rect 20312 24828 20318 24880
rect 22465 24871 22523 24877
rect 22465 24837 22477 24871
rect 22511 24868 22523 24871
rect 24118 24868 24124 24880
rect 22511 24840 24124 24868
rect 22511 24837 22523 24840
rect 22465 24831 22523 24837
rect 24118 24828 24124 24840
rect 24176 24828 24182 24880
rect 24394 24828 24400 24880
rect 24452 24828 24458 24880
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 16500 24772 17325 24800
rect 12989 24763 13047 24769
rect 17313 24769 17325 24772
rect 17359 24800 17371 24803
rect 17359 24772 18460 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 18432 24744 18460 24772
rect 18506 24760 18512 24812
rect 18564 24800 18570 24812
rect 18564 24772 18736 24800
rect 18564 24760 18570 24772
rect 9306 24692 9312 24744
rect 9364 24692 9370 24744
rect 9585 24735 9643 24741
rect 9585 24701 9597 24735
rect 9631 24732 9643 24735
rect 9674 24732 9680 24744
rect 9631 24704 9680 24732
rect 9631 24701 9643 24704
rect 9585 24695 9643 24701
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 12253 24735 12311 24741
rect 12253 24701 12265 24735
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13354 24732 13360 24744
rect 13311 24704 13360 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 10870 24624 10876 24676
rect 10928 24664 10934 24676
rect 12268 24664 12296 24695
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 14826 24692 14832 24744
rect 14884 24732 14890 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 14884 24704 17417 24732
rect 14884 24692 14890 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 18414 24692 18420 24744
rect 18472 24692 18478 24744
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18708 24732 18736 24772
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 21082 24760 21088 24812
rect 21140 24760 21146 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 23474 24800 23480 24812
rect 22603 24772 23480 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 19610 24732 19616 24744
rect 18708 24704 19616 24732
rect 18601 24695 18659 24701
rect 10928 24636 12296 24664
rect 10928 24624 10934 24636
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 18616 24664 18644 24695
rect 19610 24692 19616 24704
rect 19668 24692 19674 24744
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20438 24732 20444 24744
rect 20027 24704 20444 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22278 24732 22284 24744
rect 21499 24704 22284 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 22278 24692 22284 24704
rect 22336 24692 22342 24744
rect 22646 24692 22652 24744
rect 22704 24692 22710 24744
rect 23290 24692 23296 24744
rect 23348 24732 23354 24744
rect 23566 24732 23572 24744
rect 23348 24704 23572 24732
rect 23348 24692 23354 24704
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25130 24732 25136 24744
rect 23891 24704 25136 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 25222 24692 25228 24744
rect 25280 24732 25286 24744
rect 25317 24735 25375 24741
rect 25317 24732 25329 24735
rect 25280 24704 25329 24732
rect 25280 24692 25286 24704
rect 25317 24701 25329 24704
rect 25363 24701 25375 24735
rect 25317 24695 25375 24701
rect 17092 24636 18644 24664
rect 17092 24624 17098 24636
rect 11057 24599 11115 24605
rect 11057 24565 11069 24599
rect 11103 24596 11115 24599
rect 11146 24596 11152 24608
rect 11103 24568 11152 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 13722 24596 13728 24608
rect 11747 24568 13728 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14734 24556 14740 24608
rect 14792 24556 14798 24608
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15528 24568 16865 24596
rect 15528 24556 15534 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16853 24559 16911 24565
rect 17218 24556 17224 24608
rect 17276 24596 17282 24608
rect 17770 24596 17776 24608
rect 17276 24568 17776 24596
rect 17276 24556 17282 24568
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 19702 24556 19708 24608
rect 19760 24596 19766 24608
rect 20622 24596 20628 24608
rect 19760 24568 20628 24596
rect 19760 24556 19766 24568
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 22097 24599 22155 24605
rect 22097 24565 22109 24599
rect 22143 24596 22155 24599
rect 22186 24596 22192 24608
rect 22143 24568 22192 24596
rect 22143 24565 22155 24568
rect 22097 24559 22155 24565
rect 22186 24556 22192 24568
rect 22244 24556 22250 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 11136 24395 11194 24401
rect 11136 24361 11148 24395
rect 11182 24392 11194 24395
rect 14734 24392 14740 24404
rect 11182 24364 14740 24392
rect 11182 24361 11194 24364
rect 11136 24355 11194 24361
rect 14734 24352 14740 24364
rect 14792 24352 14798 24404
rect 21082 24352 21088 24404
rect 21140 24392 21146 24404
rect 21140 24364 23428 24392
rect 21140 24352 21146 24364
rect 23290 24284 23296 24336
rect 23348 24284 23354 24336
rect 9306 24216 9312 24268
rect 9364 24256 9370 24268
rect 10873 24259 10931 24265
rect 10873 24256 10885 24259
rect 9364 24228 10885 24256
rect 9364 24216 9370 24228
rect 10873 24225 10885 24228
rect 10919 24256 10931 24259
rect 12342 24256 12348 24268
rect 10919 24228 12348 24256
rect 10919 24225 10931 24228
rect 10873 24219 10931 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 18598 24216 18604 24268
rect 18656 24216 18662 24268
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19058 24256 19064 24268
rect 18831 24228 19064 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19426 24216 19432 24268
rect 19484 24216 19490 24268
rect 20438 24216 20444 24268
rect 20496 24256 20502 24268
rect 21177 24259 21235 24265
rect 21177 24256 21189 24259
rect 20496 24228 21189 24256
rect 20496 24216 20502 24228
rect 21177 24225 21189 24228
rect 21223 24225 21235 24259
rect 21177 24219 21235 24225
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 23308 24256 23336 24284
rect 21959 24228 23336 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 17678 24148 17684 24200
rect 17736 24148 17742 24200
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 18874 24188 18880 24200
rect 18555 24160 18880 24188
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 21082 24188 21088 24200
rect 20838 24160 21088 24188
rect 21082 24148 21088 24160
rect 21140 24148 21146 24200
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 15933 24123 15991 24129
rect 9916 24092 11638 24120
rect 9916 24080 9922 24092
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 19705 24123 19763 24129
rect 15979 24092 19656 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 9122 24012 9128 24064
rect 9180 24052 9186 24064
rect 12618 24052 12624 24064
rect 9180 24024 12624 24052
rect 9180 24012 9186 24024
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 18141 24055 18199 24061
rect 18141 24021 18153 24055
rect 18187 24052 18199 24055
rect 18322 24052 18328 24064
rect 18187 24024 18328 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18322 24012 18328 24024
rect 18380 24012 18386 24064
rect 19628 24052 19656 24092
rect 19705 24089 19717 24123
rect 19751 24120 19763 24123
rect 19978 24120 19984 24132
rect 19751 24092 19984 24120
rect 19751 24089 19763 24092
rect 19705 24083 19763 24089
rect 19978 24080 19984 24092
rect 20036 24080 20042 24132
rect 22094 24120 22100 24132
rect 21008 24092 22100 24120
rect 21008 24052 21036 24092
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22278 24120 22284 24132
rect 22235 24092 22284 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 23400 24120 23428 24364
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 24765 24395 24823 24401
rect 24765 24392 24777 24395
rect 24176 24364 24777 24392
rect 24176 24352 24182 24364
rect 24765 24361 24777 24364
rect 24811 24361 24823 24395
rect 24765 24355 24823 24361
rect 24946 24148 24952 24200
rect 25004 24188 25010 24200
rect 25406 24188 25412 24200
rect 25004 24160 25412 24188
rect 25004 24148 25010 24160
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 23566 24120 23572 24132
rect 23400 24106 23572 24120
rect 23414 24092 23572 24106
rect 23566 24080 23572 24092
rect 23624 24120 23630 24132
rect 24394 24120 24400 24132
rect 23624 24092 24400 24120
rect 23624 24080 23630 24092
rect 24394 24080 24400 24092
rect 24452 24080 24458 24132
rect 19628 24024 21036 24052
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23532 24024 23673 24052
rect 23532 24012 23538 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 9858 23848 9864 23860
rect 9416 23820 9864 23848
rect 8662 23740 8668 23792
rect 8720 23780 8726 23792
rect 9033 23783 9091 23789
rect 9033 23780 9045 23783
rect 8720 23752 9045 23780
rect 8720 23740 8726 23752
rect 9033 23749 9045 23752
rect 9079 23780 9091 23783
rect 9122 23780 9128 23792
rect 9079 23752 9128 23780
rect 9079 23749 9091 23752
rect 9033 23743 9091 23749
rect 9122 23740 9128 23752
rect 9180 23740 9186 23792
rect 9416 23780 9444 23820
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 13633 23851 13691 23857
rect 13633 23817 13645 23851
rect 13679 23848 13691 23851
rect 13679 23820 14596 23848
rect 13679 23817 13691 23820
rect 13633 23811 13691 23817
rect 9490 23780 9496 23792
rect 9416 23752 9496 23780
rect 9490 23740 9496 23752
rect 9548 23740 9554 23792
rect 12618 23740 12624 23792
rect 12676 23780 12682 23792
rect 14568 23780 14596 23820
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 15160 23820 17233 23848
rect 15160 23808 15166 23820
rect 17221 23817 17233 23820
rect 17267 23848 17279 23851
rect 19705 23851 19763 23857
rect 17267 23820 18000 23848
rect 17267 23817 17279 23820
rect 17221 23811 17279 23817
rect 15562 23780 15568 23792
rect 12676 23752 13768 23780
rect 14568 23752 15568 23780
rect 12676 23740 12682 23752
rect 13740 23712 13768 23752
rect 15562 23740 15568 23752
rect 15620 23740 15626 23792
rect 15930 23740 15936 23792
rect 15988 23780 15994 23792
rect 15988 23752 17448 23780
rect 15988 23740 15994 23752
rect 13740 23684 13860 23712
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 7892 23616 8769 23644
rect 7892 23604 7898 23616
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 8757 23607 8815 23613
rect 13722 23604 13728 23656
rect 13780 23604 13786 23656
rect 13832 23653 13860 23684
rect 13906 23672 13912 23724
rect 13964 23712 13970 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 13964 23684 14841 23712
rect 13964 23672 13970 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 13817 23647 13875 23653
rect 13817 23613 13829 23647
rect 13863 23613 13875 23647
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 13817 23607 13875 23613
rect 13924 23616 15025 23644
rect 13354 23536 13360 23588
rect 13412 23576 13418 23588
rect 13924 23576 13952 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 17420 23653 17448 23752
rect 17972 23712 18000 23820
rect 19705 23817 19717 23851
rect 19751 23848 19763 23851
rect 19886 23848 19892 23860
rect 19751 23820 19892 23848
rect 19751 23817 19763 23820
rect 19705 23811 19763 23817
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 20898 23808 20904 23860
rect 20956 23808 20962 23860
rect 20993 23851 21051 23857
rect 20993 23817 21005 23851
rect 21039 23848 21051 23851
rect 21818 23848 21824 23860
rect 21039 23820 21824 23848
rect 21039 23817 21051 23820
rect 20993 23811 21051 23817
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 24949 23851 25007 23857
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25130 23848 25136 23860
rect 24995 23820 25136 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 19518 23780 19524 23792
rect 18156 23752 19524 23780
rect 18156 23712 18184 23752
rect 19518 23740 19524 23752
rect 19576 23740 19582 23792
rect 19794 23740 19800 23792
rect 19852 23780 19858 23792
rect 19852 23752 22416 23780
rect 19852 23740 19858 23752
rect 17972 23684 18184 23712
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 22002 23712 22008 23724
rect 18233 23675 18291 23681
rect 19260 23684 22008 23712
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 17276 23616 17325 23644
rect 17276 23604 17282 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 13412 23548 13952 23576
rect 14461 23579 14519 23585
rect 13412 23536 13418 23548
rect 14461 23545 14473 23579
rect 14507 23576 14519 23579
rect 18248 23576 18276 23675
rect 14507 23548 18276 23576
rect 14507 23545 14519 23548
rect 14461 23539 14519 23545
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10502 23508 10508 23520
rect 9732 23480 10508 23508
rect 9732 23468 9738 23480
rect 10502 23468 10508 23480
rect 10560 23468 10566 23520
rect 12250 23468 12256 23520
rect 12308 23508 12314 23520
rect 13265 23511 13323 23517
rect 13265 23508 13277 23511
rect 12308 23480 13277 23508
rect 12308 23468 12314 23480
rect 13265 23477 13277 23480
rect 13311 23477 13323 23511
rect 13265 23471 13323 23477
rect 13722 23468 13728 23520
rect 13780 23508 13786 23520
rect 15286 23508 15292 23520
rect 13780 23480 15292 23508
rect 13780 23468 13786 23480
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 15838 23468 15844 23520
rect 15896 23468 15902 23520
rect 16298 23468 16304 23520
rect 16356 23508 16362 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16356 23480 16865 23508
rect 16356 23468 16362 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 16853 23471 16911 23477
rect 18049 23511 18107 23517
rect 18049 23477 18061 23511
rect 18095 23508 18107 23511
rect 19260 23508 19288 23684
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 22388 23721 22416 23752
rect 24486 23740 24492 23792
rect 24544 23740 24550 23792
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 19702 23644 19708 23656
rect 19484 23616 19708 23644
rect 19484 23604 19490 23616
rect 19702 23604 19708 23616
rect 19760 23644 19766 23656
rect 19797 23647 19855 23653
rect 19797 23644 19809 23647
rect 19760 23616 19809 23644
rect 19760 23604 19766 23616
rect 19797 23613 19809 23616
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 19978 23604 19984 23656
rect 20036 23604 20042 23656
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21085 23647 21143 23653
rect 21085 23644 21097 23647
rect 21048 23616 21097 23644
rect 21048 23604 21054 23616
rect 21085 23613 21097 23616
rect 21131 23613 21143 23647
rect 21085 23607 21143 23613
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 23474 23604 23480 23656
rect 23532 23604 23538 23656
rect 19996 23576 20024 23604
rect 22830 23576 22836 23588
rect 19996 23548 22836 23576
rect 22830 23536 22836 23548
rect 22888 23536 22894 23588
rect 18095 23480 19288 23508
rect 19337 23511 19395 23517
rect 18095 23477 18107 23480
rect 18049 23471 18107 23477
rect 19337 23477 19349 23511
rect 19383 23508 19395 23511
rect 19886 23508 19892 23520
rect 19383 23480 19892 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20530 23468 20536 23520
rect 20588 23468 20594 23520
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 22646 23508 22652 23520
rect 22235 23480 22652 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 22646 23468 22652 23480
rect 22704 23468 22710 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 9030 23264 9036 23316
rect 9088 23304 9094 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 9088 23276 9137 23304
rect 9088 23264 9094 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 14734 23264 14740 23316
rect 14792 23264 14798 23316
rect 16390 23264 16396 23316
rect 16448 23304 16454 23316
rect 17310 23304 17316 23316
rect 16448 23276 17316 23304
rect 16448 23264 16454 23276
rect 17310 23264 17316 23276
rect 17368 23264 17374 23316
rect 18230 23264 18236 23316
rect 18288 23304 18294 23316
rect 18414 23304 18420 23316
rect 18288 23276 18420 23304
rect 18288 23264 18294 23276
rect 18414 23264 18420 23276
rect 18472 23304 18478 23316
rect 20806 23304 20812 23316
rect 18472 23276 20812 23304
rect 18472 23264 18478 23276
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 20898 23264 20904 23316
rect 20956 23264 20962 23316
rect 9214 23196 9220 23248
rect 9272 23236 9278 23248
rect 9272 23208 12434 23236
rect 9272 23196 9278 23208
rect 8570 23128 8576 23180
rect 8628 23168 8634 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 8628 23140 9689 23168
rect 8628 23128 8634 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 11054 23128 11060 23180
rect 11112 23168 11118 23180
rect 11793 23171 11851 23177
rect 11793 23168 11805 23171
rect 11112 23140 11805 23168
rect 11112 23128 11118 23140
rect 11793 23137 11805 23140
rect 11839 23137 11851 23171
rect 12406 23168 12434 23208
rect 13354 23196 13360 23248
rect 13412 23236 13418 23248
rect 15102 23236 15108 23248
rect 13412 23208 15108 23236
rect 13412 23196 13418 23208
rect 15102 23196 15108 23208
rect 15160 23196 15166 23248
rect 16025 23239 16083 23245
rect 16025 23205 16037 23239
rect 16071 23236 16083 23239
rect 16574 23236 16580 23248
rect 16071 23208 16580 23236
rect 16071 23205 16083 23208
rect 16025 23199 16083 23205
rect 16574 23196 16580 23208
rect 16632 23236 16638 23248
rect 17586 23236 17592 23248
rect 16632 23208 17592 23236
rect 16632 23196 16638 23208
rect 17586 23196 17592 23208
rect 17644 23236 17650 23248
rect 21358 23236 21364 23248
rect 17644 23208 21364 23236
rect 17644 23196 17650 23208
rect 21358 23196 21364 23208
rect 21416 23196 21422 23248
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12406 23140 13553 23168
rect 11793 23131 11851 23137
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 13541 23131 13599 23137
rect 13648 23140 15301 23168
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 9490 23100 9496 23112
rect 8444 23072 9496 23100
rect 8444 23060 8450 23072
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 12802 23060 12808 23112
rect 12860 23100 12866 23112
rect 13648 23100 13676 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 18230 23128 18236 23180
rect 18288 23128 18294 23180
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 18598 23168 18604 23180
rect 18463 23140 18604 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 20438 23168 20444 23180
rect 20211 23140 20444 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 23382 23128 23388 23180
rect 23440 23168 23446 23180
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 23440 23140 23489 23168
rect 23440 23128 23446 23140
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 24854 23128 24860 23180
rect 24912 23168 24918 23180
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 24912 23140 25053 23168
rect 24912 23128 24918 23140
rect 25041 23137 25053 23140
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25314 23168 25320 23180
rect 25271 23140 25320 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 12860 23072 13676 23100
rect 15105 23103 15163 23109
rect 12860 23060 12866 23072
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15838 23100 15844 23112
rect 15151 23072 15844 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 18187 23072 18552 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 8846 22992 8852 23044
rect 8904 23032 8910 23044
rect 9585 23035 9643 23041
rect 9585 23032 9597 23035
rect 8904 23004 9597 23032
rect 8904 22992 8910 23004
rect 9585 23001 9597 23004
rect 9631 23001 9643 23035
rect 9585 22995 9643 23001
rect 11609 23035 11667 23041
rect 11609 23001 11621 23035
rect 11655 23032 11667 23035
rect 11790 23032 11796 23044
rect 11655 23004 11796 23032
rect 11655 23001 11667 23004
rect 11609 22995 11667 23001
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 17218 23032 17224 23044
rect 15120 23004 17224 23032
rect 9490 22924 9496 22976
rect 9548 22924 9554 22976
rect 10318 22924 10324 22976
rect 10376 22964 10382 22976
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 10376 22936 11253 22964
rect 10376 22924 10382 22936
rect 11241 22933 11253 22936
rect 11287 22933 11299 22967
rect 11241 22927 11299 22933
rect 12526 22924 12532 22976
rect 12584 22964 12590 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12584 22936 13001 22964
rect 12584 22924 12590 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13354 22924 13360 22976
rect 13412 22924 13418 22976
rect 13449 22967 13507 22973
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 15120 22964 15148 23004
rect 17218 22992 17224 23004
rect 17276 22992 17282 23044
rect 18414 23032 18420 23044
rect 17788 23004 18420 23032
rect 13495 22936 15148 22964
rect 15197 22967 15255 22973
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 15197 22933 15209 22967
rect 15243 22964 15255 22967
rect 16574 22964 16580 22976
rect 15243 22936 16580 22964
rect 15243 22933 15255 22936
rect 15197 22927 15255 22933
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 17788 22973 17816 23004
rect 18414 22992 18420 23004
rect 18472 22992 18478 23044
rect 18524 23032 18552 23072
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 20714 23100 20720 23112
rect 20027 23072 20720 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 21818 23060 21824 23112
rect 21876 23060 21882 23112
rect 22646 23060 22652 23112
rect 22704 23060 22710 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25866 23100 25872 23112
rect 24995 23072 25872 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 18690 23032 18696 23044
rect 18524 23004 18696 23032
rect 18690 22992 18696 23004
rect 18748 23032 18754 23044
rect 20990 23032 20996 23044
rect 18748 23004 20996 23032
rect 18748 22992 18754 23004
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 17773 22967 17831 22973
rect 17773 22933 17785 22967
rect 17819 22933 17831 22967
rect 17773 22927 17831 22933
rect 18506 22924 18512 22976
rect 18564 22964 18570 22976
rect 19521 22967 19579 22973
rect 19521 22964 19533 22967
rect 18564 22936 19533 22964
rect 18564 22924 18570 22936
rect 19521 22933 19533 22936
rect 19567 22933 19579 22967
rect 19521 22927 19579 22933
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 22646 22964 22652 22976
rect 21683 22936 22652 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 22646 22924 22652 22936
rect 22704 22924 22710 22976
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 3418 22720 3424 22772
rect 3476 22760 3482 22772
rect 12066 22760 12072 22772
rect 3476 22732 12072 22760
rect 3476 22720 3482 22732
rect 12066 22720 12072 22732
rect 12124 22720 12130 22772
rect 13446 22760 13452 22772
rect 12636 22732 13452 22760
rect 12636 22704 12664 22732
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 16853 22763 16911 22769
rect 16853 22729 16865 22763
rect 16899 22760 16911 22763
rect 21818 22760 21824 22772
rect 16899 22732 21824 22760
rect 16899 22729 16911 22732
rect 16853 22723 16911 22729
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 8444 22664 8786 22692
rect 8444 22652 8450 22664
rect 12618 22652 12624 22704
rect 12676 22652 12682 22704
rect 12710 22652 12716 22704
rect 12768 22692 12774 22704
rect 12768 22664 13110 22692
rect 12768 22652 12774 22664
rect 17218 22652 17224 22704
rect 17276 22692 17282 22704
rect 19886 22692 19892 22704
rect 17276 22664 19892 22692
rect 17276 22652 17282 22664
rect 19886 22652 19892 22664
rect 19944 22652 19950 22704
rect 21177 22695 21235 22701
rect 21177 22661 21189 22695
rect 21223 22692 21235 22695
rect 21726 22692 21732 22704
rect 21223 22664 21732 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 21726 22652 21732 22664
rect 21784 22652 21790 22704
rect 22370 22692 22376 22704
rect 22066 22664 22376 22692
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8021 22627 8079 22633
rect 8021 22624 8033 22627
rect 7892 22596 8033 22624
rect 7892 22584 7898 22596
rect 8021 22593 8033 22596
rect 8067 22593 8079 22627
rect 8021 22587 8079 22593
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 8297 22559 8355 22565
rect 8297 22525 8309 22559
rect 8343 22556 8355 22559
rect 8343 22528 9720 22556
rect 8343 22525 8355 22528
rect 8297 22519 8355 22525
rect 9692 22488 9720 22528
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 10962 22556 10968 22568
rect 9824 22528 10968 22556
rect 9824 22516 9830 22528
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 17052 22556 17080 22587
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 22066 22624 22094 22664
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 23293 22695 23351 22701
rect 23293 22661 23305 22695
rect 23339 22692 23351 22695
rect 24854 22692 24860 22704
rect 23339 22664 24860 22692
rect 23339 22661 23351 22664
rect 23293 22655 23351 22661
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 21140 22596 22094 22624
rect 22281 22627 22339 22633
rect 21140 22584 21146 22596
rect 22281 22593 22293 22627
rect 22327 22624 22339 22627
rect 23750 22624 23756 22636
rect 22327 22596 23756 22624
rect 22327 22593 22339 22596
rect 22281 22587 22339 22593
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 23934 22584 23940 22636
rect 23992 22584 23998 22636
rect 12768 22528 17080 22556
rect 21269 22559 21327 22565
rect 12768 22516 12774 22528
rect 21269 22525 21281 22559
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 10410 22488 10416 22500
rect 9692 22460 10416 22488
rect 10410 22448 10416 22460
rect 10468 22448 10474 22500
rect 20070 22448 20076 22500
rect 20128 22488 20134 22500
rect 21284 22488 21312 22519
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 20128 22460 21312 22488
rect 20128 22448 20134 22460
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 20162 22380 20168 22432
rect 20220 22380 20226 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 21082 22420 21088 22432
rect 20864 22392 21088 22420
rect 20864 22380 20870 22392
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 10502 22176 10508 22228
rect 10560 22216 10566 22228
rect 21085 22219 21143 22225
rect 10560 22188 12434 22216
rect 10560 22176 10566 22188
rect 10594 22108 10600 22160
rect 10652 22148 10658 22160
rect 11606 22148 11612 22160
rect 10652 22120 11192 22148
rect 10652 22108 10658 22120
rect 11164 22089 11192 22120
rect 11440 22120 11612 22148
rect 11440 22094 11468 22120
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 12406 22148 12434 22188
rect 21085 22185 21097 22219
rect 21131 22216 21143 22219
rect 21131 22188 23704 22216
rect 21131 22185 21143 22188
rect 21085 22179 21143 22185
rect 15746 22148 15752 22160
rect 12406 22120 12480 22148
rect 11348 22089 11468 22094
rect 11149 22083 11207 22089
rect 11149 22049 11161 22083
rect 11195 22049 11207 22083
rect 11149 22043 11207 22049
rect 11333 22083 11468 22089
rect 11333 22049 11345 22083
rect 11379 22066 11468 22083
rect 11379 22049 11391 22066
rect 11333 22043 11391 22049
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12452 22089 12480 22120
rect 15304 22120 15752 22148
rect 15304 22089 15332 22120
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 22830 22108 22836 22160
rect 22888 22148 22894 22160
rect 23293 22151 23351 22157
rect 23293 22148 23305 22151
rect 22888 22120 23305 22148
rect 22888 22108 22894 22120
rect 23293 22117 23305 22120
rect 23339 22117 23351 22151
rect 23293 22111 23351 22117
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 12308 22052 12357 22080
rect 12308 22040 12314 22052
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22049 15439 22083
rect 15381 22043 15439 22049
rect 16301 22083 16359 22089
rect 16301 22049 16313 22083
rect 16347 22080 16359 22083
rect 17034 22080 17040 22092
rect 16347 22052 17040 22080
rect 16347 22049 16359 22052
rect 16301 22043 16359 22049
rect 9858 21972 9864 22024
rect 9916 22012 9922 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9916 21984 10057 22012
rect 9916 21972 9922 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 11054 22012 11060 22024
rect 10192 21984 11060 22012
rect 10192 21972 10198 21984
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 13814 22012 13820 22024
rect 11808 21984 13820 22012
rect 11808 21944 11836 21984
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 15396 22012 15424 22043
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 20165 22083 20223 22089
rect 20165 22080 20177 22083
rect 19668 22052 20177 22080
rect 19668 22040 19674 22052
rect 20165 22049 20177 22052
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 20346 22040 20352 22092
rect 20404 22040 20410 22092
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 23198 22080 23204 22092
rect 21591 22052 23204 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 23676 22080 23704 22188
rect 23750 22176 23756 22228
rect 23808 22176 23814 22228
rect 25222 22148 25228 22160
rect 25148 22120 25228 22148
rect 23676 22052 24992 22080
rect 14148 21984 15424 22012
rect 14148 21972 14154 21984
rect 16022 21972 16028 22024
rect 16080 21972 16086 22024
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 22012 20131 22015
rect 20254 22012 20260 22024
rect 20119 21984 20260 22012
rect 20119 21981 20131 21984
rect 20073 21975 20131 21981
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 22922 21972 22928 22024
rect 22980 21972 22986 22024
rect 24964 22021 24992 22052
rect 25038 22040 25044 22092
rect 25096 22040 25102 22092
rect 25148 22089 25176 22120
rect 25222 22108 25228 22120
rect 25280 22108 25286 22160
rect 25133 22083 25191 22089
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 23937 22015 23995 22021
rect 23937 22012 23949 22015
rect 23308 21984 23949 22012
rect 12710 21944 12716 21956
rect 10704 21916 11836 21944
rect 11900 21916 12716 21944
rect 10704 21885 10732 21916
rect 10689 21879 10747 21885
rect 10689 21845 10701 21879
rect 10735 21845 10747 21879
rect 10689 21839 10747 21845
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11900 21885 11928 21916
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 16574 21904 16580 21956
rect 16632 21944 16638 21956
rect 20622 21944 20628 21956
rect 16632 21916 16790 21944
rect 19720 21916 20628 21944
rect 16632 21904 16638 21916
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21845 11943 21879
rect 11885 21839 11943 21845
rect 12250 21836 12256 21888
rect 12308 21836 12314 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 19720 21885 19748 21916
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 21818 21904 21824 21956
rect 21876 21904 21882 21956
rect 23308 21944 23336 21984
rect 23937 21981 23949 21984
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 23216 21916 23336 21944
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 17184 21848 17785 21876
rect 17184 21836 17190 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 17773 21839 17831 21845
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 22002 21836 22008 21888
rect 22060 21876 22066 21888
rect 23216 21876 23244 21916
rect 22060 21848 23244 21876
rect 22060 21836 22066 21848
rect 23382 21836 23388 21888
rect 23440 21876 23446 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23440 21848 24593 21876
rect 23440 21836 23446 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 7374 21632 7380 21684
rect 7432 21672 7438 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 7432 21644 9781 21672
rect 7432 21632 7438 21644
rect 9769 21641 9781 21644
rect 9815 21672 9827 21675
rect 10134 21672 10140 21684
rect 9815 21644 10140 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 10134 21632 10140 21644
rect 10192 21632 10198 21684
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 12250 21672 12256 21684
rect 10413 21635 10471 21641
rect 10520 21644 12256 21672
rect 8386 21564 8392 21616
rect 8444 21604 8450 21616
rect 8444 21576 8786 21604
rect 8444 21564 8450 21576
rect 7834 21496 7840 21548
rect 7892 21536 7898 21548
rect 8021 21539 8079 21545
rect 8021 21536 8033 21539
rect 7892 21508 8033 21536
rect 7892 21496 7898 21508
rect 8021 21505 8033 21508
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 10520 21468 10548 21644
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 18233 21675 18291 21681
rect 12360 21644 14688 21672
rect 10781 21607 10839 21613
rect 10781 21573 10793 21607
rect 10827 21604 10839 21607
rect 11606 21604 11612 21616
rect 10827 21576 11612 21604
rect 10827 21573 10839 21576
rect 10781 21567 10839 21573
rect 11606 21564 11612 21576
rect 11664 21564 11670 21616
rect 11790 21564 11796 21616
rect 11848 21604 11854 21616
rect 12360 21604 12388 21644
rect 11848 21576 12388 21604
rect 11848 21564 11854 21576
rect 13446 21564 13452 21616
rect 13504 21604 13510 21616
rect 13504 21576 13846 21604
rect 13504 21564 13510 21576
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 11112 21508 11897 21536
rect 11112 21496 11118 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 12342 21496 12348 21548
rect 12400 21536 12406 21548
rect 12710 21536 12716 21548
rect 12400 21508 12716 21536
rect 12400 21496 12406 21508
rect 12710 21496 12716 21508
rect 12768 21536 12774 21548
rect 13081 21539 13139 21545
rect 13081 21536 13093 21539
rect 12768 21508 13093 21536
rect 12768 21496 12774 21508
rect 13081 21505 13093 21508
rect 13127 21505 13139 21539
rect 14660 21536 14688 21644
rect 18233 21641 18245 21675
rect 18279 21641 18291 21675
rect 18233 21635 18291 21641
rect 19245 21675 19303 21681
rect 19245 21641 19257 21675
rect 19291 21672 19303 21675
rect 20162 21672 20168 21684
rect 19291 21644 20168 21672
rect 19291 21641 19303 21644
rect 19245 21635 19303 21641
rect 14826 21564 14832 21616
rect 14884 21604 14890 21616
rect 18248 21604 18276 21635
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 21818 21632 21824 21684
rect 21876 21672 21882 21684
rect 22830 21672 22836 21684
rect 21876 21644 22836 21672
rect 21876 21632 21882 21644
rect 22830 21632 22836 21644
rect 22888 21672 22894 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 22888 21644 25053 21672
rect 22888 21632 22894 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 22554 21604 22560 21616
rect 14884 21576 16574 21604
rect 18248 21576 22560 21604
rect 14884 21564 14890 21576
rect 15565 21539 15623 21545
rect 14660 21508 15056 21536
rect 13081 21499 13139 21505
rect 9364 21440 10548 21468
rect 10873 21471 10931 21477
rect 9364 21428 9370 21440
rect 10873 21437 10885 21471
rect 10919 21437 10931 21471
rect 10873 21431 10931 21437
rect 10888 21400 10916 21431
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21468 13415 21471
rect 14090 21468 14096 21480
rect 13403 21440 14096 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 14384 21440 14841 21468
rect 12158 21400 12164 21412
rect 9692 21372 10824 21400
rect 10888 21372 12164 21400
rect 8284 21335 8342 21341
rect 8284 21301 8296 21335
rect 8330 21332 8342 21335
rect 9692 21332 9720 21372
rect 8330 21304 9720 21332
rect 10796 21332 10824 21372
rect 12158 21360 12164 21372
rect 12216 21360 12222 21412
rect 11146 21332 11152 21344
rect 10796 21304 11152 21332
rect 8330 21301 8342 21304
rect 8284 21295 8342 21301
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 13354 21292 13360 21344
rect 13412 21332 13418 21344
rect 14384 21332 14412 21440
rect 14829 21437 14841 21440
rect 14875 21468 14887 21471
rect 14918 21468 14924 21480
rect 14875 21440 14924 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15028 21468 15056 21508
rect 15565 21505 15577 21539
rect 15611 21536 15623 21539
rect 16206 21536 16212 21548
rect 15611 21508 16212 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16546 21536 16574 21576
rect 22554 21564 22560 21576
rect 22612 21564 22618 21616
rect 23474 21604 23480 21616
rect 22664 21576 23480 21604
rect 18417 21539 18475 21545
rect 18417 21536 18429 21539
rect 16546 21508 18429 21536
rect 18417 21505 18429 21508
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 19426 21536 19432 21548
rect 19383 21508 19432 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19352 21468 19380 21499
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 21818 21536 21824 21548
rect 20303 21508 21824 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 15028 21440 19380 21468
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 20070 21468 20076 21480
rect 19567 21440 20076 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 22002 21468 22008 21480
rect 21315 21440 22008 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 22002 21428 22008 21440
rect 22060 21428 22066 21480
rect 22664 21477 22692 21576
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 23624 21576 24058 21604
rect 23624 21564 23630 21576
rect 23198 21496 23204 21548
rect 23256 21536 23262 21548
rect 23293 21539 23351 21545
rect 23293 21536 23305 21539
rect 23256 21508 23305 21536
rect 23256 21496 23262 21508
rect 23293 21505 23305 21508
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 22465 21471 22523 21477
rect 22465 21437 22477 21471
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 25314 21468 25320 21480
rect 23615 21440 25320 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 14642 21360 14648 21412
rect 14700 21400 14706 21412
rect 15749 21403 15807 21409
rect 15749 21400 15761 21403
rect 14700 21372 15761 21400
rect 14700 21360 14706 21372
rect 15749 21369 15761 21372
rect 15795 21369 15807 21403
rect 15749 21363 15807 21369
rect 19610 21360 19616 21412
rect 19668 21400 19674 21412
rect 19668 21372 20576 21400
rect 19668 21360 19674 21372
rect 13412 21304 14412 21332
rect 18877 21335 18935 21341
rect 13412 21292 13418 21304
rect 18877 21301 18889 21335
rect 18923 21332 18935 21335
rect 20438 21332 20444 21344
rect 18923 21304 20444 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 20548 21332 20576 21372
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 20548 21304 22017 21332
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22005 21295 22063 21301
rect 22370 21292 22376 21344
rect 22428 21332 22434 21344
rect 22480 21332 22508 21431
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 22428 21304 22508 21332
rect 22428 21292 22434 21304
rect 22922 21292 22928 21344
rect 22980 21332 22986 21344
rect 23566 21332 23572 21344
rect 22980 21304 23572 21332
rect 22980 21292 22986 21304
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 8570 21088 8576 21140
rect 8628 21088 8634 21140
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 12434 21128 12440 21140
rect 9539 21100 12440 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 16264 21100 16957 21128
rect 16264 21088 16270 21100
rect 16945 21097 16957 21100
rect 16991 21128 17003 21131
rect 17034 21128 17040 21140
rect 16991 21100 17040 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 22094 21088 22100 21140
rect 22152 21128 22158 21140
rect 23934 21128 23940 21140
rect 22152 21100 23940 21128
rect 22152 21088 22158 21100
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 20625 21063 20683 21069
rect 20625 21029 20637 21063
rect 20671 21060 20683 21063
rect 21266 21060 21272 21072
rect 20671 21032 21272 21060
rect 20671 21029 20683 21032
rect 20625 21023 20683 21029
rect 21266 21020 21272 21032
rect 21324 21020 21330 21072
rect 22186 21020 22192 21072
rect 22244 21020 22250 21072
rect 22738 21020 22744 21072
rect 22796 21060 22802 21072
rect 23382 21060 23388 21072
rect 22796 21032 23388 21060
rect 22796 21020 22802 21032
rect 23382 21020 23388 21032
rect 23440 21060 23446 21072
rect 23440 21032 25268 21060
rect 23440 21020 23446 21032
rect 7101 20995 7159 21001
rect 7101 20961 7113 20995
rect 7147 20992 7159 20995
rect 9582 20992 9588 21004
rect 7147 20964 9588 20992
rect 7147 20961 7159 20964
rect 7101 20955 7159 20961
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20992 12495 20995
rect 12618 20992 12624 21004
rect 12483 20964 12624 20992
rect 12483 20961 12495 20964
rect 12437 20955 12495 20961
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 16022 20992 16028 21004
rect 15243 20964 16028 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 16022 20952 16028 20964
rect 16080 20992 16086 21004
rect 16482 20992 16488 21004
rect 16080 20964 16488 20992
rect 16080 20952 16086 20964
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 19518 20952 19524 21004
rect 19576 20992 19582 21004
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19576 20964 19993 20992
rect 19576 20952 19582 20964
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 21082 20952 21088 21004
rect 21140 20952 21146 21004
rect 21177 20995 21235 21001
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 22370 20992 22376 21004
rect 21223 20964 22376 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 23842 20952 23848 21004
rect 23900 20992 23906 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 23900 20964 25145 20992
rect 23900 20952 23906 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 6546 20884 6552 20936
rect 6604 20924 6610 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6604 20896 6837 20924
rect 6604 20884 6610 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 9858 20884 9864 20936
rect 9916 20884 9922 20936
rect 10686 20884 10692 20936
rect 10744 20884 10750 20936
rect 16574 20884 16580 20936
rect 16632 20884 16638 20936
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19760 20896 19809 20924
rect 19760 20884 19766 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19886 20884 19892 20936
rect 19944 20884 19950 20936
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 22094 20924 22100 20936
rect 21876 20896 22100 20924
rect 21876 20884 21882 20896
rect 22094 20884 22100 20896
rect 22152 20884 22158 20936
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 24946 20884 24952 20936
rect 25004 20924 25010 20936
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 25004 20896 25053 20924
rect 25004 20884 25010 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 8478 20856 8484 20868
rect 8326 20828 8484 20856
rect 8478 20816 8484 20828
rect 8536 20816 8542 20868
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 10928 20828 10977 20856
rect 10928 20816 10934 20828
rect 10965 20825 10977 20828
rect 11011 20825 11023 20859
rect 10965 20819 11023 20825
rect 11422 20816 11428 20868
rect 11480 20816 11486 20868
rect 15473 20859 15531 20865
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15746 20856 15752 20868
rect 15519 20828 15752 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 19978 20856 19984 20868
rect 19444 20828 19984 20856
rect 9950 20748 9956 20800
rect 10008 20748 10014 20800
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 14366 20788 14372 20800
rect 13504 20760 14372 20788
rect 13504 20748 13510 20760
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 19444 20797 19472 20828
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 23845 20859 23903 20865
rect 23845 20825 23857 20859
rect 23891 20856 23903 20859
rect 25130 20856 25136 20868
rect 23891 20828 25136 20856
rect 23891 20825 23903 20828
rect 23845 20819 23903 20825
rect 25130 20816 25136 20828
rect 25188 20816 25194 20868
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20757 19487 20791
rect 19429 20751 19487 20757
rect 24581 20791 24639 20797
rect 24581 20757 24593 20791
rect 24627 20788 24639 20791
rect 24854 20788 24860 20800
rect 24627 20760 24860 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 25240 20788 25268 21032
rect 24995 20760 25268 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 9548 20556 10425 20584
rect 9548 20544 9554 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 10413 20547 10471 20553
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 14734 20584 14740 20596
rect 10827 20556 14740 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 15470 20544 15476 20596
rect 15528 20544 15534 20596
rect 19334 20584 19340 20596
rect 16868 20556 19340 20584
rect 8478 20476 8484 20528
rect 8536 20476 8542 20528
rect 9766 20476 9772 20528
rect 9824 20516 9830 20528
rect 10873 20519 10931 20525
rect 10873 20516 10885 20519
rect 9824 20488 10885 20516
rect 9824 20476 9830 20488
rect 10873 20485 10885 20488
rect 10919 20485 10931 20519
rect 10873 20479 10931 20485
rect 11422 20476 11428 20528
rect 11480 20516 11486 20528
rect 13446 20516 13452 20528
rect 11480 20488 13452 20516
rect 11480 20476 11486 20488
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 14366 20476 14372 20528
rect 14424 20516 14430 20528
rect 16574 20516 16580 20528
rect 14424 20488 16580 20516
rect 14424 20476 14430 20488
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 7742 20448 7748 20460
rect 6604 20420 7748 20448
rect 6604 20408 6610 20420
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 9640 20420 11008 20448
rect 9640 20408 9646 20420
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8570 20380 8576 20392
rect 8067 20352 8576 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10980 20389 11008 20420
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 16868 20457 16896 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 22094 20544 22100 20596
rect 22152 20544 22158 20596
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 17126 20476 17132 20528
rect 17184 20476 17190 20528
rect 17402 20476 17408 20528
rect 17460 20516 17466 20528
rect 17460 20488 17618 20516
rect 17460 20476 17466 20488
rect 23566 20476 23572 20528
rect 23624 20516 23630 20528
rect 23624 20488 24334 20516
rect 23624 20476 23630 20488
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 9769 20383 9827 20389
rect 9769 20380 9781 20383
rect 9732 20352 9781 20380
rect 9732 20340 9738 20352
rect 9769 20349 9781 20352
rect 9815 20349 9827 20383
rect 9769 20343 9827 20349
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13354 20380 13360 20392
rect 13035 20352 13360 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13354 20340 13360 20352
rect 13412 20340 13418 20392
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 15580 20312 15608 20343
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 18138 20380 18144 20392
rect 17552 20352 18144 20380
rect 17552 20340 17558 20352
rect 18138 20340 18144 20352
rect 18196 20340 18202 20392
rect 18598 20340 18604 20392
rect 18656 20340 18662 20392
rect 20088 20380 20116 20411
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 20220 20420 22293 20448
rect 20220 20408 20226 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22554 20408 22560 20460
rect 22612 20448 22618 20460
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22612 20420 22937 20448
rect 22612 20408 22618 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 21174 20380 21180 20392
rect 20088 20352 21180 20380
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20380 21327 20383
rect 22094 20380 22100 20392
rect 21315 20352 22100 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 22094 20340 22100 20352
rect 22152 20340 22158 20392
rect 22738 20340 22744 20392
rect 22796 20380 22802 20392
rect 23569 20383 23627 20389
rect 23569 20380 23581 20383
rect 22796 20352 23581 20380
rect 22796 20340 22802 20352
rect 23569 20349 23581 20352
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25130 20380 25136 20392
rect 23891 20352 25136 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 14476 20284 15608 20312
rect 14476 20256 14504 20284
rect 14458 20204 14464 20256
rect 14516 20204 14522 20256
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 17770 20244 17776 20256
rect 15059 20216 17776 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 22646 20204 22652 20256
rect 22704 20244 22710 20256
rect 22741 20247 22799 20253
rect 22741 20244 22753 20247
rect 22704 20216 22753 20244
rect 22704 20204 22710 20216
rect 22741 20213 22753 20216
rect 22787 20213 22799 20247
rect 22741 20207 22799 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 9214 20040 9220 20052
rect 8444 20012 9220 20040
rect 8444 20000 8450 20012
rect 9214 20000 9220 20012
rect 9272 20040 9278 20052
rect 9382 20043 9440 20049
rect 9382 20040 9394 20043
rect 9272 20012 9394 20040
rect 9272 20000 9278 20012
rect 9382 20009 9394 20012
rect 9428 20009 9440 20043
rect 9382 20003 9440 20009
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 13906 20040 13912 20052
rect 11379 20012 13912 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15804 20012 16037 20040
rect 15804 20000 15810 20012
rect 16025 20009 16037 20012
rect 16071 20040 16083 20043
rect 16114 20040 16120 20052
rect 16071 20012 16120 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 19334 20040 19340 20052
rect 16531 20012 19340 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 20162 20040 20168 20052
rect 19444 20012 20168 20040
rect 19444 19972 19472 20012
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 23566 20040 23572 20052
rect 20864 20012 23572 20040
rect 20864 20000 20870 20012
rect 16546 19944 19472 19972
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 7892 19876 9137 19904
rect 7892 19864 7898 19876
rect 9125 19873 9137 19876
rect 9171 19904 9183 19907
rect 10686 19904 10692 19916
rect 9171 19876 10692 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 12768 19876 14289 19904
rect 12768 19864 12774 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 14918 19864 14924 19916
rect 14976 19904 14982 19916
rect 16546 19904 16574 19944
rect 14976 19876 16574 19904
rect 14976 19864 14982 19876
rect 17126 19864 17132 19916
rect 17184 19904 17190 19916
rect 18049 19907 18107 19913
rect 18049 19904 18061 19907
rect 17184 19876 18061 19904
rect 17184 19864 17190 19876
rect 18049 19873 18061 19876
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 19889 19907 19947 19913
rect 18196 19876 19840 19904
rect 18196 19864 18202 19876
rect 16666 19796 16672 19848
rect 16724 19796 16730 19848
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17920 19808 17969 19836
rect 17920 19796 17926 19808
rect 17957 19805 17969 19808
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19150 19836 19156 19848
rect 18923 19808 19156 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 8478 19728 8484 19780
rect 8536 19768 8542 19780
rect 11422 19768 11428 19780
rect 8536 19740 9890 19768
rect 10796 19740 11428 19768
rect 8536 19728 8542 19740
rect 9784 19700 9812 19740
rect 10796 19700 10824 19740
rect 11422 19728 11428 19740
rect 11480 19728 11486 19780
rect 14553 19771 14611 19777
rect 14553 19737 14565 19771
rect 14599 19737 14611 19771
rect 16574 19768 16580 19780
rect 15778 19740 16580 19768
rect 14553 19731 14611 19737
rect 9784 19672 10824 19700
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 11882 19700 11888 19712
rect 11839 19672 11888 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 14568 19700 14596 19731
rect 16574 19728 16580 19740
rect 16632 19768 16638 19780
rect 17034 19768 17040 19780
rect 16632 19740 17040 19768
rect 16632 19728 16638 19740
rect 17034 19728 17040 19740
rect 17092 19768 17098 19780
rect 17402 19768 17408 19780
rect 17092 19740 17408 19768
rect 17092 19728 17098 19740
rect 17402 19728 17408 19740
rect 17460 19728 17466 19780
rect 19242 19768 19248 19780
rect 17512 19740 19248 19768
rect 15930 19700 15936 19712
rect 14568 19672 15936 19700
rect 15930 19660 15936 19672
rect 15988 19660 15994 19712
rect 17512 19709 17540 19740
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19669 17555 19703
rect 17497 19663 17555 19669
rect 17862 19660 17868 19712
rect 17920 19660 17926 19712
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 19150 19700 19156 19712
rect 18739 19672 19156 19700
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 19812 19700 19840 19876
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20254 19904 20260 19916
rect 19935 19876 20260 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20254 19864 20260 19876
rect 20312 19904 20318 19916
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 20312 19876 22109 19904
rect 20312 19864 20318 19876
rect 22097 19873 22109 19876
rect 22143 19904 22155 19907
rect 22738 19904 22744 19916
rect 22143 19876 22744 19904
rect 22143 19873 22155 19876
rect 22097 19867 22155 19873
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 23492 19836 23520 20012
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 23842 20000 23848 20052
rect 23900 20000 23906 20052
rect 24026 19836 24032 19848
rect 23492 19822 24032 19836
rect 23506 19808 24032 19822
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 20548 19740 20654 19768
rect 21652 19740 22385 19768
rect 20548 19700 20576 19740
rect 20806 19700 20812 19712
rect 19812 19672 20812 19700
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 20898 19660 20904 19712
rect 20956 19700 20962 19712
rect 21652 19709 21680 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 22373 19731 22431 19737
rect 21637 19703 21695 19709
rect 21637 19700 21649 19703
rect 20956 19672 21649 19700
rect 20956 19660 20962 19672
rect 21637 19669 21649 19672
rect 21683 19669 21695 19703
rect 21637 19663 21695 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 11480 19468 13032 19496
rect 11480 19456 11486 19468
rect 8478 19428 8484 19440
rect 8050 19400 8484 19428
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 12710 19428 12716 19440
rect 12452 19400 12716 19428
rect 9122 19320 9128 19372
rect 9180 19320 9186 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 10042 19360 10048 19372
rect 9263 19332 10048 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 12452 19369 12480 19400
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 13004 19428 13032 19468
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13780 19468 14044 19496
rect 13780 19456 13786 19468
rect 14016 19428 14044 19468
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14185 19499 14243 19505
rect 14185 19496 14197 19499
rect 14148 19468 14197 19496
rect 14148 19456 14154 19468
rect 14185 19465 14197 19468
rect 14231 19465 14243 19499
rect 14185 19459 14243 19465
rect 14918 19456 14924 19508
rect 14976 19456 14982 19508
rect 15565 19499 15623 19505
rect 15565 19465 15577 19499
rect 15611 19496 15623 19499
rect 15611 19468 16574 19496
rect 15611 19465 15623 19468
rect 15565 19459 15623 19465
rect 15933 19431 15991 19437
rect 15933 19428 15945 19431
rect 13004 19400 13202 19428
rect 14016 19400 15945 19428
rect 15933 19397 15945 19400
rect 15979 19397 15991 19431
rect 15933 19391 15991 19397
rect 16025 19431 16083 19437
rect 16025 19397 16037 19431
rect 16071 19428 16083 19431
rect 16298 19428 16304 19440
rect 16071 19400 16304 19428
rect 16071 19397 16083 19400
rect 16025 19391 16083 19397
rect 16298 19388 16304 19400
rect 16356 19388 16362 19440
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11756 19332 11897 19360
rect 11756 19320 11762 19332
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 15102 19320 15108 19372
rect 15160 19320 15166 19372
rect 16546 19360 16574 19468
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 16816 19468 17049 19496
rect 16816 19456 16822 19468
rect 17037 19465 17049 19468
rect 17083 19465 17095 19499
rect 17037 19459 17095 19465
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 17368 19468 17509 19496
rect 17368 19456 17374 19468
rect 17497 19465 17509 19468
rect 17543 19465 17555 19499
rect 17497 19459 17555 19465
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 16850 19388 16856 19440
rect 16908 19428 16914 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 16908 19400 17417 19428
rect 16908 19388 16914 19400
rect 17405 19397 17417 19400
rect 17451 19397 17463 19431
rect 18690 19428 18696 19440
rect 17405 19391 17463 19397
rect 17512 19400 18696 19428
rect 17512 19360 17540 19400
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 18984 19428 19012 19459
rect 20438 19456 20444 19508
rect 20496 19456 20502 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 22189 19499 22247 19505
rect 22189 19496 22201 19499
rect 20864 19468 22201 19496
rect 20864 19456 20870 19468
rect 22189 19465 22201 19468
rect 22235 19465 22247 19499
rect 22189 19459 22247 19465
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 24578 19496 24584 19508
rect 22695 19468 24584 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 23566 19428 23572 19440
rect 18984 19400 23572 19428
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23661 19431 23719 19437
rect 23661 19397 23673 19431
rect 23707 19428 23719 19431
rect 23750 19428 23756 19440
rect 23707 19400 23756 19428
rect 23707 19397 23719 19400
rect 23661 19391 23719 19397
rect 23750 19388 23756 19400
rect 23808 19388 23814 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 16546 19332 17540 19360
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 17828 19332 19165 19360
rect 17828 19320 17834 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 22557 19363 22615 19369
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19292 6978 19304
rect 7374 19292 7380 19304
rect 6972 19264 7380 19292
rect 6972 19252 6978 19264
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 14458 19292 14464 19304
rect 12759 19264 14464 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 8570 19184 8576 19236
rect 8628 19224 8634 19236
rect 9324 19224 9352 19255
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 16114 19252 16120 19304
rect 16172 19252 16178 19304
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 20625 19295 20683 19301
rect 20625 19261 20637 19295
rect 20671 19292 20683 19295
rect 20898 19292 20904 19304
rect 20671 19264 20904 19292
rect 20671 19261 20683 19264
rect 20625 19255 20683 19261
rect 8628 19196 9352 19224
rect 8628 19184 8634 19196
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 17604 19224 17632 19255
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 22572 19292 22600 19323
rect 22830 19320 22836 19372
rect 22888 19360 22894 19372
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 22888 19332 23397 19360
rect 22888 19320 22894 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 21499 19264 22600 19292
rect 22741 19295 22799 19301
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 22741 19261 22753 19295
rect 22787 19292 22799 19295
rect 22922 19292 22928 19304
rect 22787 19264 22928 19292
rect 22787 19261 22799 19264
rect 22741 19255 22799 19261
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 17368 19196 17632 19224
rect 17368 19184 17374 19196
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 23290 19224 23296 19236
rect 22336 19196 23296 19224
rect 22336 19184 22342 19196
rect 23290 19184 23296 19196
rect 23348 19184 23354 19236
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 9214 19156 9220 19168
rect 8352 19128 9220 19156
rect 8352 19116 8358 19128
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 23382 19156 23388 19168
rect 21140 19128 23388 19156
rect 21140 19116 21146 19128
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8386 18912 8392 18964
rect 8444 18912 8450 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10778 18952 10784 18964
rect 10091 18924 10784 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 16666 18952 16672 18964
rect 11563 18924 16672 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 21082 18952 21088 18964
rect 19260 18924 21088 18952
rect 10410 18844 10416 18896
rect 10468 18884 10474 18896
rect 11606 18884 11612 18896
rect 10468 18856 11612 18884
rect 10468 18844 10474 18856
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8294 18816 8300 18828
rect 6963 18788 8300 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 10612 18825 10640 18856
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 18782 18884 18788 18896
rect 16546 18856 18788 18884
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 10928 18788 12081 18816
rect 10928 18776 10934 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 12069 18779 12127 18785
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6604 18720 6653 18748
rect 6604 18708 6610 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 8478 18748 8484 18760
rect 8050 18720 8484 18748
rect 6641 18711 6699 18717
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10410 18748 10416 18760
rect 10008 18720 10416 18748
rect 10008 18708 10014 18720
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12492 18720 12909 18748
rect 12492 18708 12498 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16546 18748 16574 18856
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17770 18816 17776 18828
rect 17451 18788 17776 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 16255 18720 16574 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 16908 18720 17141 18748
rect 16908 18708 16914 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17236 18748 17264 18776
rect 17494 18748 17500 18760
rect 17236 18720 17500 18748
rect 17129 18711 17187 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 8220 18652 11897 18680
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 8220 18612 8248 18652
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 11885 18643 11943 18649
rect 11977 18683 12035 18689
rect 11977 18649 11989 18683
rect 12023 18680 12035 18683
rect 12526 18680 12532 18692
rect 12023 18652 12532 18680
rect 12023 18649 12035 18652
rect 11977 18643 12035 18649
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 19260 18680 19288 18924
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 21174 18912 21180 18964
rect 21232 18952 21238 18964
rect 21637 18955 21695 18961
rect 21637 18952 21649 18955
rect 21232 18924 21649 18952
rect 21232 18912 21238 18924
rect 21637 18921 21649 18924
rect 21683 18921 21695 18955
rect 21637 18915 21695 18921
rect 20257 18887 20315 18893
rect 20257 18853 20269 18887
rect 20303 18884 20315 18887
rect 22554 18884 22560 18896
rect 20303 18856 22560 18884
rect 20303 18853 20315 18856
rect 20257 18847 20315 18853
rect 22554 18844 22560 18856
rect 22612 18844 22618 18896
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19392 18788 21864 18816
rect 19392 18776 19398 18788
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 12728 18652 19288 18680
rect 19628 18680 19656 18711
rect 20438 18708 20444 18760
rect 20496 18708 20502 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21450 18748 21456 18760
rect 21131 18720 21456 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21836 18757 21864 18788
rect 23842 18776 23848 18828
rect 23900 18776 23906 18828
rect 21821 18751 21879 18757
rect 21821 18717 21833 18751
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 23624 18720 24777 18748
rect 23624 18708 23630 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 21910 18680 21916 18692
rect 19628 18652 21916 18680
rect 7616 18584 8248 18612
rect 7616 18572 7622 18584
rect 10502 18572 10508 18624
rect 10560 18572 10566 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 12728 18612 12756 18652
rect 21910 18640 21916 18652
rect 21968 18640 21974 18692
rect 22002 18640 22008 18692
rect 22060 18680 22066 18692
rect 25498 18680 25504 18692
rect 22060 18652 25504 18680
rect 22060 18640 22066 18652
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 10928 18584 12756 18612
rect 10928 18572 10934 18584
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 16025 18615 16083 18621
rect 16025 18612 16037 18615
rect 15712 18584 16037 18612
rect 15712 18572 15718 18584
rect 16025 18581 16037 18584
rect 16071 18581 16083 18615
rect 16025 18575 16083 18581
rect 16758 18572 16764 18624
rect 16816 18572 16822 18624
rect 18782 18572 18788 18624
rect 18840 18612 18846 18624
rect 19429 18615 19487 18621
rect 19429 18612 19441 18615
rect 18840 18584 19441 18612
rect 18840 18572 18846 18584
rect 19429 18581 19441 18584
rect 19475 18581 19487 18615
rect 19429 18575 19487 18581
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 20901 18615 20959 18621
rect 20901 18612 20913 18615
rect 20772 18584 20913 18612
rect 20772 18572 20778 18584
rect 20901 18581 20913 18584
rect 20947 18581 20959 18615
rect 20901 18575 20959 18581
rect 24118 18572 24124 18624
rect 24176 18612 24182 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 24176 18584 24593 18612
rect 24176 18572 24182 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 9582 18408 9588 18420
rect 9447 18380 9588 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 10318 18368 10324 18420
rect 10376 18368 10382 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 13725 18411 13783 18417
rect 13725 18408 13737 18411
rect 10560 18380 13737 18408
rect 10560 18368 10566 18380
rect 13725 18377 13737 18380
rect 13771 18377 13783 18411
rect 13725 18371 13783 18377
rect 14093 18411 14151 18417
rect 14093 18377 14105 18411
rect 14139 18408 14151 18411
rect 17218 18408 17224 18420
rect 14139 18380 17224 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 8478 18300 8484 18352
rect 8536 18300 8542 18352
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 9272 18312 10456 18340
rect 9272 18300 9278 18312
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 10192 18244 10241 18272
rect 10192 18232 10198 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 6546 18164 6552 18216
rect 6604 18204 6610 18216
rect 10428 18213 10456 18312
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 12802 18340 12808 18352
rect 10836 18312 12808 18340
rect 10836 18300 10842 18312
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 13265 18343 13323 18349
rect 13265 18309 13277 18343
rect 13311 18340 13323 18343
rect 14108 18340 14136 18371
rect 17218 18368 17224 18380
rect 17276 18408 17282 18420
rect 22002 18408 22008 18420
rect 17276 18380 22008 18408
rect 17276 18368 17282 18380
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 25682 18408 25688 18420
rect 22664 18380 25688 18408
rect 13311 18312 14136 18340
rect 13311 18309 13323 18312
rect 13265 18303 13323 18309
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 22664 18349 22692 18380
rect 25682 18368 25688 18380
rect 25740 18368 25746 18420
rect 22649 18343 22707 18349
rect 17092 18312 17618 18340
rect 17092 18300 17098 18312
rect 22649 18309 22661 18343
rect 22695 18309 22707 18343
rect 22649 18303 22707 18309
rect 23569 18343 23627 18349
rect 23569 18309 23581 18343
rect 23615 18340 23627 18343
rect 23658 18340 23664 18352
rect 23615 18312 23664 18340
rect 23615 18309 23627 18312
rect 23569 18303 23627 18309
rect 23658 18300 23664 18312
rect 23716 18300 23722 18352
rect 24026 18300 24032 18352
rect 24084 18300 24090 18352
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 12584 18244 14320 18272
rect 12584 18232 12590 18244
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 6604 18176 7665 18204
rect 6604 18164 6610 18176
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18204 7987 18207
rect 10413 18207 10471 18213
rect 7975 18176 9812 18204
rect 7975 18173 7987 18176
rect 7929 18167 7987 18173
rect 7668 18068 7696 18167
rect 9582 18136 9588 18148
rect 8956 18108 9588 18136
rect 8956 18068 8984 18108
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 7668 18040 8984 18068
rect 9784 18068 9812 18176
rect 10413 18173 10425 18207
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 14182 18164 14188 18216
rect 14240 18164 14246 18216
rect 14292 18213 14320 18244
rect 16482 18232 16488 18284
rect 16540 18272 16546 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16540 18244 16865 18272
rect 16540 18232 16546 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 19300 18244 20545 18272
rect 19300 18232 19306 18244
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16448 18176 17141 18204
rect 16448 18164 16454 18176
rect 17129 18173 17141 18176
rect 17175 18204 17187 18207
rect 18598 18204 18604 18216
rect 17175 18176 18604 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 21192 18204 21220 18235
rect 22738 18232 22744 18284
rect 22796 18272 22802 18284
rect 23293 18275 23351 18281
rect 23293 18272 23305 18275
rect 22796 18244 23305 18272
rect 22796 18232 22802 18244
rect 23293 18241 23305 18244
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 24210 18204 24216 18216
rect 21192 18176 24216 18204
rect 24210 18164 24216 18176
rect 24268 18164 24274 18216
rect 25314 18164 25320 18216
rect 25372 18164 25378 18216
rect 9861 18139 9919 18145
rect 9861 18105 9873 18139
rect 9907 18136 9919 18139
rect 15102 18136 15108 18148
rect 9907 18108 15108 18136
rect 9907 18105 9919 18108
rect 9861 18099 9919 18105
rect 15102 18096 15108 18108
rect 15160 18096 15166 18148
rect 20349 18139 20407 18145
rect 20349 18105 20361 18139
rect 20395 18136 20407 18139
rect 23290 18136 23296 18148
rect 20395 18108 23296 18136
rect 20395 18105 20407 18108
rect 20349 18099 20407 18105
rect 23290 18096 23296 18108
rect 23348 18096 23354 18148
rect 10778 18068 10784 18080
rect 9784 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 18598 18028 18604 18080
rect 18656 18028 18662 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20956 18040 21005 18068
rect 20956 18028 20962 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 20993 18031 21051 18037
rect 22738 18028 22744 18080
rect 22796 18028 22802 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7708 17836 7849 17864
rect 7708 17824 7714 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 12526 17864 12532 17876
rect 7837 17827 7895 17833
rect 11072 17836 12532 17864
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7800 17700 8401 17728
rect 7800 17688 7806 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9732 17700 10057 17728
rect 9732 17688 9738 17700
rect 10045 17697 10057 17700
rect 10091 17728 10103 17731
rect 11072 17728 11100 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12894 17864 12900 17876
rect 12676 17836 12900 17864
rect 12676 17824 12682 17836
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 13538 17824 13544 17876
rect 13596 17864 13602 17876
rect 14274 17864 14280 17876
rect 13596 17836 14280 17864
rect 13596 17824 13602 17836
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 20162 17824 20168 17876
rect 20220 17864 20226 17876
rect 21177 17867 21235 17873
rect 21177 17864 21189 17867
rect 20220 17836 21189 17864
rect 20220 17824 20226 17836
rect 21177 17833 21189 17836
rect 21223 17833 21235 17867
rect 21177 17827 21235 17833
rect 12802 17796 12808 17808
rect 10091 17700 11100 17728
rect 11164 17768 12808 17796
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 7374 17620 7380 17672
rect 7432 17620 7438 17672
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17660 9367 17663
rect 9398 17660 9404 17672
rect 9355 17632 9404 17660
rect 9355 17629 9367 17632
rect 9309 17623 9367 17629
rect 9398 17620 9404 17632
rect 9456 17620 9462 17672
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9640 17632 9781 17660
rect 9640 17620 9646 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 11164 17646 11192 17768
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 25774 17796 25780 17808
rect 22020 17768 25780 17796
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11664 17700 11805 17728
rect 11664 17688 11670 17700
rect 11793 17697 11805 17700
rect 11839 17728 11851 17731
rect 12250 17728 12256 17740
rect 11839 17700 12256 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12768 17700 13093 17728
rect 12768 17688 12774 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 18414 17688 18420 17740
rect 18472 17688 18478 17740
rect 18598 17688 18604 17740
rect 18656 17688 18662 17740
rect 12345 17663 12403 17669
rect 9769 17623 9827 17629
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12391 17632 13216 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 9214 17592 9220 17604
rect 8251 17564 9220 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 8297 17527 8355 17533
rect 8297 17493 8309 17527
rect 8343 17524 8355 17527
rect 9950 17524 9956 17536
rect 8343 17496 9956 17524
rect 8343 17493 8355 17496
rect 8297 17487 8355 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 10226 17484 10232 17536
rect 10284 17524 10290 17536
rect 10962 17524 10968 17536
rect 10284 17496 10968 17524
rect 10284 17484 10290 17496
rect 10962 17484 10968 17496
rect 11020 17524 11026 17536
rect 12360 17524 12388 17623
rect 13188 17592 13216 17632
rect 13630 17620 13636 17672
rect 13688 17620 13694 17672
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17660 15899 17663
rect 16114 17660 16120 17672
rect 15887 17632 16120 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17660 16911 17663
rect 16942 17660 16948 17672
rect 16899 17632 16948 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 22020 17669 22048 17768
rect 25774 17756 25780 17768
rect 25832 17756 25838 17808
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 25041 17731 25099 17737
rect 25041 17728 25053 17731
rect 25004 17700 25053 17728
rect 25004 17688 25010 17700
rect 25041 17697 25053 17700
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 22649 17663 22707 17669
rect 22649 17660 22661 17663
rect 22612 17632 22661 17660
rect 22612 17620 22618 17632
rect 22649 17629 22661 17632
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 17218 17592 17224 17604
rect 13188 17564 17224 17592
rect 17218 17552 17224 17564
rect 17276 17592 17282 17604
rect 17678 17592 17684 17604
rect 17276 17564 17684 17592
rect 17276 17552 17282 17564
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 18325 17595 18383 17601
rect 18325 17561 18337 17595
rect 18371 17592 18383 17595
rect 18874 17592 18880 17604
rect 18371 17564 18880 17592
rect 18371 17561 18383 17564
rect 18325 17555 18383 17561
rect 18874 17552 18880 17564
rect 18932 17552 18938 17604
rect 18966 17552 18972 17604
rect 19024 17592 19030 17604
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 19024 17564 19717 17592
rect 19024 17552 19030 17564
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 20990 17592 20996 17604
rect 20930 17564 20996 17592
rect 19705 17555 19763 17561
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 21818 17592 21824 17604
rect 21100 17564 21824 17592
rect 11020 17496 12388 17524
rect 11020 17484 11026 17496
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 15194 17524 15200 17536
rect 12676 17496 15200 17524
rect 12676 17484 12682 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 16669 17527 16727 17533
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 16850 17524 16856 17536
rect 16715 17496 16856 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 17957 17527 18015 17533
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 21100 17524 21128 17564
rect 21818 17552 21824 17564
rect 21876 17552 21882 17604
rect 18003 17496 21128 17524
rect 22097 17527 22155 17533
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22646 17524 22652 17536
rect 22143 17496 22652 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22646 17484 22652 17496
rect 22704 17484 22710 17536
rect 22830 17484 22836 17536
rect 22888 17524 22894 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 22888 17496 24593 17524
rect 22888 17484 22894 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7432 17292 8033 17320
rect 7432 17280 7438 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9033 17323 9091 17329
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9306 17320 9312 17332
rect 9079 17292 9312 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 11790 17320 11796 17332
rect 9508 17292 11796 17320
rect 9508 17252 9536 17292
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12345 17323 12403 17329
rect 12345 17289 12357 17323
rect 12391 17320 12403 17323
rect 12434 17320 12440 17332
rect 12391 17292 12440 17320
rect 12391 17289 12403 17292
rect 12345 17283 12403 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13630 17320 13636 17332
rect 13219 17292 13636 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 16482 17320 16488 17332
rect 14476 17292 16488 17320
rect 6886 17224 9536 17252
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 6886 17184 6914 17224
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 9640 17224 10977 17252
rect 9640 17212 9646 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 14182 17252 14188 17264
rect 10965 17215 11023 17221
rect 12452 17224 14188 17252
rect 3568 17156 6914 17184
rect 3568 17144 3574 17156
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 8720 17156 9628 17184
rect 8720 17144 8726 17156
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 3384 17088 8125 17116
rect 3384 17076 3390 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8938 17116 8944 17128
rect 8343 17088 8944 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9600 17125 9628 17156
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 12452 17193 12480 17224
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 11664 17156 12449 17184
rect 11664 17144 11670 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13630 17184 13636 17196
rect 13311 17156 13636 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 14476 17193 14504 17292
rect 16482 17280 16488 17292
rect 16540 17320 16546 17332
rect 16574 17320 16580 17332
rect 16540 17292 16580 17320
rect 16540 17280 16546 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 18877 17323 18935 17329
rect 18877 17289 18889 17323
rect 18923 17320 18935 17323
rect 20438 17320 20444 17332
rect 18923 17292 20444 17320
rect 18923 17289 18935 17292
rect 18877 17283 18935 17289
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 21177 17323 21235 17329
rect 21177 17289 21189 17323
rect 21223 17320 21235 17323
rect 24302 17320 24308 17332
rect 21223 17292 24308 17320
rect 21223 17289 21235 17292
rect 21177 17283 21235 17289
rect 24302 17280 24308 17292
rect 24360 17280 24366 17332
rect 15962 17224 16712 17252
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17153 14519 17187
rect 16684 17184 16712 17224
rect 16942 17212 16948 17264
rect 17000 17212 17006 17264
rect 18233 17255 18291 17261
rect 18233 17221 18245 17255
rect 18279 17252 18291 17255
rect 18506 17252 18512 17264
rect 18279 17224 18512 17252
rect 18279 17221 18291 17224
rect 18233 17215 18291 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 18690 17212 18696 17264
rect 18748 17252 18754 17264
rect 23293 17255 23351 17261
rect 18748 17224 20024 17252
rect 18748 17212 18754 17224
rect 17034 17184 17040 17196
rect 16684 17156 17040 17184
rect 14461 17147 14519 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 19996 17193 20024 17224
rect 20088 17224 21404 17252
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9456 17088 9505 17116
rect 9456 17076 9462 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 12894 17116 12900 17128
rect 12575 17088 12900 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13354 17076 13360 17128
rect 13412 17076 13418 17128
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 15470 17116 15476 17128
rect 14783 17088 15476 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 19076 17116 19104 17147
rect 20088 17116 20116 17224
rect 21082 17144 21088 17196
rect 21140 17144 21146 17196
rect 21376 17125 21404 17224
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 24854 17252 24860 17264
rect 23339 17224 24860 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 22186 17144 22192 17196
rect 22244 17144 22250 17196
rect 24118 17144 24124 17196
rect 24176 17144 24182 17196
rect 25314 17184 25320 17196
rect 24228 17156 25320 17184
rect 16080 17088 19104 17116
rect 19168 17088 20116 17116
rect 21361 17119 21419 17125
rect 16080 17076 16086 17088
rect 7466 17008 7472 17060
rect 7524 17048 7530 17060
rect 7653 17051 7711 17057
rect 7653 17048 7665 17051
rect 7524 17020 7665 17048
rect 7524 17008 7530 17020
rect 7653 17017 7665 17020
rect 7699 17017 7711 17051
rect 7653 17011 7711 17017
rect 11977 17051 12035 17057
rect 11977 17017 11989 17051
rect 12023 17048 12035 17051
rect 12618 17048 12624 17060
rect 12023 17020 12624 17048
rect 12023 17017 12035 17020
rect 11977 17011 12035 17017
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 15930 17008 15936 17060
rect 15988 17048 15994 17060
rect 16209 17051 16267 17057
rect 16209 17048 16221 17051
rect 15988 17020 16221 17048
rect 15988 17008 15994 17020
rect 16209 17017 16221 17020
rect 16255 17017 16267 17051
rect 16209 17011 16267 17017
rect 17126 17008 17132 17060
rect 17184 17008 17190 17060
rect 19168 17048 19196 17088
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 24228 17116 24256 17156
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 21407 17088 24256 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 24762 17076 24768 17128
rect 24820 17076 24826 17128
rect 17328 17020 19196 17048
rect 19797 17051 19855 17057
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 15378 16980 15384 16992
rect 12851 16952 15384 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 16390 16940 16396 16992
rect 16448 16980 16454 16992
rect 17328 16980 17356 17020
rect 19797 17017 19809 17051
rect 19843 17048 19855 17051
rect 22002 17048 22008 17060
rect 19843 17020 22008 17048
rect 19843 17017 19855 17020
rect 19797 17011 19855 17017
rect 22002 17008 22008 17020
rect 22060 17008 22066 17060
rect 22462 17008 22468 17060
rect 22520 17048 22526 17060
rect 22646 17048 22652 17060
rect 22520 17020 22652 17048
rect 22520 17008 22526 17020
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 16448 16952 17356 16980
rect 16448 16940 16454 16952
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18012 16952 18337 16980
rect 18012 16940 18018 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 20438 16940 20444 16992
rect 20496 16980 20502 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20496 16952 20729 16980
rect 20496 16940 20502 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 24026 16940 24032 16992
rect 24084 16980 24090 16992
rect 24762 16980 24768 16992
rect 24084 16952 24768 16980
rect 24084 16940 24090 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 9030 16776 9036 16788
rect 8536 16748 9036 16776
rect 8536 16736 8542 16748
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 12710 16776 12716 16788
rect 11900 16748 12716 16776
rect 9490 16600 9496 16652
rect 9548 16640 9554 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 9548 16612 10977 16640
rect 9548 16600 9554 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 11900 16640 11928 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 14090 16776 14096 16788
rect 13464 16748 14096 16776
rect 11839 16612 11928 16640
rect 12069 16643 12127 16649
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 13464 16640 13492 16748
rect 14090 16736 14096 16748
rect 14148 16776 14154 16788
rect 15102 16776 15108 16788
rect 14148 16748 15108 16776
rect 14148 16736 14154 16748
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 17494 16776 17500 16788
rect 17092 16748 17500 16776
rect 17092 16736 17098 16748
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 24765 16779 24823 16785
rect 24765 16776 24777 16779
rect 21140 16748 24777 16776
rect 21140 16736 21146 16748
rect 24765 16745 24777 16748
rect 24811 16745 24823 16779
rect 24765 16739 24823 16745
rect 14734 16668 14740 16720
rect 14792 16708 14798 16720
rect 17954 16708 17960 16720
rect 14792 16680 17960 16708
rect 14792 16668 14798 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 15105 16643 15163 16649
rect 15105 16640 15117 16643
rect 12115 16612 13492 16640
rect 13556 16612 15117 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 9030 16572 9036 16584
rect 7524 16544 9036 16572
rect 7524 16532 7530 16544
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 10781 16507 10839 16513
rect 10781 16473 10793 16507
rect 10827 16504 10839 16507
rect 11422 16504 11428 16516
rect 10827 16476 11428 16504
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 12802 16464 12808 16516
rect 12860 16464 12866 16516
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 8904 16408 10425 16436
rect 8904 16396 8910 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11146 16436 11152 16448
rect 10919 16408 11152 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13556 16445 13584 16612
rect 15105 16609 15117 16612
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 16206 16600 16212 16652
rect 16264 16600 16270 16652
rect 16298 16600 16304 16652
rect 16356 16600 16362 16652
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 18325 16643 18383 16649
rect 18325 16640 18337 16643
rect 16632 16612 18337 16640
rect 16632 16600 16638 16612
rect 18325 16609 18337 16612
rect 18371 16640 18383 16643
rect 19426 16640 19432 16652
rect 18371 16612 19432 16640
rect 18371 16609 18383 16612
rect 18325 16603 18383 16609
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 20254 16600 20260 16652
rect 20312 16600 20318 16652
rect 16022 16572 16028 16584
rect 14568 16544 16028 16572
rect 14568 16445 14596 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 17862 16572 17868 16584
rect 16546 16544 17868 16572
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15013 16507 15071 16513
rect 15013 16504 15025 16507
rect 14884 16476 15025 16504
rect 14884 16464 14890 16476
rect 15013 16473 15025 16476
rect 15059 16473 15071 16507
rect 15013 16467 15071 16473
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13504 16408 13553 16436
rect 13504 16396 13510 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 13541 16399 13599 16405
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 14921 16439 14979 16445
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 15654 16436 15660 16448
rect 14967 16408 15660 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 16546 16436 16574 16544
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 20438 16572 20444 16584
rect 19852 16544 20444 16572
rect 19852 16532 19858 16544
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 17218 16464 17224 16516
rect 17276 16504 17282 16516
rect 17497 16507 17555 16513
rect 17497 16504 17509 16507
rect 17276 16476 17509 16504
rect 17276 16464 17282 16476
rect 17497 16473 17509 16476
rect 17543 16504 17555 16507
rect 19429 16507 19487 16513
rect 19429 16504 19441 16507
rect 17543 16476 19441 16504
rect 17543 16473 17555 16476
rect 17497 16467 17555 16473
rect 17788 16448 17816 16476
rect 19429 16473 19441 16476
rect 19475 16473 19487 16507
rect 19429 16467 19487 16473
rect 20162 16464 20168 16516
rect 20220 16504 20226 16516
rect 21008 16504 21036 16535
rect 21082 16532 21088 16584
rect 21140 16572 21146 16584
rect 21450 16572 21456 16584
rect 21140 16544 21456 16572
rect 21140 16532 21146 16544
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16572 21695 16575
rect 22278 16572 22284 16584
rect 21683 16544 22284 16572
rect 21683 16541 21695 16544
rect 21637 16535 21695 16541
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22649 16575 22707 16581
rect 22649 16572 22661 16575
rect 22428 16544 22661 16572
rect 22428 16532 22434 16544
rect 22649 16541 22661 16544
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22094 16504 22100 16516
rect 20220 16476 20852 16504
rect 21008 16476 22100 16504
rect 20220 16464 20226 16476
rect 15795 16408 16574 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 17770 16396 17776 16448
rect 17828 16396 17834 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 20530 16436 20536 16448
rect 19392 16408 20536 16436
rect 19392 16396 19398 16408
rect 20530 16396 20536 16408
rect 20588 16396 20594 16448
rect 20824 16445 20852 16476
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 23845 16507 23903 16513
rect 23845 16473 23857 16507
rect 23891 16504 23903 16507
rect 24854 16504 24860 16516
rect 23891 16476 24860 16504
rect 23891 16473 23903 16476
rect 23845 16467 23903 16473
rect 24854 16464 24860 16476
rect 24912 16464 24918 16516
rect 20809 16439 20867 16445
rect 20809 16405 20821 16439
rect 20855 16405 20867 16439
rect 20809 16399 20867 16405
rect 21453 16439 21511 16445
rect 21453 16405 21465 16439
rect 21499 16436 21511 16439
rect 21542 16436 21548 16448
rect 21499 16408 21548 16436
rect 21499 16405 21511 16408
rect 21453 16399 21511 16405
rect 21542 16396 21548 16408
rect 21600 16396 21606 16448
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 9824 16204 10241 16232
rect 9824 16192 9830 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 10502 16192 10508 16244
rect 10560 16232 10566 16244
rect 11882 16232 11888 16244
rect 10560 16204 11888 16232
rect 10560 16192 10566 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12158 16192 12164 16244
rect 12216 16192 12222 16244
rect 12529 16235 12587 16241
rect 12529 16201 12541 16235
rect 12575 16232 12587 16235
rect 14366 16232 14372 16244
rect 12575 16204 14372 16232
rect 12575 16201 12587 16204
rect 12529 16195 12587 16201
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 14826 16232 14832 16244
rect 14599 16204 14832 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 15013 16235 15071 16241
rect 15013 16201 15025 16235
rect 15059 16232 15071 16235
rect 17402 16232 17408 16244
rect 15059 16204 17408 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 17402 16192 17408 16204
rect 17460 16232 17466 16244
rect 17460 16204 17724 16232
rect 17460 16192 17466 16204
rect 7466 16124 7472 16176
rect 7524 16124 7530 16176
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 10735 16136 12848 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 12618 16056 12624 16108
rect 12676 16056 12682 16108
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7834 16028 7840 16040
rect 6871 16000 7840 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7834 15988 7840 16000
rect 7892 16028 7898 16040
rect 9582 16028 9588 16040
rect 7892 16000 9588 16028
rect 7892 15988 7898 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 11882 16028 11888 16040
rect 10836 16000 11888 16028
rect 10836 15988 10842 16000
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12308 16000 12725 16028
rect 12308 15988 12314 16000
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 12820 15960 12848 16136
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 17221 16167 17279 16173
rect 13596 16136 13952 16164
rect 13596 16124 13602 16136
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13556 16068 13737 16096
rect 13357 15963 13415 15969
rect 13357 15960 13369 15963
rect 8220 15932 8984 15960
rect 12820 15932 13369 15960
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 8220 15892 8248 15932
rect 5224 15864 8248 15892
rect 5224 15852 5230 15864
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8570 15892 8576 15904
rect 8352 15864 8576 15892
rect 8352 15852 8358 15864
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 8956 15892 8984 15932
rect 13357 15929 13369 15932
rect 13403 15929 13415 15963
rect 13556 15960 13584 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 13924 16037 13952 16136
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 17586 16164 17592 16176
rect 17267 16136 17592 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 17586 16124 17592 16136
rect 17644 16124 17650 16176
rect 17696 16164 17724 16204
rect 17862 16192 17868 16244
rect 17920 16232 17926 16244
rect 20162 16232 20168 16244
rect 17920 16204 20168 16232
rect 17920 16192 17926 16204
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 21358 16232 21364 16244
rect 20272 16204 21364 16232
rect 20272 16164 20300 16204
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 22646 16192 22652 16244
rect 22704 16192 22710 16244
rect 23290 16192 23296 16244
rect 23348 16232 23354 16244
rect 23348 16204 25084 16232
rect 23348 16192 23354 16204
rect 21450 16164 21456 16176
rect 17696 16136 20300 16164
rect 21206 16136 21456 16164
rect 21450 16124 21456 16136
rect 21508 16164 21514 16176
rect 22664 16164 22692 16192
rect 21508 16136 22692 16164
rect 21508 16124 21514 16136
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15712 16068 15945 16096
rect 15712 16056 15718 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18322 16096 18328 16108
rect 18095 16068 18328 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19334 16096 19340 16108
rect 18739 16068 19340 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19484 16068 19717 16096
rect 19484 16056 19490 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 24397 16099 24455 16105
rect 19705 16059 19763 16065
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13688 16000 13829 16028
rect 13688 15988 13694 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 19981 16031 20039 16037
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 20070 16028 20076 16040
rect 20027 16000 20076 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 20070 15988 20076 16000
rect 20128 15988 20134 16040
rect 20346 15988 20352 16040
rect 20404 16028 20410 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 20404 16000 22017 16028
rect 20404 15988 20410 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22281 16031 22339 16037
rect 22281 16028 22293 16031
rect 22005 15991 22063 15997
rect 22112 16000 22293 16028
rect 18138 15960 18144 15972
rect 13556 15932 18144 15960
rect 13357 15923 13415 15929
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 11606 15892 11612 15904
rect 8956 15864 11612 15892
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 16356 15864 17325 15892
rect 16356 15852 16362 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 17313 15855 17371 15861
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17460 15864 17877 15892
rect 17460 15852 17466 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 18509 15895 18567 15901
rect 18509 15892 18521 15895
rect 18472 15864 18521 15892
rect 18472 15852 18478 15864
rect 18509 15861 18521 15864
rect 18555 15861 18567 15895
rect 18509 15855 18567 15861
rect 20530 15852 20536 15904
rect 20588 15892 20594 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 20588 15864 21465 15892
rect 20588 15852 20594 15864
rect 21453 15861 21465 15864
rect 21499 15892 21511 15895
rect 22112 15892 22140 16000
rect 22281 15997 22293 16000
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 23400 16028 23428 16082
rect 24397 16065 24409 16099
rect 24443 16096 24455 16099
rect 24670 16096 24676 16108
rect 24443 16068 24676 16096
rect 24443 16065 24455 16068
rect 24397 16059 24455 16065
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 25056 16105 25084 16204
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 23658 16028 23664 16040
rect 22704 16000 23664 16028
rect 22704 15988 22710 16000
rect 23658 15988 23664 16000
rect 23716 16028 23722 16040
rect 24762 16028 24768 16040
rect 23716 16000 24768 16028
rect 23716 15988 23722 16000
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 21499 15864 22140 15892
rect 21499 15861 21511 15864
rect 21453 15855 21511 15861
rect 22646 15852 22652 15904
rect 22704 15892 22710 15904
rect 23753 15895 23811 15901
rect 23753 15892 23765 15895
rect 22704 15864 23765 15892
rect 22704 15852 22710 15864
rect 23753 15861 23765 15864
rect 23799 15861 23811 15895
rect 23753 15855 23811 15861
rect 24026 15852 24032 15904
rect 24084 15892 24090 15904
rect 24857 15895 24915 15901
rect 24857 15892 24869 15895
rect 24084 15864 24869 15892
rect 24084 15852 24090 15864
rect 24857 15861 24869 15864
rect 24903 15861 24915 15895
rect 24857 15855 24915 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9122 15648 9128 15700
rect 9180 15648 9186 15700
rect 11698 15648 11704 15700
rect 11756 15648 11762 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 14182 15688 14188 15700
rect 12676 15660 14188 15688
rect 12676 15648 12682 15660
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 16564 15691 16622 15697
rect 16564 15657 16576 15691
rect 16610 15688 16622 15691
rect 18598 15688 18604 15700
rect 16610 15660 18604 15688
rect 16610 15657 16622 15660
rect 16564 15651 16622 15657
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 22060 15660 24808 15688
rect 22060 15648 22066 15660
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 13630 15620 13636 15632
rect 11388 15592 13636 15620
rect 11388 15580 11394 15592
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 17678 15580 17684 15632
rect 17736 15620 17742 15632
rect 17736 15592 17908 15620
rect 17736 15580 17742 15592
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9640 15524 9689 15552
rect 9640 15512 9646 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 12250 15512 12256 15564
rect 12308 15512 12314 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 15194 15552 15200 15564
rect 12860 15524 15200 15552
rect 12860 15512 12866 15524
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15552 16359 15555
rect 16574 15552 16580 15564
rect 16347 15524 16580 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16574 15512 16580 15524
rect 16632 15512 16638 15564
rect 14458 15444 14464 15496
rect 14516 15444 14522 15496
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 17644 15456 17710 15484
rect 17644 15444 17650 15456
rect 12069 15419 12127 15425
rect 12069 15385 12081 15419
rect 12115 15416 12127 15419
rect 12618 15416 12624 15428
rect 12115 15388 12624 15416
rect 12115 15385 12127 15388
rect 12069 15379 12127 15385
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 9490 15308 9496 15360
rect 9548 15308 9554 15360
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10594 15348 10600 15360
rect 10284 15320 10600 15348
rect 10284 15308 10290 15320
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 12161 15351 12219 15357
rect 12161 15317 12173 15351
rect 12207 15348 12219 15351
rect 12802 15348 12808 15360
rect 12207 15320 12808 15348
rect 12207 15317 12219 15320
rect 12161 15311 12219 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 17880 15348 17908 15592
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20254 15552 20260 15564
rect 19475 15524 20260 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20254 15512 20260 15524
rect 20312 15552 20318 15564
rect 22278 15552 22284 15564
rect 20312 15524 22284 15552
rect 20312 15512 20318 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 22646 15552 22652 15564
rect 22603 15524 22652 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 23290 15512 23296 15564
rect 23348 15552 23354 15564
rect 24029 15555 24087 15561
rect 24029 15552 24041 15555
rect 23348 15524 24041 15552
rect 23348 15512 23354 15524
rect 24029 15521 24041 15524
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 23658 15444 23664 15496
rect 23716 15444 23722 15496
rect 24780 15493 24808 15660
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 19702 15416 19708 15428
rect 19536 15388 19708 15416
rect 19536 15360 19564 15388
rect 19702 15376 19708 15388
rect 19760 15376 19766 15428
rect 21450 15416 21456 15428
rect 20930 15388 21456 15416
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 22554 15416 22560 15428
rect 22152 15388 22560 15416
rect 22152 15376 22158 15388
rect 22554 15376 22560 15388
rect 22612 15376 22618 15428
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 17552 15320 18061 15348
rect 17552 15308 17558 15320
rect 18049 15317 18061 15320
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 20128 15320 21189 15348
rect 20128 15308 20134 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 23474 15348 23480 15360
rect 21683 15320 23480 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 24578 15308 24584 15360
rect 24636 15308 24642 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 13722 15144 13728 15156
rect 13679 15116 13728 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14458 15144 14464 15156
rect 14047 15116 14464 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15896 15116 15945 15144
rect 15896 15104 15902 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 19978 15104 19984 15156
rect 20036 15104 20042 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20680 15116 21189 15144
rect 20680 15104 20686 15116
rect 21177 15113 21189 15116
rect 21223 15113 21235 15147
rect 21177 15107 21235 15113
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22244 15116 22293 15144
rect 22244 15104 22250 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22281 15107 22339 15113
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 23290 15144 23296 15156
rect 22612 15116 23296 15144
rect 22612 15104 22618 15116
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 7524 15048 8418 15076
rect 7524 15036 7530 15048
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 10505 15079 10563 15085
rect 10505 15045 10517 15079
rect 10551 15076 10563 15079
rect 11974 15076 11980 15088
rect 10551 15048 11980 15076
rect 10551 15045 10563 15048
rect 10505 15039 10563 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 18693 15079 18751 15085
rect 18693 15045 18705 15079
rect 18739 15076 18751 15079
rect 20162 15076 20168 15088
rect 18739 15048 20168 15076
rect 18739 15045 18751 15048
rect 18693 15039 18751 15045
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 9692 15008 9720 15036
rect 10597 15011 10655 15017
rect 9692 14980 9812 15008
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 6420 14912 7665 14940
rect 6420 14900 6426 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8294 14940 8300 14952
rect 7975 14912 8300 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 7668 14804 7696 14903
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9784 14940 9812 14980
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 11606 15008 11612 15020
rect 10643 14980 11612 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 19392 14980 19901 15008
rect 19392 14968 19398 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 21048 14980 21097 15008
rect 21048 14968 21054 14980
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 22060 14980 22477 15008
rect 22060 14968 22066 14980
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 22612 14980 23949 15008
rect 22612 14968 22618 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 9784 14912 10701 14940
rect 9677 14903 9735 14909
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 9030 14832 9036 14884
rect 9088 14872 9094 14884
rect 9692 14872 9720 14903
rect 14090 14900 14096 14952
rect 14148 14900 14154 14952
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 15746 14940 15752 14952
rect 14323 14912 15752 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 16022 14900 16028 14952
rect 16080 14900 16086 14952
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16482 14940 16488 14952
rect 16255 14912 16488 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 22646 14940 22652 14952
rect 21407 14912 22652 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 13630 14872 13636 14884
rect 9088 14844 13636 14872
rect 9088 14832 9094 14844
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 18874 14872 18880 14884
rect 15611 14844 18880 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 19521 14875 19579 14881
rect 19521 14841 19533 14875
rect 19567 14872 19579 14875
rect 21910 14872 21916 14884
rect 19567 14844 21916 14872
rect 19567 14841 19579 14844
rect 19521 14835 19579 14841
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 9950 14804 9956 14816
rect 7668 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 16390 14804 16396 14816
rect 12308 14776 16396 14804
rect 12308 14764 12314 14776
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 18785 14807 18843 14813
rect 18785 14804 18797 14807
rect 18748 14776 18797 14804
rect 18748 14764 18754 14776
rect 18785 14773 18797 14776
rect 18831 14773 18843 14807
rect 18785 14767 18843 14773
rect 20717 14807 20775 14813
rect 20717 14773 20729 14807
rect 20763 14804 20775 14807
rect 23566 14804 23572 14816
rect 20763 14776 23572 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7800 14572 8125 14600
rect 7800 14560 7806 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 19518 14600 19524 14612
rect 8113 14563 8171 14569
rect 13372 14572 19524 14600
rect 6362 14424 6368 14476
rect 6420 14424 6426 14476
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14464 6699 14467
rect 9306 14464 9312 14476
rect 6687 14436 9312 14464
rect 6687 14433 6699 14436
rect 6641 14427 6699 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11940 14436 11989 14464
rect 11940 14424 11946 14436
rect 11977 14433 11989 14436
rect 12023 14464 12035 14467
rect 12066 14464 12072 14476
rect 12023 14436 12072 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 13372 14405 13400 14572
rect 19518 14560 19524 14572
rect 19576 14600 19582 14612
rect 26694 14600 26700 14612
rect 19576 14572 26700 14600
rect 19576 14560 19582 14572
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 16482 14492 16488 14544
rect 16540 14532 16546 14544
rect 17862 14532 17868 14544
rect 16540 14504 17868 14532
rect 16540 14492 16546 14504
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 13630 14424 13636 14476
rect 13688 14464 13694 14476
rect 15378 14464 15384 14476
rect 13688 14436 15384 14464
rect 13688 14424 13694 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 15528 14436 16957 14464
rect 15528 14424 15534 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 22278 14424 22284 14476
rect 22336 14424 22342 14476
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 12575 14368 13369 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 16807 14368 17785 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 19668 14368 20453 14396
rect 19668 14356 19674 14368
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 23658 14356 23664 14408
rect 23716 14356 23722 14408
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 7374 14288 7380 14340
rect 7432 14288 7438 14340
rect 10229 14331 10287 14337
rect 10229 14297 10241 14331
rect 10275 14297 10287 14331
rect 10229 14291 10287 14297
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 10244 14260 10272 14291
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 13538 14328 13544 14340
rect 11532 14300 13544 14328
rect 11532 14260 11560 14300
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 20346 14328 20352 14340
rect 16546 14300 20352 14328
rect 9824 14232 11560 14260
rect 9824 14220 9830 14232
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12768 14232 13001 14260
rect 12768 14220 12774 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 12989 14223 13047 14229
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13449 14263 13507 14269
rect 13449 14260 13461 14263
rect 13320 14232 13461 14260
rect 13320 14220 13326 14232
rect 13449 14229 13461 14232
rect 13495 14260 13507 14263
rect 14918 14260 14924 14272
rect 13495 14232 14924 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 16393 14263 16451 14269
rect 16393 14229 16405 14263
rect 16439 14260 16451 14263
rect 16546 14260 16574 14300
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 22278 14288 22284 14340
rect 22336 14328 22342 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 22336 14300 22569 14328
rect 22336 14288 22342 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 22557 14291 22615 14297
rect 16439 14232 16574 14260
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16724 14232 16865 14260
rect 16724 14220 16730 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20036 14232 20269 14260
rect 20036 14220 20042 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23348 14232 24041 14260
rect 23348 14220 23354 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24029 14223 24087 14229
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 24176 14232 24593 14260
rect 24176 14220 24182 14232
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 7524 14028 8432 14056
rect 7524 14016 7530 14028
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 8021 13991 8079 13997
rect 8021 13988 8033 13991
rect 7800 13960 8033 13988
rect 7800 13948 7806 13960
rect 8021 13957 8033 13960
rect 8067 13957 8079 13991
rect 8404 13988 8432 14028
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 12989 14059 13047 14065
rect 8904 14028 12940 14056
rect 8904 14016 8910 14028
rect 8478 13988 8484 14000
rect 8404 13960 8484 13988
rect 8021 13951 8079 13957
rect 8478 13948 8484 13960
rect 8536 13948 8542 14000
rect 9766 13948 9772 14000
rect 9824 13948 9830 14000
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10965 13991 11023 13997
rect 10965 13988 10977 13991
rect 10008 13960 10977 13988
rect 10008 13948 10014 13960
rect 10965 13957 10977 13960
rect 11011 13957 11023 13991
rect 12912 13988 12940 14028
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 18601 14059 18659 14065
rect 13035 14028 18460 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13262 13988 13268 14000
rect 12912 13960 13268 13988
rect 10965 13951 11023 13957
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 17586 13988 17592 14000
rect 16868 13960 17592 13988
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 11882 13920 11888 13932
rect 10275 13892 11888 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10980 13864 11008 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 16114 13920 16120 13932
rect 15252 13892 16120 13920
rect 15252 13880 15258 13892
rect 16114 13880 16120 13892
rect 16172 13920 16178 13932
rect 16868 13920 16896 13960
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 18432 13988 18460 14028
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18966 14056 18972 14068
rect 18647 14028 18972 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 24762 14056 24768 14068
rect 20211 14028 24768 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 19242 13988 19248 14000
rect 18432 13960 19248 13988
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 19521 13991 19579 13997
rect 19521 13957 19533 13991
rect 19567 13988 19579 13991
rect 21634 13988 21640 14000
rect 19567 13960 21640 13988
rect 19567 13957 19579 13960
rect 19521 13951 19579 13957
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 24578 13988 24584 14000
rect 22296 13960 24584 13988
rect 16172 13892 16896 13920
rect 16172 13880 16178 13892
rect 20346 13880 20352 13932
rect 20404 13880 20410 13932
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 22296 13929 22324 13960
rect 24578 13948 24584 13960
rect 24636 13948 24642 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20864 13892 21097 13920
rect 20864 13880 20870 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 24118 13880 24124 13932
rect 24176 13880 24182 13932
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7340 13824 7757 13852
rect 7340 13812 7346 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8536 13824 9628 13852
rect 8536 13812 8542 13824
rect 9600 13784 9628 13824
rect 10962 13812 10968 13864
rect 11020 13812 11026 13864
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12584 13824 13093 13852
rect 12584 13812 12590 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 11238 13784 11244 13796
rect 9600 13756 11244 13784
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 13280 13784 13308 13815
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 15528 13824 15577 13852
rect 15528 13812 15534 13824
rect 15565 13821 15577 13824
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 19058 13852 19064 13864
rect 17644 13824 19064 13852
rect 17644 13812 17650 13824
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 19702 13812 19708 13864
rect 19760 13812 19766 13864
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13852 23351 13855
rect 24854 13852 24860 13864
rect 23339 13824 24860 13852
rect 23339 13821 23351 13824
rect 23293 13815 23351 13821
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 20901 13787 20959 13793
rect 11572 13756 13216 13784
rect 13280 13756 13952 13784
rect 11572 13744 11578 13756
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11112 13688 11897 13716
rect 11112 13676 11118 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 11885 13679 11943 13685
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12492 13688 12633 13716
rect 12492 13676 12498 13688
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 13188 13716 13216 13756
rect 13924 13728 13952 13756
rect 18156 13756 20300 13784
rect 13630 13716 13636 13728
rect 13188 13688 13636 13716
rect 12621 13679 12679 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13906 13676 13912 13728
rect 13964 13676 13970 13728
rect 14080 13719 14138 13725
rect 14080 13685 14092 13719
rect 14126 13716 14138 13719
rect 14274 13716 14280 13728
rect 14126 13688 14280 13716
rect 14126 13685 14138 13688
rect 14080 13679 14138 13685
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 18156 13716 18184 13756
rect 17368 13688 18184 13716
rect 17368 13676 17374 13688
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 20162 13716 20168 13728
rect 18380 13688 20168 13716
rect 18380 13676 18386 13688
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 20272 13716 20300 13756
rect 20901 13753 20913 13787
rect 20947 13784 20959 13787
rect 21818 13784 21824 13796
rect 20947 13756 21824 13784
rect 20947 13753 20959 13756
rect 20901 13747 20959 13753
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 21082 13716 21088 13728
rect 20272 13688 21088 13716
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 7892 13484 8217 13512
rect 7892 13472 7898 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8205 13475 8263 13481
rect 9214 13472 9220 13524
rect 9272 13472 9278 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 9364 13484 9996 13512
rect 9364 13472 9370 13484
rect 9858 13444 9864 13456
rect 9692 13416 9864 13444
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6420 13348 6469 13376
rect 6420 13336 6426 13348
rect 6457 13345 6469 13348
rect 6503 13376 6515 13379
rect 7282 13376 7288 13388
rect 6503 13348 7288 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 9692 13385 9720 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9968 13376 9996 13484
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 11204 13484 13001 13512
rect 11204 13472 11210 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14918 13512 14924 13524
rect 13964 13484 14924 13512
rect 13964 13472 13970 13484
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15528 13484 19334 13512
rect 15528 13472 15534 13484
rect 13814 13444 13820 13456
rect 11716 13416 13820 13444
rect 9815 13348 9996 13376
rect 10413 13379 10471 13385
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 11716 13376 11744 13416
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 15654 13444 15660 13456
rect 15304 13416 15660 13444
rect 10459 13348 11744 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 10428 13308 10456 13339
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 12124 13348 13553 13376
rect 12124 13336 12130 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 15304 13376 15332 13416
rect 15654 13404 15660 13416
rect 15712 13444 15718 13456
rect 16206 13444 16212 13456
rect 15712 13416 16212 13444
rect 15712 13404 15718 13416
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 19306 13444 19334 13484
rect 19886 13444 19892 13456
rect 19306 13416 19892 13444
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 26050 13444 26056 13456
rect 20220 13416 26056 13444
rect 20220 13404 20226 13416
rect 26050 13404 26056 13416
rect 26108 13404 26114 13456
rect 13688 13348 15332 13376
rect 13688 13336 13694 13348
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15746 13376 15752 13388
rect 15436 13348 15752 13376
rect 15436 13336 15442 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 21269 13379 21327 13385
rect 17696 13348 21220 13376
rect 13446 13308 13452 13320
rect 9180 13280 10456 13308
rect 12084 13280 13452 13308
rect 9180 13268 9186 13280
rect 6733 13243 6791 13249
rect 6733 13209 6745 13243
rect 6779 13240 6791 13243
rect 6779 13212 6914 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 6886 13172 6914 13212
rect 7466 13200 7472 13252
rect 7524 13200 7530 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 10594 13240 10600 13252
rect 9631 13212 10600 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 10689 13243 10747 13249
rect 10689 13209 10701 13243
rect 10735 13209 10747 13243
rect 10689 13203 10747 13209
rect 9766 13172 9772 13184
rect 6886 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 10704 13172 10732 13203
rect 11238 13200 11244 13252
rect 11296 13200 11302 13252
rect 12084 13172 12112 13280
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 15565 13311 15623 13317
rect 14516 13280 15516 13308
rect 14516 13268 14522 13280
rect 13357 13243 13415 13249
rect 13357 13209 13369 13243
rect 13403 13240 13415 13243
rect 14550 13240 14556 13252
rect 13403 13212 14556 13240
rect 13403 13209 13415 13212
rect 13357 13203 13415 13209
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 15488 13240 15516 13280
rect 15565 13277 15577 13311
rect 15611 13308 15623 13311
rect 17310 13308 17316 13320
rect 15611 13280 17316 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 17696 13240 17724 13348
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 21192 13317 21220 13348
rect 21269 13345 21281 13379
rect 21315 13376 21327 13379
rect 21358 13376 21364 13388
rect 21315 13348 21364 13376
rect 21315 13345 21327 13348
rect 21269 13339 21327 13345
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 21453 13379 21511 13385
rect 21453 13345 21465 13379
rect 21499 13376 21511 13379
rect 23382 13376 23388 13388
rect 21499 13348 23388 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 23532 13348 24808 13376
rect 23532 13336 23538 13348
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 17828 13280 19441 13308
rect 17828 13268 17834 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 21177 13311 21235 13317
rect 21177 13277 21189 13311
rect 21223 13277 21235 13311
rect 21177 13271 21235 13277
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 24026 13308 24032 13320
rect 22879 13280 24032 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 15488 13212 17724 13240
rect 17862 13200 17868 13252
rect 17920 13200 17926 13252
rect 18049 13243 18107 13249
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18506 13240 18512 13252
rect 18095 13212 18512 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18598 13200 18604 13252
rect 18656 13200 18662 13252
rect 20254 13200 20260 13252
rect 20312 13200 20318 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 22204 13240 22232 13271
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24780 13317 24808 13348
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 20404 13212 22232 13240
rect 23845 13243 23903 13249
rect 20404 13200 20410 13212
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 24946 13240 24952 13252
rect 23891 13212 24952 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 10704 13144 12112 13172
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 13630 13172 13636 13184
rect 13495 13144 13636 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14642 13172 14648 13184
rect 14056 13144 14648 13172
rect 14056 13132 14062 13144
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 15654 13132 15660 13184
rect 15712 13132 15718 13184
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 16632 13144 18705 13172
rect 16632 13132 16638 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13172 20867 13175
rect 21174 13172 21180 13184
rect 20855 13144 21180 13172
rect 20855 13141 20867 13144
rect 20809 13135 20867 13141
rect 21174 13132 21180 13144
rect 21232 13132 21238 13184
rect 24578 13132 24584 13184
rect 24636 13132 24642 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6687 12940 7512 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 6972 12872 7236 12900
rect 6972 12860 6978 12872
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 7208 12773 7236 12872
rect 7484 12832 7512 12940
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7616 12940 7849 12968
rect 7616 12928 7622 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 7837 12931 7895 12937
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9582 12968 9588 12980
rect 9079 12940 9588 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11054 12968 11060 12980
rect 10827 12940 11060 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 8205 12903 8263 12909
rect 8205 12869 8217 12903
rect 8251 12900 8263 12903
rect 8294 12900 8300 12912
rect 8251 12872 8300 12900
rect 8251 12869 8263 12872
rect 8205 12863 8263 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 9490 12860 9496 12912
rect 9548 12900 9554 12912
rect 10428 12900 10456 12931
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 13725 12971 13783 12977
rect 11808 12940 12572 12968
rect 9548 12872 10456 12900
rect 10873 12903 10931 12909
rect 9548 12860 9554 12872
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 11808 12900 11836 12940
rect 10919 12872 11836 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 11882 12860 11888 12912
rect 11940 12860 11946 12912
rect 7484 12804 8524 12832
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 4212 12736 7113 12764
rect 4212 12724 4218 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7193 12727 7251 12733
rect 7392 12736 8309 12764
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 7392 12696 7420 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8386 12724 8392 12776
rect 8444 12724 8450 12776
rect 4304 12668 7420 12696
rect 8496 12696 8524 12804
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 12434 12832 12440 12844
rect 9508 12804 12440 12832
rect 9508 12773 9536 12804
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9766 12764 9772 12776
rect 9723 12736 9772 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 10962 12764 10968 12776
rect 9824 12736 10968 12764
rect 9824 12724 9830 12736
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 12544 12764 12572 12940
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 15010 12968 15016 12980
rect 13771 12940 15016 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15289 12971 15347 12977
rect 15289 12937 15301 12971
rect 15335 12968 15347 12971
rect 15335 12940 15516 12968
rect 15335 12937 15347 12940
rect 15289 12931 15347 12937
rect 12713 12903 12771 12909
rect 12713 12869 12725 12903
rect 12759 12900 12771 12903
rect 13814 12900 13820 12912
rect 12759 12872 13820 12900
rect 12759 12869 12771 12872
rect 12713 12863 12771 12869
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 13906 12860 13912 12912
rect 13964 12900 13970 12912
rect 13964 12872 14780 12900
rect 13964 12860 13970 12872
rect 13722 12792 13728 12844
rect 13780 12832 13786 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13780 12804 14105 12832
rect 13780 12792 13786 12804
rect 14093 12801 14105 12804
rect 14139 12801 14151 12835
rect 14752 12832 14780 12872
rect 15102 12860 15108 12912
rect 15160 12900 15166 12912
rect 15381 12903 15439 12909
rect 15381 12900 15393 12903
rect 15160 12872 15393 12900
rect 15160 12860 15166 12872
rect 15381 12869 15393 12872
rect 15427 12869 15439 12903
rect 15488 12900 15516 12940
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 16666 12968 16672 12980
rect 15712 12940 16672 12968
rect 15712 12928 15718 12940
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 16816 12940 17325 12968
rect 16816 12928 16822 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18693 12971 18751 12977
rect 18095 12940 18644 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18322 12900 18328 12912
rect 15488 12872 18328 12900
rect 15381 12863 15439 12869
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 14752 12804 17233 12832
rect 14093 12795 14151 12801
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17460 12804 18245 12832
rect 17460 12792 17466 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18616 12832 18644 12940
rect 18693 12937 18705 12971
rect 18739 12937 18751 12971
rect 18693 12931 18751 12937
rect 19061 12971 19119 12977
rect 19061 12937 19073 12971
rect 19107 12968 19119 12971
rect 20346 12968 20352 12980
rect 19107 12940 20352 12968
rect 19107 12937 19119 12940
rect 19061 12931 19119 12937
rect 18708 12900 18736 12931
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 21177 12971 21235 12977
rect 21177 12937 21189 12971
rect 21223 12968 21235 12971
rect 21266 12968 21272 12980
rect 21223 12940 21272 12968
rect 21223 12937 21235 12940
rect 21177 12931 21235 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 22554 12968 22560 12980
rect 22051 12940 22560 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 20990 12900 20996 12912
rect 18708 12872 20996 12900
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 23290 12900 23296 12912
rect 21376 12872 23296 12900
rect 18616 12804 19288 12832
rect 18233 12795 18291 12801
rect 13814 12764 13820 12776
rect 11756 12736 12480 12764
rect 12544 12736 13820 12764
rect 11756 12724 11762 12736
rect 10318 12696 10324 12708
rect 8496 12668 10324 12696
rect 4304 12656 4310 12668
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 12342 12696 12348 12708
rect 10652 12668 12348 12696
rect 10652 12656 10658 12668
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 12452 12696 12480 12736
rect 13814 12724 13820 12736
rect 13872 12764 13878 12776
rect 13998 12764 14004 12776
rect 13872 12736 14004 12764
rect 13872 12724 13878 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12733 14243 12767
rect 14185 12727 14243 12733
rect 13906 12696 13912 12708
rect 12452 12668 13912 12696
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 14200 12696 14228 12727
rect 14274 12724 14280 12776
rect 14332 12724 14338 12776
rect 14918 12724 14924 12776
rect 14976 12764 14982 12776
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 14976 12736 15485 12764
rect 14976 12724 14982 12736
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 17497 12767 17555 12773
rect 16080 12736 17264 12764
rect 16080 12724 16086 12736
rect 16758 12696 16764 12708
rect 14200 12668 15332 12696
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 14921 12631 14979 12637
rect 14921 12628 14933 12631
rect 12492 12600 14933 12628
rect 12492 12588 12498 12600
rect 14921 12597 14933 12600
rect 14967 12597 14979 12631
rect 15304 12628 15332 12668
rect 16546 12668 16764 12696
rect 16546 12628 16574 12668
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 17236 12696 17264 12736
rect 17497 12733 17509 12767
rect 17543 12764 17555 12767
rect 18966 12764 18972 12776
rect 17543 12736 18972 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 19153 12767 19211 12773
rect 19153 12733 19165 12767
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19168 12696 19196 12727
rect 17236 12668 19196 12696
rect 15304 12600 16574 12628
rect 16853 12631 16911 12637
rect 14921 12591 14979 12597
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 18874 12628 18880 12640
rect 16899 12600 18880 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19260 12628 19288 12804
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19852 12804 20085 12832
rect 19852 12792 19858 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20772 12804 21097 12832
rect 20772 12792 20778 12804
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 20530 12764 20536 12776
rect 19383 12736 20536 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 21376 12773 21404 12872
rect 23290 12860 23296 12872
rect 23348 12860 23354 12912
rect 23750 12860 23756 12912
rect 23808 12860 23814 12912
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 22830 12724 22836 12776
rect 22888 12764 22894 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22888 12736 23029 12764
rect 22888 12724 22894 12736
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 24670 12764 24676 12776
rect 23017 12727 23075 12733
rect 23124 12736 24676 12764
rect 19886 12656 19892 12708
rect 19944 12656 19950 12708
rect 20717 12699 20775 12705
rect 20717 12665 20729 12699
rect 20763 12696 20775 12699
rect 23124 12696 23152 12736
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 20763 12668 23152 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 22094 12628 22100 12640
rect 19260 12600 22100 12628
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 23382 12588 23388 12640
rect 23440 12628 23446 12640
rect 24765 12631 24823 12637
rect 24765 12628 24777 12631
rect 23440 12600 24777 12628
rect 23440 12588 23446 12600
rect 24765 12597 24777 12600
rect 24811 12597 24823 12631
rect 24765 12591 24823 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7064 12396 7573 12424
rect 7064 12384 7070 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 7561 12387 7619 12393
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 8352 12396 8401 12424
rect 8352 12384 8358 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 8389 12387 8447 12393
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10100 12396 10241 12424
rect 10100 12384 10106 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12618 12384 12624 12436
rect 12676 12384 12682 12436
rect 14366 12384 14372 12436
rect 14424 12384 14430 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 18598 12424 18604 12436
rect 14884 12396 18604 12424
rect 14884 12384 14890 12396
rect 18598 12384 18604 12396
rect 18656 12424 18662 12436
rect 20990 12424 20996 12436
rect 18656 12396 20996 12424
rect 18656 12384 18662 12396
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10502 12356 10508 12368
rect 10192 12328 10508 12356
rect 10192 12316 10198 12328
rect 10502 12316 10508 12328
rect 10560 12316 10566 12368
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 12526 12356 12532 12368
rect 11848 12328 12532 12356
rect 11848 12316 11854 12328
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 15102 12356 15108 12368
rect 14608 12328 15108 12356
rect 14608 12316 14614 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 17034 12356 17040 12368
rect 16724 12328 17040 12356
rect 16724 12316 16730 12328
rect 17034 12316 17040 12328
rect 17092 12356 17098 12368
rect 17218 12356 17224 12368
rect 17092 12328 17224 12356
rect 17092 12316 17098 12328
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17678 12356 17684 12368
rect 17368 12328 17684 12356
rect 17368 12316 17374 12328
rect 17678 12316 17684 12328
rect 17736 12316 17742 12368
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 9272 12260 10793 12288
rect 9272 12248 9278 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13354 12288 13360 12300
rect 13311 12260 13360 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13354 12248 13360 12260
rect 13412 12288 13418 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 13412 12260 14933 12288
rect 13412 12248 13418 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 19150 12288 19156 12300
rect 14921 12251 14979 12257
rect 17144 12260 19156 12288
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 17034 12220 17040 12232
rect 13035 12192 17040 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 17034 12180 17040 12192
rect 17092 12220 17098 12232
rect 17144 12220 17172 12260
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20312 12260 20361 12288
rect 20312 12248 20318 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 24578 12288 24584 12300
rect 20349 12251 20407 12257
rect 22848 12260 24584 12288
rect 17092 12192 17172 12220
rect 17221 12223 17279 12229
rect 17092 12180 17098 12192
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17770 12220 17776 12232
rect 17267 12192 17776 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 19242 12220 19248 12232
rect 18739 12192 19248 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19518 12180 19524 12232
rect 19576 12180 19582 12232
rect 22094 12180 22100 12232
rect 22152 12220 22158 12232
rect 22278 12220 22284 12232
rect 22152 12192 22284 12220
rect 22152 12180 22158 12192
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22848 12229 22876 12260
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 23624 12192 24777 12220
rect 23624 12180 23630 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 12526 12152 12532 12164
rect 11839 12124 12532 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 12952 12124 13093 12152
rect 12952 12112 12958 12124
rect 13081 12121 13093 12124
rect 13127 12152 13139 12155
rect 13722 12152 13728 12164
rect 13127 12124 13728 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 14458 12112 14464 12164
rect 14516 12152 14522 12164
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14516 12124 14841 12152
rect 14516 12112 14522 12124
rect 14829 12121 14841 12124
rect 14875 12121 14887 12155
rect 14829 12115 14887 12121
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 17957 12155 18015 12161
rect 17957 12152 17969 12155
rect 16908 12124 17969 12152
rect 16908 12112 16914 12124
rect 17957 12121 17969 12124
rect 18003 12121 18015 12155
rect 17957 12115 18015 12121
rect 18877 12155 18935 12161
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 19150 12152 19156 12164
rect 18923 12124 19156 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 20625 12155 20683 12161
rect 20625 12121 20637 12155
rect 20671 12152 20683 12155
rect 20714 12152 20720 12164
rect 20671 12124 20720 12152
rect 20671 12121 20683 12124
rect 20625 12115 20683 12121
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 23658 12152 23664 12164
rect 21850 12124 23664 12152
rect 23658 12112 23664 12124
rect 23716 12112 23722 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12618 12084 12624 12096
rect 11931 12056 12624 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 14700 12056 14749 12084
rect 14700 12044 14706 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 17494 12084 17500 12096
rect 15068 12056 17500 12084
rect 15068 12044 15074 12056
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 18564 12056 19625 12084
rect 18564 12044 18570 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 19702 12044 19708 12096
rect 19760 12084 19766 12096
rect 22097 12087 22155 12093
rect 22097 12084 22109 12087
rect 19760 12056 22109 12084
rect 19760 12044 19766 12056
rect 22097 12053 22109 12056
rect 22143 12053 22155 12087
rect 22097 12047 22155 12053
rect 23474 12044 23480 12096
rect 23532 12084 23538 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 23532 12056 24593 12084
rect 23532 12044 23538 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 9033 11883 9091 11889
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 9214 11880 9220 11892
rect 9079 11852 9220 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 9858 11880 9864 11892
rect 9815 11852 9864 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12345 11883 12403 11889
rect 12345 11849 12357 11883
rect 12391 11880 12403 11883
rect 12434 11880 12440 11892
rect 12391 11852 12440 11880
rect 12391 11849 12403 11852
rect 12345 11843 12403 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 13173 11883 13231 11889
rect 13173 11880 13185 11883
rect 12860 11852 13185 11880
rect 12860 11840 12866 11852
rect 13173 11849 13185 11852
rect 13219 11849 13231 11883
rect 13173 11843 13231 11849
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13320 11852 13645 11880
rect 13320 11840 13326 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14240 11852 14381 11880
rect 14240 11840 14246 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 14826 11880 14832 11892
rect 14783 11852 14832 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 16666 11880 16672 11892
rect 15212 11852 16672 11880
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 12710 11812 12716 11824
rect 10275 11784 12716 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 13354 11772 13360 11824
rect 13412 11812 13418 11824
rect 13722 11812 13728 11824
rect 13412 11784 13728 11812
rect 13412 11772 13418 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 15212 11812 15240 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 17000 11852 17325 11880
rect 17000 11840 17006 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 19334 11880 19340 11892
rect 18095 11852 19340 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 20622 11880 20628 11892
rect 19659 11852 20628 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 22186 11880 22192 11892
rect 20732 11852 22192 11880
rect 13832 11784 15240 11812
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9858 11744 9864 11756
rect 8628 11716 9864 11744
rect 8628 11704 8634 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10134 11704 10140 11756
rect 10192 11704 10198 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 13541 11747 13599 11753
rect 12483 11716 13492 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 7607 11648 10333 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 10321 11645 10333 11648
rect 10367 11676 10379 11679
rect 11054 11676 11060 11688
rect 10367 11648 11060 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 12066 11608 12072 11620
rect 11020 11580 12072 11608
rect 11020 11568 11026 11580
rect 12066 11568 12072 11580
rect 12124 11608 12130 11620
rect 12544 11608 12572 11639
rect 13262 11608 13268 11620
rect 12124 11580 12572 11608
rect 12728 11580 13268 11608
rect 12124 11568 12130 11580
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12728 11540 12756 11580
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 13464 11608 13492 11716
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 13832 11744 13860 11784
rect 15286 11772 15292 11824
rect 15344 11812 15350 11824
rect 15344 11784 17356 11812
rect 15344 11772 15350 11784
rect 13587 11716 13860 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 14148 11716 14872 11744
rect 14148 11704 14154 11716
rect 14844 11688 14872 11716
rect 15120 11716 17233 11744
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 13780 11648 14780 11676
rect 13780 11636 13786 11648
rect 14550 11608 14556 11620
rect 13464 11580 14556 11608
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 14752 11608 14780 11648
rect 14826 11636 14832 11688
rect 14884 11636 14890 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 14936 11608 14964 11639
rect 14752 11580 14964 11608
rect 12492 11512 12756 11540
rect 12492 11500 12498 11512
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13446 11540 13452 11552
rect 12860 11512 13452 11540
rect 12860 11500 12866 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 15120 11540 15148 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17328 11744 17356 11784
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 20732 11812 20760 11852
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 17460 11784 20760 11812
rect 20901 11815 20959 11821
rect 17460 11772 17466 11784
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 21082 11812 21088 11824
rect 20947 11784 21088 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 22370 11772 22376 11824
rect 22428 11772 22434 11824
rect 23382 11772 23388 11824
rect 23440 11772 23446 11824
rect 23658 11772 23664 11824
rect 23716 11812 23722 11824
rect 23716 11784 23874 11812
rect 23716 11772 23722 11784
rect 18417 11747 18475 11753
rect 17328 11716 17540 11744
rect 17221 11707 17279 11713
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16356 11648 17417 11676
rect 16356 11636 16362 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17512 11676 17540 11716
rect 18417 11713 18429 11747
rect 18463 11744 18475 11747
rect 19610 11744 19616 11756
rect 18463 11716 19616 11744
rect 18463 11713 18475 11716
rect 18417 11707 18475 11713
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11744 20039 11747
rect 21634 11744 21640 11756
rect 20027 11716 21640 11744
rect 20027 11713 20039 11716
rect 19981 11707 20039 11713
rect 21634 11704 21640 11716
rect 21692 11704 21698 11756
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22278 11704 22284 11756
rect 22336 11744 22342 11756
rect 22830 11744 22836 11756
rect 22336 11716 22836 11744
rect 22336 11704 22342 11716
rect 22830 11704 22836 11716
rect 22888 11744 22894 11756
rect 23109 11747 23167 11753
rect 23109 11744 23121 11747
rect 22888 11716 23121 11744
rect 22888 11704 22894 11716
rect 23109 11713 23121 11716
rect 23155 11713 23167 11747
rect 23109 11707 23167 11713
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17512 11648 18521 11676
rect 17405 11639 17463 11645
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19426 11676 19432 11688
rect 18739 11648 19432 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19628 11648 20085 11676
rect 16853 11611 16911 11617
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 19518 11608 19524 11620
rect 16899 11580 19524 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 13780 11512 15148 11540
rect 13780 11500 13786 11512
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 19628 11540 19656 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 20303 11648 21128 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 17828 11512 19656 11540
rect 17828 11500 17834 11512
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 19852 11512 21005 11540
rect 19852 11500 19858 11512
rect 20993 11509 21005 11512
rect 21039 11509 21051 11543
rect 21100 11540 21128 11648
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 22646 11608 22652 11620
rect 21600 11580 22652 11608
rect 21600 11568 21606 11580
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 22094 11540 22100 11552
rect 21100 11512 22100 11540
rect 20993 11503 21051 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 24854 11500 24860 11552
rect 24912 11500 24918 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 10652 11308 12633 11336
rect 10652 11296 10658 11308
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 12621 11299 12679 11305
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13722 11336 13728 11348
rect 13044 11308 13728 11336
rect 13044 11296 13050 11308
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 15194 11336 15200 11348
rect 14108 11308 15200 11336
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 9447 11172 11989 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 11977 11169 11989 11172
rect 12023 11200 12035 11203
rect 12158 11200 12164 11212
rect 12023 11172 12164 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12406 11172 13277 11200
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 12406 11132 12434 11172
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13538 11200 13544 11212
rect 13311 11172 13544 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 11112 11104 12434 11132
rect 12989 11135 13047 11141
rect 11112 11092 11118 11104
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 14108 11132 14136 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 17402 11336 17408 11348
rect 17267 11308 17408 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 19610 11296 19616 11348
rect 19668 11296 19674 11348
rect 21634 11296 21640 11348
rect 21692 11296 21698 11348
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 22370 11336 22376 11348
rect 22143 11308 22376 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 24581 11339 24639 11345
rect 24581 11336 24593 11339
rect 23348 11308 24593 11336
rect 23348 11296 23354 11308
rect 24581 11305 24593 11308
rect 24627 11305 24639 11339
rect 24581 11299 24639 11305
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 16485 11271 16543 11277
rect 16485 11268 16497 11271
rect 16356 11240 16497 11268
rect 16356 11228 16362 11240
rect 16485 11237 16497 11240
rect 16531 11237 16543 11271
rect 16485 11231 16543 11237
rect 17865 11271 17923 11277
rect 17865 11237 17877 11271
rect 17911 11268 17923 11271
rect 20809 11271 20867 11277
rect 17911 11240 20760 11268
rect 17911 11237 17923 11240
rect 17865 11231 17923 11237
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11200 14795 11203
rect 16850 11200 16856 11212
rect 14783 11172 16856 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 18322 11160 18328 11212
rect 18380 11160 18386 11212
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 19610 11200 19616 11212
rect 18555 11172 19616 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 20732 11200 20760 11240
rect 20809 11237 20821 11271
rect 20855 11268 20867 11271
rect 23842 11268 23848 11280
rect 20855 11240 23848 11268
rect 20855 11237 20867 11240
rect 20809 11231 20867 11237
rect 23842 11228 23848 11240
rect 23900 11228 23906 11280
rect 21174 11200 21180 11212
rect 20732 11172 21180 11200
rect 21174 11160 21180 11172
rect 21232 11160 21238 11212
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 23569 11203 23627 11209
rect 23569 11200 23581 11203
rect 21324 11172 23581 11200
rect 21324 11160 21330 11172
rect 23569 11169 23581 11172
rect 23615 11169 23627 11203
rect 23569 11163 23627 11169
rect 13035 11104 14136 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16172 11104 16896 11132
rect 16172 11092 16178 11104
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12802 11064 12808 11076
rect 11931 11036 12808 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 13127 11036 14964 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10870 10996 10876 11008
rect 9732 10968 10876 10996
rect 9732 10956 9738 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11422 10956 11428 11008
rect 11480 10956 11486 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 13722 10996 13728 11008
rect 12676 10968 13728 10996
rect 12676 10956 12682 10968
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 14936 10996 14964 11036
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 16868 11064 16896 11104
rect 17402 11092 17408 11144
rect 17460 11092 17466 11144
rect 18598 11132 18604 11144
rect 17512 11104 18604 11132
rect 17512 11064 17540 11104
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 20162 11092 20168 11144
rect 20220 11092 20226 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20272 11104 21005 11132
rect 16868 11036 17540 11064
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 18233 11067 18291 11073
rect 18233 11064 18245 11067
rect 18012 11036 18245 11064
rect 18012 11024 18018 11036
rect 18233 11033 18245 11036
rect 18279 11033 18291 11067
rect 18233 11027 18291 11033
rect 18432 11036 19104 11064
rect 15194 10996 15200 11008
rect 14936 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15654 10956 15660 11008
rect 15712 10996 15718 11008
rect 18432 10996 18460 11036
rect 15712 10968 18460 10996
rect 19076 10996 19104 11036
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 20272 11064 20300 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 22281 11135 22339 11141
rect 22281 11101 22293 11135
rect 22327 11132 22339 11135
rect 22738 11132 22744 11144
rect 22327 11104 22744 11132
rect 22327 11101 22339 11104
rect 22281 11095 22339 11101
rect 22738 11092 22744 11104
rect 22796 11092 22802 11144
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 19576 11036 20300 11064
rect 20349 11067 20407 11073
rect 19576 11024 19582 11036
rect 20349 11033 20361 11067
rect 20395 11064 20407 11067
rect 20438 11064 20444 11076
rect 20395 11036 20444 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 22940 11064 22968 11095
rect 24670 11092 24676 11144
rect 24728 11132 24734 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24728 11104 24777 11132
rect 24728 11092 24734 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 21968 11036 22968 11064
rect 21968 11024 21974 11036
rect 22002 10996 22008 11008
rect 19076 10968 22008 10996
rect 15712 10956 15718 10968
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22738 10956 22744 11008
rect 22796 10956 22802 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9824 10764 9965 10792
rect 9824 10752 9830 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 13722 10752 13728 10804
rect 13780 10752 13786 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15160 10764 15577 10792
rect 15160 10752 15166 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 17678 10792 17684 10804
rect 15565 10755 15623 10761
rect 15856 10764 17684 10792
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 7156 10696 8493 10724
rect 7156 10684 7162 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 9858 10724 9864 10736
rect 9706 10696 9864 10724
rect 8481 10687 8539 10693
rect 9858 10684 9864 10696
rect 9916 10724 9922 10736
rect 10594 10724 10600 10736
rect 9916 10696 10600 10724
rect 9916 10684 9922 10696
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 12406 10696 13001 10724
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 8202 10588 8208 10600
rect 7340 10560 8208 10588
rect 7340 10548 7346 10560
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 12406 10588 12434 10696
rect 12989 10693 13001 10696
rect 13035 10724 13047 10727
rect 13998 10724 14004 10736
rect 13035 10696 14004 10724
rect 13035 10693 13047 10696
rect 12989 10687 13047 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 14093 10727 14151 10733
rect 14093 10693 14105 10727
rect 14139 10724 14151 10727
rect 15856 10724 15884 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 24026 10792 24032 10804
rect 18708 10764 24032 10792
rect 14139 10696 15884 10724
rect 14139 10693 14151 10696
rect 14093 10687 14151 10693
rect 15930 10684 15936 10736
rect 15988 10684 15994 10736
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 15562 10656 15568 10668
rect 12943 10628 15568 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 18708 10665 18736 10764
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 19610 10684 19616 10736
rect 19668 10724 19674 10736
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 19668 10696 19993 10724
rect 19668 10684 19674 10696
rect 19981 10693 19993 10696
rect 20027 10693 20039 10727
rect 19981 10687 20039 10693
rect 21358 10684 21364 10736
rect 21416 10724 21422 10736
rect 23201 10727 23259 10733
rect 23201 10724 23213 10727
rect 21416 10696 23213 10724
rect 21416 10684 21422 10696
rect 23201 10693 23213 10696
rect 23247 10693 23259 10727
rect 23201 10687 23259 10693
rect 17497 10659 17555 10665
rect 15764 10628 17448 10656
rect 8996 10560 12434 10588
rect 13173 10591 13231 10597
rect 8996 10548 9002 10560
rect 13173 10557 13185 10591
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13188 10520 13216 10551
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13964 10560 14197 10588
rect 13964 10548 13970 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 13446 10520 13452 10532
rect 13188 10492 13452 10520
rect 13446 10480 13452 10492
rect 13504 10520 13510 10532
rect 14384 10520 14412 10551
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 15764 10588 15792 10628
rect 14884 10560 15792 10588
rect 14884 10548 14890 10560
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15896 10560 16037 10588
rect 15896 10548 15902 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 17310 10588 17316 10600
rect 16224 10560 17316 10588
rect 16132 10520 16160 10548
rect 13504 10492 16160 10520
rect 13504 10480 13510 10492
rect 11146 10412 11152 10464
rect 11204 10412 11210 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 12032 10424 12081 10452
rect 12032 10412 12038 10424
rect 12069 10421 12081 10424
rect 12115 10421 12127 10455
rect 12069 10415 12127 10421
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 16224 10452 16252 10560
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17420 10588 17448 10628
rect 17497 10625 17509 10659
rect 17543 10656 17555 10659
rect 18693 10659 18751 10665
rect 17543 10628 18644 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 18046 10588 18052 10600
rect 17420 10560 18052 10588
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 18616 10588 18644 10628
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 22066 10628 22201 10656
rect 18782 10588 18788 10600
rect 18616 10560 18788 10588
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 19720 10520 19748 10551
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 21450 10588 21456 10600
rect 20772 10560 21456 10588
rect 20772 10548 20778 10560
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 22066 10520 22094 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22554 10616 22560 10668
rect 22612 10656 22618 10668
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22612 10628 23121 10656
rect 22612 10616 22618 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10656 24179 10659
rect 24578 10656 24584 10668
rect 24167 10628 24584 10656
rect 24167 10625 24179 10628
rect 24121 10619 24179 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 24854 10656 24860 10668
rect 24688 10628 24860 10656
rect 22646 10548 22652 10600
rect 22704 10588 22710 10600
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 22704 10560 23397 10588
rect 22704 10548 22710 10560
rect 23385 10557 23397 10560
rect 23431 10588 23443 10591
rect 24688 10588 24716 10628
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 23431 10560 24716 10588
rect 23431 10557 23443 10560
rect 23385 10551 23443 10557
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 23474 10520 23480 10532
rect 16908 10492 19748 10520
rect 21008 10492 22094 10520
rect 22204 10492 23480 10520
rect 16908 10480 16914 10492
rect 13412 10424 16252 10452
rect 13412 10412 13418 10424
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 16448 10424 17601 10452
rect 16448 10412 16454 10424
rect 17589 10421 17601 10424
rect 17635 10421 17647 10455
rect 17589 10415 17647 10421
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 21008 10452 21036 10492
rect 19392 10424 21036 10452
rect 19392 10412 19398 10424
rect 22002 10412 22008 10464
rect 22060 10412 22066 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22204 10452 22232 10492
rect 23474 10480 23480 10492
rect 23532 10480 23538 10532
rect 22152 10424 22232 10452
rect 22741 10455 22799 10461
rect 22152 10412 22158 10424
rect 22741 10421 22753 10455
rect 22787 10452 22799 10455
rect 23566 10452 23572 10464
rect 22787 10424 23572 10452
rect 22787 10421 22799 10424
rect 22741 10415 22799 10421
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 13354 10248 13360 10260
rect 11655 10220 13360 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13446 10208 13452 10260
rect 13504 10208 13510 10260
rect 14550 10208 14556 10260
rect 14608 10208 14614 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 22554 10248 22560 10260
rect 18012 10220 22560 10248
rect 18012 10208 18018 10220
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 24578 10208 24584 10260
rect 24636 10208 24642 10260
rect 10870 10140 10876 10192
rect 10928 10180 10934 10192
rect 10928 10152 12204 10180
rect 10928 10140 10934 10152
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8260 10084 9321 10112
rect 8260 10072 8266 10084
rect 9309 10081 9321 10084
rect 9355 10112 9367 10115
rect 9582 10112 9588 10124
rect 9355 10084 9588 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 11422 10072 11428 10124
rect 11480 10112 11486 10124
rect 12176 10121 12204 10152
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 12805 10183 12863 10189
rect 12805 10180 12817 10183
rect 12400 10152 12817 10180
rect 12400 10140 12406 10152
rect 12805 10149 12817 10152
rect 12851 10149 12863 10183
rect 13464 10180 13492 10208
rect 15470 10180 15476 10192
rect 12805 10143 12863 10149
rect 13280 10152 15476 10180
rect 13280 10121 13308 10152
rect 15470 10140 15476 10152
rect 15528 10140 15534 10192
rect 18141 10183 18199 10189
rect 18141 10149 18153 10183
rect 18187 10149 18199 10183
rect 18141 10143 18199 10149
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11480 10084 12081 10112
rect 11480 10072 11486 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 14976 10084 15117 10112
rect 14976 10072 14982 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 17862 10112 17868 10124
rect 17368 10084 17868 10112
rect 17368 10072 17374 10084
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 18156 10112 18184 10143
rect 18230 10140 18236 10192
rect 18288 10140 18294 10192
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 22094 10180 22100 10192
rect 18472 10152 22100 10180
rect 18472 10140 18478 10152
rect 22094 10140 22100 10152
rect 22152 10140 22158 10192
rect 18064 10084 18184 10112
rect 18248 10112 18276 10140
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18248 10084 18613 10112
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 17681 10047 17739 10053
rect 17681 10044 17693 10047
rect 13780 10016 17693 10044
rect 13780 10004 13786 10016
rect 17681 10013 17693 10016
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9088 9948 9597 9976
rect 9088 9936 9094 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 10594 9936 10600 9988
rect 10652 9936 10658 9988
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 11204 9948 13185 9976
rect 11204 9936 11210 9948
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 13173 9939 13231 9945
rect 15013 9979 15071 9985
rect 15013 9945 15025 9979
rect 15059 9976 15071 9979
rect 15286 9976 15292 9988
rect 15059 9948 15292 9976
rect 15059 9945 15071 9948
rect 15013 9939 15071 9945
rect 15286 9936 15292 9948
rect 15344 9936 15350 9988
rect 16853 9979 16911 9985
rect 16853 9945 16865 9979
rect 16899 9976 16911 9979
rect 17586 9976 17592 9988
rect 16899 9948 17592 9976
rect 16899 9945 16911 9948
rect 16853 9939 16911 9945
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 18064 9976 18092 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 20070 10112 20076 10124
rect 18831 10084 20076 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 21361 10115 21419 10121
rect 21361 10112 21373 10115
rect 21232 10084 21373 10112
rect 21232 10072 21238 10084
rect 21361 10081 21373 10084
rect 21407 10081 21419 10115
rect 21361 10075 21419 10081
rect 21450 10072 21456 10124
rect 21508 10072 21514 10124
rect 22278 10072 22284 10124
rect 22336 10072 22342 10124
rect 22557 10115 22615 10121
rect 22557 10081 22569 10115
rect 22603 10112 22615 10115
rect 22646 10112 22652 10124
rect 22603 10084 22652 10112
rect 22603 10081 22615 10084
rect 22557 10075 22615 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20806 10044 20812 10056
rect 20303 10016 20812 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 21266 10004 21272 10056
rect 21324 10004 21330 10056
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23842 10004 23848 10056
rect 23900 10044 23906 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 23900 10016 24777 10044
rect 23900 10004 23906 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 19426 9976 19432 9988
rect 18064 9948 19432 9976
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 19521 9979 19579 9985
rect 19521 9945 19533 9979
rect 19567 9976 19579 9979
rect 20530 9976 20536 9988
rect 19567 9948 20536 9976
rect 19567 9945 19579 9948
rect 19521 9939 19579 9945
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 22646 9976 22652 9988
rect 20916 9948 22652 9976
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 14826 9908 14832 9920
rect 7156 9880 14832 9908
rect 7156 9868 7162 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15102 9908 15108 9920
rect 14967 9880 15108 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15102 9868 15108 9880
rect 15160 9908 15166 9920
rect 16482 9908 16488 9920
rect 15160 9880 16488 9908
rect 15160 9868 15166 9880
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17494 9868 17500 9920
rect 17552 9868 17558 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 18104 9880 18521 9908
rect 18104 9868 18110 9880
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18509 9871 18567 9877
rect 18782 9868 18788 9920
rect 18840 9908 18846 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 18840 9880 19625 9908
rect 18840 9868 18846 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 20916 9917 20944 9948
rect 22646 9936 22652 9948
rect 22704 9936 22710 9988
rect 20349 9911 20407 9917
rect 20349 9908 20361 9911
rect 19760 9880 20361 9908
rect 19760 9868 19766 9880
rect 20349 9877 20361 9880
rect 20395 9877 20407 9911
rect 20349 9871 20407 9877
rect 20901 9911 20959 9917
rect 20901 9877 20913 9911
rect 20947 9877 20959 9911
rect 20901 9871 20959 9877
rect 22830 9868 22836 9920
rect 22888 9908 22894 9920
rect 24029 9911 24087 9917
rect 24029 9908 24041 9911
rect 22888 9880 24041 9908
rect 22888 9868 22894 9880
rect 24029 9877 24041 9880
rect 24075 9877 24087 9911
rect 24029 9871 24087 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 15286 9704 15292 9716
rect 9824 9676 15292 9704
rect 9824 9664 9830 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 17310 9704 17316 9716
rect 17144 9676 17316 9704
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 14369 9639 14427 9645
rect 10652 9608 12466 9636
rect 10652 9596 10658 9608
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 14550 9636 14556 9648
rect 14415 9608 14556 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 15657 9639 15715 9645
rect 15657 9636 15669 9639
rect 15028 9608 15669 9636
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 10836 9472 11713 9500
rect 10836 9460 10842 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12526 9500 12532 9512
rect 12023 9472 12532 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 14274 9500 14280 9512
rect 13495 9472 14280 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 14918 9500 14924 9512
rect 14691 9472 14924 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15028 9432 15056 9608
rect 15657 9605 15669 9608
rect 15703 9636 15715 9639
rect 17144 9636 17172 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 22186 9704 22192 9716
rect 17552 9676 22192 9704
rect 17552 9664 17558 9676
rect 22186 9664 22192 9676
rect 22244 9664 22250 9716
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 24394 9704 24400 9716
rect 22704 9676 24400 9704
rect 22704 9664 22710 9676
rect 24394 9664 24400 9676
rect 24452 9664 24458 9716
rect 17862 9636 17868 9648
rect 15703 9608 17172 9636
rect 17236 9608 17868 9636
rect 15703 9605 15715 9608
rect 15657 9599 15715 9605
rect 17236 9577 17264 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 18598 9596 18604 9648
rect 18656 9596 18662 9648
rect 19978 9596 19984 9648
rect 20036 9636 20042 9648
rect 20346 9636 20352 9648
rect 20036 9608 20352 9636
rect 20036 9596 20042 9608
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 17221 9571 17279 9577
rect 15611 9540 17172 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 17144 9500 17172 9540
rect 17221 9537 17233 9571
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19300 9540 20269 9568
rect 19300 9528 19306 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 23382 9568 23388 9580
rect 22327 9540 23388 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 24118 9528 24124 9580
rect 24176 9528 24182 9580
rect 17494 9500 17500 9512
rect 17144 9472 17500 9500
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17681 9503 17739 9509
rect 17681 9469 17693 9503
rect 17727 9469 17739 9503
rect 17681 9463 17739 9469
rect 17957 9503 18015 9509
rect 17957 9469 17969 9503
rect 18003 9500 18015 9503
rect 20162 9500 20168 9512
rect 18003 9472 20168 9500
rect 18003 9469 18015 9472
rect 17957 9463 18015 9469
rect 13924 9404 15056 9432
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 13924 9364 13952 9404
rect 15194 9392 15200 9444
rect 15252 9392 15258 9444
rect 15764 9432 15792 9460
rect 17310 9432 17316 9444
rect 15764 9404 17316 9432
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 12400 9336 13952 9364
rect 12400 9324 12406 9336
rect 13998 9324 14004 9376
rect 14056 9324 14062 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 17126 9364 17132 9376
rect 14792 9336 17132 9364
rect 14792 9324 14798 9336
rect 17126 9324 17132 9336
rect 17184 9364 17190 9376
rect 17494 9364 17500 9376
rect 17184 9336 17500 9364
rect 17184 9324 17190 9336
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17696 9364 17724 9463
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 20349 9503 20407 9509
rect 20349 9469 20361 9503
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 22554 9500 22560 9512
rect 20579 9472 22560 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 20254 9432 20260 9444
rect 18984 9404 20260 9432
rect 18984 9364 19012 9404
rect 20254 9392 20260 9404
rect 20312 9392 20318 9444
rect 20364 9432 20392 9463
rect 22554 9460 22560 9472
rect 22612 9500 22618 9512
rect 22830 9500 22836 9512
rect 22612 9472 22836 9500
rect 22612 9460 22618 9472
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 23293 9503 23351 9509
rect 23293 9469 23305 9503
rect 23339 9500 23351 9503
rect 23566 9500 23572 9512
rect 23339 9472 23572 9500
rect 23339 9469 23351 9472
rect 23293 9463 23351 9469
rect 23566 9460 23572 9472
rect 23624 9460 23630 9512
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 20622 9432 20628 9444
rect 20364 9404 20628 9432
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 22370 9432 22376 9444
rect 22244 9404 22376 9432
rect 22244 9392 22250 9404
rect 22370 9392 22376 9404
rect 22428 9392 22434 9444
rect 17696 9336 19012 9364
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19116 9336 19441 9364
rect 19116 9324 19122 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 19886 9324 19892 9376
rect 19944 9324 19950 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20036 9336 21281 9364
rect 20036 9324 20042 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11606 9120 11612 9172
rect 11664 9120 11670 9172
rect 16482 9160 16488 9172
rect 13280 9132 16488 9160
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 10744 9064 13001 9092
rect 10744 9052 10750 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 10778 9024 10784 9036
rect 9180 8996 10784 9024
rect 9180 8984 9186 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 12124 8996 12173 9024
rect 12124 8984 12130 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 13280 9024 13308 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 19242 9160 19248 9172
rect 16724 9132 19248 9160
rect 16724 9120 16730 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 19886 9120 19892 9172
rect 19944 9160 19950 9172
rect 21726 9160 21732 9172
rect 19944 9132 21732 9160
rect 19944 9120 19950 9132
rect 21726 9120 21732 9132
rect 21784 9120 21790 9172
rect 13354 9052 13360 9104
rect 13412 9092 13418 9104
rect 17129 9095 17187 9101
rect 17129 9092 17141 9095
rect 13412 9064 17141 9092
rect 13412 9052 13418 9064
rect 17129 9061 17141 9064
rect 17175 9061 17187 9095
rect 17129 9055 17187 9061
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 18693 9095 18751 9101
rect 17368 9064 17724 9092
rect 17368 9052 17374 9064
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 13280 8996 13461 9024
rect 12161 8987 12219 8993
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 13688 8996 14872 9024
rect 13688 8984 13694 8996
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 13998 8956 14004 8968
rect 12023 8928 14004 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14844 8956 14872 8996
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 16114 8984 16120 9036
rect 16172 9024 16178 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16172 8996 16497 9024
rect 16172 8984 16178 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 17696 9033 17724 9064
rect 18693 9061 18705 9095
rect 18739 9092 18751 9095
rect 24670 9092 24676 9104
rect 18739 9064 24676 9092
rect 18739 9061 18751 9064
rect 18693 9055 18751 9061
rect 24670 9052 24676 9064
rect 24728 9052 24734 9104
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17552 8996 17601 9024
rect 17552 8984 17558 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 17681 9027 17739 9033
rect 17681 8993 17693 9027
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 20073 9027 20131 9033
rect 20073 9024 20085 9027
rect 19484 8996 20085 9024
rect 19484 8984 19490 8996
rect 20073 8993 20085 8996
rect 20119 8993 20131 9027
rect 20073 8987 20131 8993
rect 20162 8984 20168 9036
rect 20220 8984 20226 9036
rect 15930 8956 15936 8968
rect 14844 8928 15936 8956
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 17126 8956 17132 8968
rect 16347 8928 17132 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 18874 8916 18880 8968
rect 18932 8916 18938 8968
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19300 8928 19932 8956
rect 19300 8916 19306 8928
rect 18877 8915 18935 8916
rect 9401 8891 9459 8897
rect 9401 8857 9413 8891
rect 9447 8888 9459 8891
rect 9674 8888 9680 8900
rect 9447 8860 9680 8888
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 10686 8888 10692 8900
rect 10626 8860 10692 8888
rect 10686 8848 10692 8860
rect 10744 8848 10750 8900
rect 12069 8891 12127 8897
rect 12069 8857 12081 8891
rect 12115 8888 12127 8891
rect 12115 8860 14320 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 10870 8780 10876 8832
rect 10928 8780 10934 8832
rect 13354 8780 13360 8832
rect 13412 8780 13418 8832
rect 14292 8829 14320 8860
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 14516 8860 14749 8888
rect 14516 8848 14522 8860
rect 14737 8857 14749 8860
rect 14783 8857 14795 8891
rect 14737 8851 14795 8857
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19518 8888 19524 8900
rect 19116 8860 19524 8888
rect 19116 8848 19122 8860
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8789 14335 8823
rect 14277 8783 14335 8789
rect 14642 8780 14648 8832
rect 14700 8780 14706 8832
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8820 16451 8823
rect 16666 8820 16672 8832
rect 16439 8792 16672 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 17497 8823 17555 8829
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 19242 8820 19248 8832
rect 17543 8792 19248 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19484 8792 19625 8820
rect 19484 8780 19490 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19904 8820 19932 8928
rect 19978 8916 19984 8968
rect 20036 8916 20042 8968
rect 20806 8916 20812 8968
rect 20864 8916 20870 8968
rect 20898 8916 20904 8968
rect 20956 8956 20962 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 20956 8928 22661 8956
rect 20956 8916 20962 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 22738 8916 22744 8968
rect 22796 8956 22802 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 22796 8928 24777 8956
rect 22796 8916 22802 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 21818 8848 21824 8900
rect 21876 8848 21882 8900
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 22002 8820 22008 8832
rect 19904 8792 22008 8820
rect 19613 8783 19671 8789
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 24578 8780 24584 8832
rect 24636 8780 24642 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 14090 8616 14096 8628
rect 12216 8588 14096 8616
rect 12216 8576 12222 8588
rect 14090 8576 14096 8588
rect 14148 8616 14154 8628
rect 14458 8616 14464 8628
rect 14148 8588 14464 8616
rect 14148 8576 14154 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 18877 8619 18935 8625
rect 18877 8616 18889 8619
rect 16899 8588 18889 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 18877 8585 18889 8588
rect 18923 8585 18935 8619
rect 18877 8579 18935 8585
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21453 8619 21511 8625
rect 21453 8616 21465 8619
rect 20220 8588 21465 8616
rect 20220 8576 20226 8588
rect 21453 8585 21465 8588
rect 21499 8585 21511 8619
rect 21453 8579 21511 8585
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 11514 8548 11520 8560
rect 7708 8520 11520 8548
rect 7708 8508 7714 8520
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 13872 8520 13921 8548
rect 13872 8508 13878 8520
rect 13909 8517 13921 8520
rect 13955 8517 13967 8551
rect 19886 8548 19892 8560
rect 13909 8511 13967 8517
rect 17052 8520 19564 8548
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11195 8452 12081 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 14734 8480 14740 8492
rect 12069 8443 12127 8449
rect 12360 8452 14740 8480
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 12360 8421 12388 8452
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 14826 8440 14832 8492
rect 14884 8440 14890 8492
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 17052 8480 17080 8520
rect 15151 8452 17080 8480
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 17184 8452 17233 8480
rect 17184 8440 17190 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17678 8480 17684 8492
rect 17552 8452 17684 8480
rect 17552 8440 17558 8452
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 2280 8384 12173 8412
rect 2280 8372 2286 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 16666 8412 16672 8424
rect 12345 8375 12403 8381
rect 14016 8384 16672 8412
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 14016 8344 14044 8384
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 17000 8384 17325 8412
rect 17000 8372 17006 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 11204 8316 14044 8344
rect 11204 8304 11210 8316
rect 14090 8304 14096 8356
rect 14148 8304 14154 8356
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 14700 8316 16313 8344
rect 14700 8304 14706 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 16301 8307 16359 8313
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 17420 8344 17448 8375
rect 18800 8344 18828 8443
rect 18966 8372 18972 8424
rect 19024 8372 19030 8424
rect 19536 8412 19564 8520
rect 19720 8520 19892 8548
rect 19720 8489 19748 8520
rect 19886 8508 19892 8520
rect 19944 8548 19950 8560
rect 20254 8548 20260 8560
rect 19944 8520 20260 8548
rect 19944 8508 19950 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22462 8480 22468 8492
rect 22327 8452 22468 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23532 8452 23949 8480
rect 23532 8440 23538 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 20714 8412 20720 8424
rect 19536 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 21100 8412 21128 8440
rect 21266 8412 21272 8424
rect 21100 8384 21272 8412
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 22370 8372 22376 8424
rect 22428 8412 22434 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22428 8384 22569 8412
rect 22428 8372 22434 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 19334 8344 19340 8356
rect 17184 8316 17448 8344
rect 17972 8316 18828 8344
rect 18892 8316 19340 8344
rect 17184 8304 17190 8316
rect 13354 8236 13360 8288
rect 13412 8236 13418 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 17972 8276 18000 8316
rect 13504 8248 18000 8276
rect 18417 8279 18475 8285
rect 13504 8236 13510 8248
rect 18417 8245 18429 8279
rect 18463 8276 18475 8279
rect 18892 8276 18920 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 19978 8285 19984 8288
rect 18463 8248 18920 8276
rect 19968 8279 19984 8285
rect 18463 8245 18475 8248
rect 18417 8239 18475 8245
rect 19968 8245 19980 8279
rect 19968 8239 19984 8245
rect 19978 8236 19984 8239
rect 20036 8236 20042 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 13722 8072 13728 8084
rect 11839 8044 13728 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14323 8044 15884 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 10321 8007 10379 8013
rect 10321 7973 10333 8007
rect 10367 8004 10379 8007
rect 12066 8004 12072 8016
rect 10367 7976 12072 8004
rect 10367 7973 10379 7976
rect 10321 7967 10379 7973
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 15856 8004 15884 8044
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 16761 8075 16819 8081
rect 16761 8072 16773 8075
rect 16540 8044 16773 8072
rect 16540 8032 16546 8044
rect 16761 8041 16773 8044
rect 16807 8041 16819 8075
rect 16761 8035 16819 8041
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18874 8072 18880 8084
rect 18380 8044 18880 8072
rect 18380 8032 18386 8044
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 22186 8072 22192 8084
rect 22066 8044 22192 8072
rect 17402 8004 17408 8016
rect 12584 7976 14872 8004
rect 15856 7976 17408 8004
rect 12584 7964 12590 7976
rect 10870 7896 10876 7948
rect 10928 7896 10934 7948
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 14844 7945 14872 7976
rect 17402 7964 17408 7976
rect 17460 7964 17466 8016
rect 18141 8007 18199 8013
rect 18141 7973 18153 8007
rect 18187 8004 18199 8007
rect 20990 8004 20996 8016
rect 18187 7976 20996 8004
rect 18187 7973 18199 7976
rect 18141 7967 18199 7973
rect 20990 7964 20996 7976
rect 21048 7964 21054 8016
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 11020 7908 12357 7936
rect 11020 7896 11026 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 13633 7939 13691 7945
rect 12345 7899 12403 7905
rect 13280 7908 13492 7936
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 13280 7868 13308 7908
rect 10827 7840 13308 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13464 7868 13492 7908
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14829 7939 14887 7945
rect 13679 7908 14780 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14458 7868 14464 7880
rect 13464 7840 14464 7868
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 14752 7868 14780 7908
rect 14829 7905 14841 7939
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7936 15531 7939
rect 16206 7936 16212 7948
rect 15519 7908 16212 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 17310 7896 17316 7948
rect 17368 7896 17374 7948
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7936 18843 7939
rect 19518 7936 19524 7948
rect 18831 7908 19524 7936
rect 18831 7905 18843 7908
rect 18785 7899 18843 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 22066 7936 22094 8044
rect 22186 8032 22192 8044
rect 22244 8072 22250 8084
rect 22244 8044 23612 8072
rect 22244 8032 22250 8044
rect 23584 8004 23612 8044
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24176 8044 24685 8072
rect 24176 8032 24182 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 24210 8004 24216 8016
rect 23584 7976 24216 8004
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 19628 7908 22094 7936
rect 15010 7868 15016 7880
rect 14752 7840 15016 7868
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15746 7828 15752 7880
rect 15804 7828 15810 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 19628 7868 19656 7908
rect 22278 7896 22284 7948
rect 22336 7896 22342 7948
rect 22554 7896 22560 7948
rect 22612 7896 22618 7948
rect 23842 7936 23848 7948
rect 23676 7908 23848 7936
rect 23676 7880 23704 7908
rect 23842 7896 23848 7908
rect 23900 7896 23906 7948
rect 17175 7840 19656 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 20732 7840 21772 7868
rect 5258 7760 5264 7812
rect 5316 7800 5322 7812
rect 11330 7800 11336 7812
rect 5316 7772 11336 7800
rect 5316 7760 5322 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7800 12219 7803
rect 12207 7772 12434 7800
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10318 7732 10324 7744
rect 10100 7704 10324 7732
rect 10100 7692 10106 7704
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10502 7692 10508 7744
rect 10560 7732 10566 7744
rect 10689 7735 10747 7741
rect 10689 7732 10701 7735
rect 10560 7704 10701 7732
rect 10560 7692 10566 7704
rect 10689 7701 10701 7704
rect 10735 7701 10747 7735
rect 10689 7695 10747 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12124 7704 12265 7732
rect 12124 7692 12130 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12406 7732 12434 7772
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 13449 7803 13507 7809
rect 13449 7800 13461 7803
rect 12768 7772 13461 7800
rect 12768 7760 12774 7772
rect 13449 7769 13461 7772
rect 13495 7769 13507 7803
rect 13449 7763 13507 7769
rect 14274 7760 14280 7812
rect 14332 7800 14338 7812
rect 16942 7800 16948 7812
rect 14332 7772 16948 7800
rect 14332 7760 14338 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 18509 7803 18567 7809
rect 18509 7800 18521 7803
rect 17328 7772 18521 7800
rect 17328 7744 17356 7772
rect 18509 7769 18521 7772
rect 18555 7769 18567 7803
rect 18509 7763 18567 7769
rect 18874 7760 18880 7812
rect 18932 7800 18938 7812
rect 19521 7803 19579 7809
rect 19521 7800 19533 7803
rect 18932 7772 19533 7800
rect 18932 7760 18938 7772
rect 19521 7769 19533 7772
rect 19567 7769 19579 7803
rect 19521 7763 19579 7769
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 20162 7800 20168 7812
rect 19751 7772 20168 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 12802 7732 12808 7744
rect 12406 7704 12808 7732
rect 12253 7695 12311 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12952 7704 13001 7732
rect 12952 7692 12958 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 17221 7735 17279 7741
rect 17221 7701 17233 7735
rect 17267 7732 17279 7735
rect 17310 7732 17316 7744
rect 17267 7704 17316 7732
rect 17267 7701 17279 7704
rect 17221 7695 17279 7701
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 18601 7735 18659 7741
rect 18601 7732 18613 7735
rect 17552 7704 18613 7732
rect 17552 7692 17558 7704
rect 18601 7701 18613 7704
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 20732 7732 20760 7840
rect 21634 7760 21640 7812
rect 21692 7760 21698 7812
rect 21744 7800 21772 7840
rect 23658 7828 23664 7880
rect 23716 7828 23722 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 23860 7840 24869 7868
rect 21744 7772 22508 7800
rect 19392 7704 20760 7732
rect 22480 7732 22508 7772
rect 23860 7732 23888 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 22480 7704 23888 7732
rect 19392 7692 19398 7704
rect 24026 7692 24032 7744
rect 24084 7692 24090 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 10689 7531 10747 7537
rect 6788 7500 10548 7528
rect 6788 7488 6794 7500
rect 10520 7460 10548 7500
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 10962 7528 10968 7540
rect 10735 7500 10968 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 14734 7528 14740 7540
rect 11747 7500 14740 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 15804 7500 23980 7528
rect 15804 7488 15810 7500
rect 12069 7463 12127 7469
rect 12069 7460 12081 7463
rect 10520 7432 12081 7460
rect 12069 7429 12081 7432
rect 12115 7429 12127 7463
rect 12069 7423 12127 7429
rect 12161 7463 12219 7469
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 14274 7460 14280 7472
rect 12207 7432 14280 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 15010 7420 15016 7472
rect 15068 7420 15074 7472
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 16117 7463 16175 7469
rect 16117 7460 16129 7463
rect 15620 7432 16129 7460
rect 15620 7420 15626 7432
rect 16117 7429 16129 7432
rect 16163 7429 16175 7463
rect 16117 7423 16175 7429
rect 17034 7420 17040 7472
rect 17092 7420 17098 7472
rect 18414 7420 18420 7472
rect 18472 7420 18478 7472
rect 10686 7392 10692 7404
rect 10350 7364 10692 7392
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13446 7392 13452 7404
rect 13311 7364 13452 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 17494 7392 17500 7404
rect 15804 7364 17500 7392
rect 15804 7352 15810 7364
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19300 7364 20085 7392
rect 19300 7352 19306 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 23952 7401 23980 7500
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 20772 7364 22109 7392
rect 20772 7352 20778 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9217 7327 9275 7333
rect 8987 7296 9076 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9048 7188 9076 7296
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 10870 7324 10876 7336
rect 9263 7296 10876 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11698 7324 11704 7336
rect 11112 7296 11704 7324
rect 11112 7284 11118 7296
rect 11698 7284 11704 7296
rect 11756 7324 11762 7336
rect 12253 7327 12311 7333
rect 12253 7324 12265 7327
rect 11756 7296 12265 7324
rect 11756 7284 11762 7296
rect 12253 7293 12265 7296
rect 12299 7293 12311 7327
rect 12253 7287 12311 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 14001 7327 14059 7333
rect 13771 7296 13860 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 9582 7188 9588 7200
rect 9048 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 13832 7188 13860 7296
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 16298 7324 16304 7336
rect 14047 7296 16304 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 16908 7296 17693 7324
rect 16908 7284 16914 7296
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7324 18015 7327
rect 18598 7324 18604 7336
rect 18003 7296 18604 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 18598 7284 18604 7296
rect 18656 7324 18662 7336
rect 18966 7324 18972 7336
rect 18656 7296 18972 7324
rect 18656 7284 18662 7296
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7324 19487 7327
rect 19610 7324 19616 7336
rect 19475 7296 19616 7324
rect 19475 7293 19487 7296
rect 19429 7287 19487 7293
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21910 7324 21916 7336
rect 21315 7296 21916 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21910 7284 21916 7296
rect 21968 7284 21974 7336
rect 23290 7284 23296 7336
rect 23348 7284 23354 7336
rect 16868 7256 16896 7284
rect 15028 7228 16896 7256
rect 15028 7188 15056 7228
rect 17218 7216 17224 7268
rect 17276 7216 17282 7268
rect 20622 7216 20628 7268
rect 20680 7256 20686 7268
rect 24854 7256 24860 7268
rect 20680 7228 24860 7256
rect 20680 7216 20686 7228
rect 24854 7216 24860 7228
rect 24912 7216 24918 7268
rect 13832 7160 15056 7188
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15160 7160 15485 7188
rect 15160 7148 15166 7160
rect 15473 7157 15485 7160
rect 15519 7157 15531 7191
rect 15473 7151 15531 7157
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 16482 7188 16488 7200
rect 16255 7160 16488 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 18690 7188 18696 7200
rect 18380 7160 18696 7188
rect 18380 7148 18386 7160
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 19242 6984 19248 6996
rect 13872 6956 19248 6984
rect 13872 6944 13878 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20152 6987 20210 6993
rect 20152 6953 20164 6987
rect 20198 6984 20210 6987
rect 21450 6984 21456 6996
rect 20198 6956 21456 6984
rect 20198 6953 20210 6956
rect 20152 6947 20210 6953
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 22094 6984 22100 6996
rect 22066 6944 22100 6984
rect 22152 6944 22158 6996
rect 22360 6987 22418 6993
rect 22360 6953 22372 6987
rect 22406 6984 22418 6987
rect 24026 6984 24032 6996
rect 22406 6956 24032 6984
rect 22406 6953 22418 6956
rect 22360 6947 22418 6953
rect 24026 6944 24032 6956
rect 24084 6944 24090 6996
rect 15102 6916 15108 6928
rect 13648 6888 15108 6916
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 8846 6848 8852 6860
rect 5500 6820 8852 6848
rect 5500 6808 5506 6820
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 11054 6808 11060 6860
rect 11112 6808 11118 6860
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13648 6857 13676 6888
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13412 6820 13645 6848
rect 13412 6808 13418 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 14384 6820 15424 6848
rect 10778 6740 10784 6792
rect 10836 6740 10842 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13722 6780 13728 6792
rect 13495 6752 13728 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 10744 6684 11546 6712
rect 12406 6684 13369 6712
rect 10744 6672 10750 6684
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 12406 6644 12434 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13357 6675 13415 6681
rect 9732 6616 12434 6644
rect 12989 6647 13047 6653
rect 9732 6604 9738 6616
rect 12989 6613 13001 6647
rect 13035 6644 13047 6647
rect 13262 6644 13268 6656
rect 13035 6616 13268 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14384 6653 14412 6820
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15286 6780 15292 6792
rect 14599 6752 15292 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 15396 6780 15424 6820
rect 15470 6808 15476 6860
rect 15528 6848 15534 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15528 6820 15577 6848
rect 15528 6808 15534 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17034 6848 17040 6860
rect 16991 6820 17040 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 18690 6848 18696 6860
rect 17696 6820 18696 6848
rect 17696 6789 17724 6820
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 19886 6808 19892 6860
rect 19944 6848 19950 6860
rect 22066 6857 22094 6944
rect 24044 6916 24072 6944
rect 24044 6888 25176 6916
rect 25148 6857 25176 6888
rect 22066 6851 22144 6857
rect 22066 6848 22098 6851
rect 19944 6820 22098 6848
rect 19944 6808 19950 6820
rect 22086 6817 22098 6820
rect 22132 6817 22144 6851
rect 22086 6811 22144 6817
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 17681 6783 17739 6789
rect 15396 6752 17632 6780
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 15028 6684 16773 6712
rect 15028 6653 15056 6684
rect 16761 6681 16773 6684
rect 16807 6681 16819 6715
rect 17604 6712 17632 6752
rect 17681 6749 17693 6783
rect 17727 6749 17739 6783
rect 19334 6780 19340 6792
rect 17681 6743 17739 6749
rect 18248 6752 19340 6780
rect 18248 6712 18276 6752
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 23658 6780 23664 6792
rect 23506 6752 23664 6780
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 17604 6684 18276 6712
rect 18693 6715 18751 6721
rect 16761 6675 16819 6681
rect 18693 6681 18705 6715
rect 18739 6712 18751 6715
rect 20438 6712 20444 6724
rect 18739 6684 20444 6712
rect 18739 6681 18751 6684
rect 18693 6675 18751 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 25041 6715 25099 6721
rect 25041 6712 25053 6715
rect 23676 6684 25053 6712
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6613 15071 6647
rect 15013 6607 15071 6613
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 15252 6616 15393 6644
rect 15252 6604 15258 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15381 6607 15439 6613
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 15562 6644 15568 6656
rect 15519 6616 15568 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 16022 6604 16028 6656
rect 16080 6644 16086 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16080 6616 16313 6644
rect 16080 6604 16086 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 16669 6647 16727 6653
rect 16669 6613 16681 6647
rect 16715 6644 16727 6647
rect 19242 6644 19248 6656
rect 16715 6616 19248 6644
rect 16715 6613 16727 6616
rect 16669 6607 16727 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 21637 6647 21695 6653
rect 21637 6644 21649 6647
rect 20036 6616 21649 6644
rect 20036 6604 20042 6616
rect 21637 6613 21649 6616
rect 21683 6613 21695 6647
rect 21637 6607 21695 6613
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 23676 6644 23704 6684
rect 25041 6681 25053 6684
rect 25087 6681 25099 6715
rect 25041 6675 25099 6681
rect 21784 6616 23704 6644
rect 21784 6604 21790 6616
rect 23842 6604 23848 6656
rect 23900 6604 23906 6656
rect 24026 6604 24032 6656
rect 24084 6644 24090 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 24084 6616 24593 6644
rect 24084 6604 24090 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 24946 6604 24952 6656
rect 25004 6604 25010 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 13722 6440 13728 6452
rect 12492 6412 13728 6440
rect 12492 6400 12498 6412
rect 13722 6400 13728 6412
rect 13780 6440 13786 6452
rect 15194 6440 15200 6452
rect 13780 6412 15200 6440
rect 13780 6400 13786 6412
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17460 6412 18552 6440
rect 17460 6400 17466 6412
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 15749 6375 15807 6381
rect 15749 6372 15761 6375
rect 13320 6344 15761 6372
rect 13320 6332 13326 6344
rect 15749 6341 15761 6344
rect 15795 6341 15807 6375
rect 18414 6372 18420 6384
rect 18354 6344 18420 6372
rect 15749 6335 15807 6341
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 12802 6264 12808 6316
rect 12860 6304 12866 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12860 6276 13001 6304
rect 12860 6264 12866 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 13814 6304 13820 6316
rect 13771 6276 13820 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 18524 6304 18552 6412
rect 18598 6400 18604 6452
rect 18656 6400 18662 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 23842 6440 23848 6452
rect 19576 6412 23848 6440
rect 19576 6400 19582 6412
rect 23842 6400 23848 6412
rect 23900 6400 23906 6452
rect 21269 6375 21327 6381
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 22554 6372 22560 6384
rect 21315 6344 22560 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 25130 6332 25136 6384
rect 25188 6332 25194 6384
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 18524 6276 19257 6304
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 21726 6264 21732 6316
rect 21784 6304 21790 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21784 6276 22017 6304
rect 21784 6264 21790 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 24578 6304 24584 6316
rect 24167 6276 24584 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 13446 6196 13452 6248
rect 13504 6196 13510 6248
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 14884 6208 15853 6236
rect 14884 6196 14890 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 16850 6196 16856 6248
rect 16908 6196 16914 6248
rect 17126 6196 17132 6248
rect 17184 6196 17190 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22152 6208 22477 6236
rect 22152 6196 22158 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 24026 6168 24032 6180
rect 18984 6140 24032 6168
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 18984 6100 19012 6140
rect 24026 6128 24032 6140
rect 24084 6128 24090 6180
rect 14516 6072 19012 6100
rect 19061 6103 19119 6109
rect 14516 6060 14522 6072
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 20346 6100 20352 6112
rect 19107 6072 20352 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 22830 6100 22836 6112
rect 20496 6072 22836 6100
rect 20496 6060 20502 6072
rect 22830 6060 22836 6072
rect 22888 6060 22894 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11698 5856 11704 5908
rect 11756 5856 11762 5908
rect 21726 5856 21732 5908
rect 21784 5896 21790 5908
rect 24673 5899 24731 5905
rect 24673 5896 24685 5899
rect 21784 5868 24685 5896
rect 21784 5856 21790 5868
rect 24673 5865 24685 5868
rect 24719 5865 24731 5899
rect 24673 5859 24731 5865
rect 20070 5828 20076 5840
rect 16776 5800 20076 5828
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 10962 5760 10968 5772
rect 10275 5732 10968 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 16776 5769 16804 5800
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5729 16819 5763
rect 20438 5760 20444 5772
rect 16761 5723 16819 5729
rect 17512 5732 20444 5760
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9640 5664 9965 5692
rect 9640 5652 9646 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13596 5664 13737 5692
rect 13596 5652 13602 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14936 5692 14964 5720
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14936 5664 15025 5692
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16114 5692 16120 5704
rect 15887 5664 16120 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 10686 5624 10692 5636
rect 10612 5596 10692 5624
rect 10612 5556 10640 5596
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 15197 5627 15255 5633
rect 12406 5596 15056 5624
rect 12406 5556 12434 5596
rect 15028 5568 15056 5596
rect 15197 5593 15209 5627
rect 15243 5624 15255 5627
rect 17512 5624 17540 5732
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22336 5732 22661 5760
rect 22336 5720 22342 5732
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 22649 5723 22707 5729
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 18598 5692 18604 5704
rect 17727 5664 18604 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5692 18751 5695
rect 19610 5692 19616 5704
rect 18739 5664 19616 5692
rect 18739 5661 18751 5664
rect 18693 5655 18751 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 20346 5652 20352 5704
rect 20404 5652 20410 5704
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 25038 5692 25044 5704
rect 24903 5664 25044 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 15243 5596 17540 5624
rect 15243 5593 15255 5596
rect 15197 5587 15255 5593
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 17644 5596 19533 5624
rect 17644 5584 17650 5596
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 19705 5627 19763 5633
rect 19705 5593 19717 5627
rect 19751 5624 19763 5627
rect 20622 5624 20628 5636
rect 19751 5596 20628 5624
rect 19751 5593 19763 5596
rect 19705 5587 19763 5593
rect 20622 5584 20628 5596
rect 20680 5584 20686 5636
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5593 21327 5627
rect 21269 5587 21327 5593
rect 10612 5528 12434 5556
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 14182 5556 14188 5568
rect 13587 5528 14188 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14274 5516 14280 5568
rect 14332 5516 14338 5568
rect 15010 5516 15016 5568
rect 15068 5516 15074 5568
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 21284 5556 21312 5587
rect 20404 5528 21312 5556
rect 20404 5516 20410 5528
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 14826 5312 14832 5364
rect 14884 5312 14890 5364
rect 22738 5352 22744 5364
rect 16868 5324 22744 5352
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 10410 5284 10416 5296
rect 3936 5256 10416 5284
rect 3936 5244 3942 5256
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 13354 5244 13360 5296
rect 13412 5244 13418 5296
rect 15010 5284 15016 5296
rect 14582 5256 15016 5284
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 16868 5216 16896 5324
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17129 5287 17187 5293
rect 17129 5284 17141 5287
rect 17092 5256 17141 5284
rect 17092 5244 17098 5256
rect 17129 5253 17141 5256
rect 17175 5253 17187 5287
rect 18414 5284 18420 5296
rect 18354 5256 18420 5284
rect 17129 5247 17187 5253
rect 18414 5244 18420 5256
rect 18472 5244 18478 5296
rect 19886 5284 19892 5296
rect 19720 5256 19892 5284
rect 15519 5188 16896 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 19242 5176 19248 5228
rect 19300 5176 19306 5228
rect 19720 5225 19748 5256
rect 19886 5244 19892 5256
rect 19944 5244 19950 5296
rect 21266 5284 21272 5296
rect 21206 5256 21272 5284
rect 21266 5244 21272 5256
rect 21324 5244 21330 5296
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 10836 5120 13093 5148
rect 10836 5108 10842 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 13096 5012 13124 5111
rect 15764 5080 15792 5111
rect 16850 5108 16856 5160
rect 16908 5108 16914 5160
rect 17126 5108 17132 5160
rect 17184 5148 17190 5160
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 17184 5120 18613 5148
rect 17184 5108 17190 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19576 5120 19993 5148
rect 19576 5108 19582 5120
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 20622 5108 20628 5160
rect 20680 5148 20686 5160
rect 22112 5148 22140 5179
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 20680 5120 22140 5148
rect 22465 5151 22523 5157
rect 20680 5108 20686 5120
rect 22465 5117 22477 5151
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 15764 5052 16988 5080
rect 13906 5012 13912 5024
rect 13096 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 15930 5012 15936 5024
rect 14516 4984 15936 5012
rect 14516 4972 14522 4984
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 16960 5012 16988 5052
rect 21450 5040 21456 5092
rect 21508 5040 21514 5092
rect 20622 5012 20628 5024
rect 16960 4984 20628 5012
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 22480 5012 22508 5111
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 21324 4984 22508 5012
rect 21324 4972 21330 4984
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 14737 4811 14795 4817
rect 14737 4777 14749 4811
rect 14783 4808 14795 4811
rect 15654 4808 15660 4820
rect 14783 4780 15660 4808
rect 14783 4777 14795 4780
rect 14737 4771 14795 4777
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16945 4811 17003 4817
rect 16264 4780 16896 4808
rect 16264 4768 16270 4780
rect 16868 4740 16896 4780
rect 16945 4777 16957 4811
rect 16991 4808 17003 4811
rect 17034 4808 17040 4820
rect 16991 4780 17040 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 23293 4811 23351 4817
rect 23293 4777 23305 4811
rect 23339 4808 23351 4811
rect 23382 4808 23388 4820
rect 23339 4780 23388 4808
rect 23339 4777 23351 4780
rect 23293 4771 23351 4777
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 23845 4743 23903 4749
rect 23845 4740 23857 4743
rect 16868 4712 23857 4740
rect 23845 4709 23857 4712
rect 23891 4709 23903 4743
rect 23845 4703 23903 4709
rect 24854 4700 24860 4752
rect 24912 4700 24918 4752
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9582 4672 9588 4684
rect 5123 4644 9588 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13630 4672 13636 4684
rect 13219 4644 13636 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 16850 4672 16856 4684
rect 15243 4644 16856 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17552 4644 17877 4672
rect 17552 4632 17558 4644
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 24394 4672 24400 4684
rect 20956 4644 22094 4672
rect 20956 4632 20962 4644
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12483 4576 12909 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 18782 4604 18788 4616
rect 17635 4576 18788 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 5350 4496 5356 4548
rect 5408 4496 5414 4548
rect 10686 4536 10692 4548
rect 6578 4508 10692 4536
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 12912 4536 12940 4567
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 19794 4604 19800 4616
rect 19659 4576 19800 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 21542 4604 21548 4616
rect 21499 4576 21548 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 22066 4604 22094 4644
rect 24136 4644 24400 4672
rect 23201 4607 23259 4613
rect 23201 4604 23213 4607
rect 22066 4576 23213 4604
rect 23201 4573 23213 4576
rect 23247 4573 23259 4607
rect 23201 4567 23259 4573
rect 24029 4607 24087 4613
rect 24029 4573 24041 4607
rect 24075 4604 24087 4607
rect 24136 4604 24164 4644
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 24075 4576 24164 4604
rect 24075 4573 24087 4576
rect 24029 4567 24087 4573
rect 24210 4564 24216 4616
rect 24268 4604 24274 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24268 4576 24685 4604
rect 24268 4564 24274 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 15378 4536 15384 4548
rect 12912 4508 15384 4536
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15470 4496 15476 4548
rect 15528 4496 15534 4548
rect 18414 4536 18420 4548
rect 16698 4508 18420 4536
rect 15010 4428 15016 4480
rect 15068 4468 15074 4480
rect 16776 4468 16804 4508
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 22189 4539 22247 4545
rect 22189 4536 22201 4539
rect 21140 4508 22201 4536
rect 21140 4496 21146 4508
rect 22189 4505 22201 4508
rect 22235 4505 22247 4539
rect 22189 4499 22247 4505
rect 15068 4440 16804 4468
rect 15068 4428 15074 4440
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 22462 4468 22468 4480
rect 19484 4440 22468 4468
rect 19484 4428 19490 4440
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 15528 4236 15669 4264
rect 15528 4224 15534 4236
rect 15657 4233 15669 4236
rect 15703 4233 15715 4267
rect 15657 4227 15715 4233
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 20220 4236 23888 4264
rect 20220 4224 20226 4236
rect 14918 4156 14924 4208
rect 14976 4156 14982 4208
rect 20898 4156 20904 4208
rect 20956 4156 20962 4208
rect 22646 4196 22652 4208
rect 22112 4168 22652 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1544 4100 1777 4128
rect 1544 4088 1550 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1912 4100 2421 4128
rect 1912 4088 1918 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 5960 4100 6745 4128
rect 5960 4088 5966 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16632 4100 16865 4128
rect 16632 4088 16638 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 17276 4100 18705 4128
rect 17276 4088 17282 4100
rect 18693 4097 18705 4100
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 22112 4137 22140 4168
rect 22646 4156 22652 4168
rect 22704 4156 22710 4208
rect 23860 4137 23888 4236
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14826 4060 14832 4072
rect 14231 4032 14832 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 2222 3952 2228 4004
rect 2280 3952 2286 4004
rect 4154 3952 4160 4004
rect 4212 3952 4218 4004
rect 6549 3995 6607 4001
rect 6549 3961 6561 3995
rect 6595 3992 6607 3995
rect 11790 3992 11796 4004
rect 6595 3964 11796 3992
rect 6595 3961 6607 3964
rect 6549 3955 6607 3961
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 5350 3924 5356 3936
rect 1627 3896 5356 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 13280 3924 13308 4023
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18380 4032 19165 4060
rect 18380 4020 18386 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 21450 4060 21456 4072
rect 21223 4032 21456 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22066 4032 22477 4060
rect 16114 3952 16120 4004
rect 16172 3952 16178 4004
rect 16850 3952 16856 4004
rect 16908 3992 16914 4004
rect 17678 3992 17684 4004
rect 16908 3964 17684 3992
rect 16908 3952 16914 3964
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 19978 3952 19984 4004
rect 20036 3992 20042 4004
rect 22066 3992 22094 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 20036 3964 22094 3992
rect 20036 3952 20042 3964
rect 18046 3924 18052 3936
rect 13280 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 18196 3896 20545 3924
rect 18196 3884 18202 3896
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20533 3887 20591 3893
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 24320 3924 24348 4023
rect 21048 3896 24348 3924
rect 21048 3884 21054 3896
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3326 3720 3332 3732
rect 2915 3692 3332 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4246 3680 4252 3732
rect 4304 3680 4310 3732
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 7800 3692 8217 3720
rect 7800 3680 7806 3692
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 8205 3683 8263 3689
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 13814 3720 13820 3732
rect 9723 3692 13820 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 17957 3723 18015 3729
rect 17957 3720 17969 3723
rect 16356 3692 17969 3720
rect 16356 3680 16362 3692
rect 17957 3689 17969 3692
rect 18003 3689 18015 3723
rect 17957 3683 18015 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 25130 3720 25136 3732
rect 18104 3692 25136 3720
rect 18104 3680 18110 3692
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 9398 3652 9404 3664
rect 1872 3624 9404 3652
rect 1872 3593 1900 3624
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 10413 3655 10471 3661
rect 10413 3621 10425 3655
rect 10459 3652 10471 3655
rect 15838 3652 15844 3664
rect 10459 3624 15844 3652
rect 10459 3621 10471 3624
rect 10413 3615 10471 3621
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 19886 3652 19892 3664
rect 18840 3624 19892 3652
rect 18840 3612 18846 3624
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 12526 3584 12532 3596
rect 11103 3556 12532 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 17736 3556 19993 3584
rect 17736 3544 17742 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1596 3448 1624 3479
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2280 3488 3065 3516
rect 2280 3476 2286 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4856 3488 4905 3516
rect 4856 3476 4862 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6696 3488 6929 3516
rect 6696 3476 6702 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 7892 3488 8401 3516
rect 7892 3476 7898 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9640 3488 9873 3516
rect 9640 3476 9646 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 10686 3516 10692 3528
rect 10643 3488 10692 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 12158 3516 12164 3528
rect 11379 3488 12164 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 16390 3516 16396 3528
rect 16347 3488 16396 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 19702 3516 19708 3528
rect 19659 3488 19708 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20772 3488 21281 3516
rect 20772 3476 20778 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 3602 3448 3608 3460
rect 1596 3420 3608 3448
rect 3602 3408 3608 3420
rect 3660 3408 3666 3460
rect 10042 3448 10048 3460
rect 3712 3420 10048 3448
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3712 3380 3740 3420
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 18693 3451 18751 3457
rect 18693 3448 18705 3451
rect 14608 3420 18705 3448
rect 14608 3408 14614 3420
rect 18693 3417 18705 3420
rect 18739 3417 18751 3451
rect 18693 3411 18751 3417
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 21744 3448 21772 3547
rect 23474 3544 23480 3596
rect 23532 3544 23538 3596
rect 23198 3476 23204 3528
rect 23256 3476 23262 3528
rect 24670 3476 24676 3528
rect 24728 3476 24734 3528
rect 19208 3420 21772 3448
rect 19208 3408 19214 3420
rect 24854 3408 24860 3460
rect 24912 3408 24918 3460
rect 3292 3352 3740 3380
rect 3292 3340 3298 3352
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 13722 3380 13728 3392
rect 9180 3352 13728 3380
rect 9180 3340 9186 3352
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 21082 3380 21088 3392
rect 19576 3352 21088 3380
rect 19576 3340 19582 3352
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9674 3176 9680 3188
rect 8435 3148 9680 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 7116 3108 7144 3139
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10962 3136 10968 3188
rect 11020 3136 11026 3188
rect 12618 3176 12624 3188
rect 11072 3148 12624 3176
rect 11072 3108 11100 3148
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16080 3148 20208 3176
rect 16080 3136 16086 3148
rect 14366 3108 14372 3120
rect 7116 3080 11100 3108
rect 12406 3080 14372 3108
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 2590 3040 2596 3052
rect 2179 3012 2596 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 3743 3012 6960 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 3234 2972 3240 2984
rect 2455 2944 3240 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3384 2944 3433 2972
rect 3384 2932 3390 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 5316 2944 5457 2972
rect 5316 2932 5322 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 6932 2972 6960 3012
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7064 3012 7297 3040
rect 7064 3000 7070 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8478 3040 8484 3052
rect 7975 3012 8484 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8846 3040 8852 3052
rect 8619 3012 8852 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 9214 3000 9220 3052
rect 9272 3000 9278 3052
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10318 3040 10324 3052
rect 9907 3012 10324 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 11054 3040 11060 3052
rect 10551 3012 11060 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11790 3040 11796 3052
rect 11195 3012 11796 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12406 3040 12434 3080
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 20180 3108 20208 3148
rect 20254 3136 20260 3188
rect 20312 3176 20318 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 20312 3148 20637 3176
rect 20312 3136 20318 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 20625 3139 20683 3145
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 23198 3176 23204 3188
rect 21315 3148 23204 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 23658 3136 23664 3188
rect 23716 3176 23722 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 23716 3148 24869 3176
rect 23716 3136 23722 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 16632 3080 19196 3108
rect 20180 3080 21496 3108
rect 16632 3068 16638 3080
rect 12023 3012 12434 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14148 3012 14841 3040
rect 14148 3000 14154 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 18414 3040 18420 3052
rect 17083 3012 18420 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 18564 3012 18705 3040
rect 18564 3000 18570 3012
rect 18693 3009 18705 3012
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 10134 2972 10140 2984
rect 6932 2944 10140 2972
rect 5445 2935 5503 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10336 2944 11376 2972
rect 10336 2913 10364 2944
rect 7745 2907 7803 2913
rect 7745 2873 7757 2907
rect 7791 2904 7803 2907
rect 10321 2907 10379 2913
rect 7791 2876 10088 2904
rect 7791 2873 7803 2876
rect 7745 2867 7803 2873
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 9122 2836 9128 2848
rect 9079 2808 9128 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9677 2839 9735 2845
rect 9677 2805 9689 2839
rect 9723 2836 9735 2839
rect 9766 2836 9772 2848
rect 9723 2808 9772 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10060 2836 10088 2876
rect 10321 2873 10333 2907
rect 10367 2873 10379 2907
rect 11348 2904 11376 2944
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11480 2944 11713 2972
rect 11480 2932 11486 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 19168 2981 19196 3080
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 21468 3049 21496 3080
rect 22002 3068 22008 3120
rect 22060 3108 22066 3120
rect 22097 3111 22155 3117
rect 22097 3108 22109 3111
rect 22060 3080 22109 3108
rect 22060 3068 22066 3080
rect 22097 3077 22109 3080
rect 22143 3077 22155 3111
rect 22097 3071 22155 3077
rect 22278 3068 22284 3120
rect 22336 3068 22342 3120
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20772 3012 20821 3040
rect 20772 3000 20778 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22462 3000 22468 3052
rect 22520 3040 22526 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22520 3012 22937 3040
rect 22520 3000 22526 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 23569 3043 23627 3049
rect 23569 3009 23581 3043
rect 23615 3040 23627 3043
rect 24302 3040 24308 3052
rect 23615 3012 24308 3040
rect 23615 3009 23627 3012
rect 23569 3003 23627 3009
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 16850 2904 16856 2916
rect 11348 2876 16856 2904
rect 10321 2867 10379 2873
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 16942 2864 16948 2916
rect 17000 2904 17006 2916
rect 19886 2904 19892 2916
rect 17000 2876 19892 2904
rect 17000 2864 17006 2876
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 21266 2904 21272 2916
rect 20680 2876 21272 2904
rect 20680 2864 20686 2876
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 21358 2864 21364 2916
rect 21416 2904 21422 2916
rect 22186 2904 22192 2916
rect 21416 2876 22192 2904
rect 21416 2864 21422 2876
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 22646 2904 22652 2916
rect 22336 2876 22652 2904
rect 22336 2864 22342 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 22738 2864 22744 2916
rect 22796 2864 22802 2916
rect 12710 2836 12716 2848
rect 10060 2808 12716 2836
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 17310 2836 17316 2848
rect 15160 2808 17316 2836
rect 15160 2796 15166 2808
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 22094 2836 22100 2848
rect 18472 2808 22100 2836
rect 18472 2796 18478 2808
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 2823 2635 2881 2641
rect 2823 2601 2835 2635
rect 2869 2632 2881 2635
rect 7101 2635 7159 2641
rect 2869 2604 6914 2632
rect 2869 2601 2881 2604
rect 2823 2595 2881 2601
rect 6886 2564 6914 2604
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 9030 2632 9036 2644
rect 7147 2604 9036 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 11701 2635 11759 2641
rect 9171 2604 10732 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 10226 2564 10232 2576
rect 6886 2536 10232 2564
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10704 2564 10732 2604
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 17126 2632 17132 2644
rect 11747 2604 17132 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 18690 2592 18696 2644
rect 18748 2592 18754 2644
rect 20898 2592 20904 2644
rect 20956 2632 20962 2644
rect 21453 2635 21511 2641
rect 21453 2632 21465 2635
rect 20956 2604 21465 2632
rect 20956 2592 20962 2604
rect 21453 2601 21465 2604
rect 21499 2601 21511 2635
rect 21453 2595 21511 2601
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 23198 2632 23204 2644
rect 21692 2604 23204 2632
rect 21692 2592 21698 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 24765 2635 24823 2641
rect 24765 2601 24777 2635
rect 24811 2632 24823 2635
rect 24946 2632 24952 2644
rect 24811 2604 24952 2632
rect 24811 2601 24823 2604
rect 24765 2595 24823 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 12342 2564 12348 2576
rect 10704 2536 12348 2564
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 16540 2536 22048 2564
rect 16540 2524 16546 2536
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 2958 2496 2964 2508
rect 2639 2468 2964 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5534 2496 5540 2508
rect 5215 2468 5540 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7708 2468 8033 2496
rect 7708 2456 7714 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 17310 2456 17316 2508
rect 17368 2456 17374 2508
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4724 2360 4752 2391
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7374 2428 7380 2440
rect 7331 2400 7380 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 6270 2360 6276 2372
rect 4724 2332 6276 2360
rect 6270 2320 6276 2332
rect 6328 2320 6334 2372
rect 9324 2360 9352 2391
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12158 2428 12164 2440
rect 11931 2400 12164 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12894 2428 12900 2440
rect 12575 2400 12900 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14240 2400 14473 2428
rect 14240 2388 14246 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 16853 2391 16911 2397
rect 17512 2400 18889 2428
rect 9950 2360 9956 2372
rect 9324 2332 9956 2360
rect 9950 2320 9956 2332
rect 10008 2320 10014 2372
rect 10962 2320 10968 2372
rect 11020 2320 11026 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 17512 2360 17540 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 22020 2437 22048 2536
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22152 2468 22477 2496
rect 22152 2456 22158 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19116 2400 19441 2428
rect 19116 2388 19122 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23808 2400 24041 2428
rect 23808 2388 23814 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 14332 2332 17540 2360
rect 18616 2332 18920 2360
rect 14332 2320 14338 2332
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2292 4583 2295
rect 10502 2292 10508 2304
rect 4571 2264 10508 2292
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 18616 2292 18644 2332
rect 13504 2264 18644 2292
rect 18892 2292 18920 2332
rect 19610 2320 19616 2372
rect 19668 2360 19674 2372
rect 22830 2360 22836 2372
rect 19668 2332 22836 2360
rect 19668 2320 19674 2332
rect 22830 2320 22836 2332
rect 22888 2320 22894 2372
rect 23845 2295 23903 2301
rect 23845 2292 23857 2295
rect 18892 2264 23857 2292
rect 13504 2252 13510 2264
rect 23845 2261 23857 2264
rect 23891 2261 23903 2295
rect 23845 2255 23903 2261
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 9858 1980 9864 2032
rect 9916 2020 9922 2032
rect 24854 2020 24860 2032
rect 9916 1992 24860 2020
rect 9916 1980 9922 1992
rect 24854 1980 24860 1992
rect 24912 1980 24918 2032
rect 10962 1912 10968 1964
rect 11020 1952 11026 1964
rect 22094 1952 22100 1964
rect 11020 1924 22100 1952
rect 11020 1912 11026 1924
rect 22094 1912 22100 1924
rect 22152 1912 22158 1964
rect 3418 1844 3424 1896
rect 3476 1884 3482 1896
rect 8754 1884 8760 1896
rect 3476 1856 8760 1884
rect 3476 1844 3482 1856
rect 8754 1844 8760 1856
rect 8812 1844 8818 1896
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 18604 54272 18656 54324
rect 8576 54204 8628 54256
rect 4068 54136 4120 54188
rect 4804 54179 4856 54188
rect 4804 54145 4813 54179
rect 4813 54145 4847 54179
rect 4847 54145 4856 54179
rect 4804 54136 4856 54145
rect 7380 54179 7432 54188
rect 7380 54145 7389 54179
rect 7389 54145 7423 54179
rect 7423 54145 7432 54179
rect 7380 54136 7432 54145
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 11704 54136 11756 54188
rect 13728 54136 13780 54188
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 18972 54136 19024 54188
rect 20628 54136 20680 54188
rect 21732 54136 21784 54188
rect 23112 54136 23164 54188
rect 24492 54136 24544 54188
rect 2412 54068 2464 54120
rect 5172 54111 5224 54120
rect 5172 54077 5181 54111
rect 5181 54077 5215 54111
rect 5215 54077 5224 54111
rect 5172 54068 5224 54077
rect 7840 54111 7892 54120
rect 7840 54077 7849 54111
rect 7849 54077 7883 54111
rect 7883 54077 7892 54111
rect 7840 54068 7892 54077
rect 9312 54068 9364 54120
rect 12348 54068 12400 54120
rect 15844 54000 15896 54052
rect 12440 53932 12492 53984
rect 14924 53975 14976 53984
rect 14924 53941 14933 53975
rect 14933 53941 14967 53975
rect 14967 53941 14976 53975
rect 14924 53932 14976 53941
rect 16120 53932 16172 53984
rect 17684 53975 17736 53984
rect 17684 53941 17693 53975
rect 17693 53941 17727 53975
rect 17727 53941 17736 53975
rect 17684 53932 17736 53941
rect 20904 53975 20956 53984
rect 20904 53941 20913 53975
rect 20913 53941 20947 53975
rect 20947 53941 20956 53975
rect 20904 53932 20956 53941
rect 24676 53932 24728 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 10692 53660 10744 53712
rect 1032 53592 1084 53644
rect 3792 53592 3844 53644
rect 6552 53592 6604 53644
rect 6644 53524 6696 53576
rect 7840 53524 7892 53576
rect 10692 53524 10744 53576
rect 23296 53524 23348 53576
rect 23756 53567 23808 53576
rect 23756 53533 23765 53567
rect 23765 53533 23799 53567
rect 23799 53533 23808 53567
rect 23756 53524 23808 53533
rect 25044 53567 25096 53576
rect 25044 53533 25053 53567
rect 25053 53533 25087 53567
rect 25087 53533 25096 53567
rect 25044 53524 25096 53533
rect 5540 53456 5592 53508
rect 22100 53388 22152 53440
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 26516 53388 26568 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 4068 53184 4120 53236
rect 7748 53048 7800 53100
rect 23388 53048 23440 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 19984 52844 20036 52896
rect 25780 52844 25832 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 25964 52436 26016 52488
rect 24952 52411 25004 52420
rect 24952 52377 24961 52411
rect 24961 52377 24995 52411
rect 24995 52377 25004 52411
rect 24952 52368 25004 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 6644 52139 6696 52148
rect 6644 52105 6653 52139
rect 6653 52105 6687 52139
rect 6687 52105 6696 52139
rect 6644 52096 6696 52105
rect 9404 51960 9456 52012
rect 25872 51960 25924 52012
rect 24124 51756 24176 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 7380 51552 7432 51604
rect 7840 51484 7892 51536
rect 4804 51348 4856 51400
rect 8484 51391 8536 51400
rect 8484 51357 8493 51391
rect 8493 51357 8527 51391
rect 8527 51357 8536 51391
rect 8484 51348 8536 51357
rect 10508 51348 10560 51400
rect 10600 51280 10652 51332
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 25044 51255 25096 51264
rect 25044 51221 25053 51255
rect 25053 51221 25087 51255
rect 25087 51221 25096 51255
rect 25044 51212 25096 51221
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 24952 50915 25004 50924
rect 24952 50881 24961 50915
rect 24961 50881 24995 50915
rect 24995 50881 25004 50915
rect 24952 50872 25004 50881
rect 17592 50668 17644 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 8392 50464 8444 50516
rect 9588 50507 9640 50516
rect 9588 50473 9597 50507
rect 9597 50473 9631 50507
rect 9631 50473 9640 50507
rect 9588 50464 9640 50473
rect 7748 50396 7800 50448
rect 8300 50396 8352 50448
rect 8576 50260 8628 50312
rect 9588 50260 9640 50312
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 24860 49784 24912 49836
rect 19800 49716 19852 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 10692 49351 10744 49360
rect 10692 49317 10701 49351
rect 10701 49317 10735 49351
rect 10735 49317 10744 49351
rect 10692 49308 10744 49317
rect 11704 49351 11756 49360
rect 11704 49317 11713 49351
rect 11713 49317 11747 49351
rect 11747 49317 11756 49351
rect 11704 49308 11756 49317
rect 10140 49104 10192 49156
rect 10876 49104 10928 49156
rect 25136 49147 25188 49156
rect 25136 49113 25145 49147
rect 25145 49113 25179 49147
rect 25179 49113 25188 49147
rect 25136 49104 25188 49113
rect 25228 49079 25280 49088
rect 25228 49045 25237 49079
rect 25237 49045 25271 49079
rect 25271 49045 25280 49079
rect 25228 49036 25280 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 8392 48875 8444 48884
rect 8392 48841 8401 48875
rect 8401 48841 8435 48875
rect 8435 48841 8444 48875
rect 8392 48832 8444 48841
rect 9956 48764 10008 48816
rect 9496 48628 9548 48680
rect 9128 48560 9180 48612
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 8300 48084 8352 48136
rect 25136 48059 25188 48068
rect 25136 48025 25145 48059
rect 25145 48025 25179 48059
rect 25179 48025 25188 48059
rect 25136 48016 25188 48025
rect 12348 47948 12400 48000
rect 21456 47948 21508 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9220 47744 9272 47796
rect 9404 47744 9456 47796
rect 8576 47608 8628 47660
rect 10232 47608 10284 47660
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 15936 47540 15988 47592
rect 22100 47540 22152 47592
rect 9496 47447 9548 47456
rect 9496 47413 9505 47447
rect 9505 47413 9539 47447
rect 9539 47413 9548 47447
rect 9496 47404 9548 47413
rect 25412 47404 25464 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 14924 47064 14976 47116
rect 9220 46996 9272 47048
rect 21088 46928 21140 46980
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 9772 46656 9824 46708
rect 10600 46656 10652 46708
rect 12348 46631 12400 46640
rect 12348 46597 12357 46631
rect 12357 46597 12391 46631
rect 12391 46597 12400 46631
rect 12348 46588 12400 46597
rect 8300 46563 8352 46572
rect 8300 46529 8309 46563
rect 8309 46529 8343 46563
rect 8343 46529 8352 46563
rect 8300 46520 8352 46529
rect 10232 46563 10284 46572
rect 10232 46529 10241 46563
rect 10241 46529 10275 46563
rect 10275 46529 10284 46563
rect 10232 46520 10284 46529
rect 16120 46588 16172 46640
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 7840 46452 7892 46504
rect 12440 46452 12492 46504
rect 13728 46495 13780 46504
rect 13728 46461 13737 46495
rect 13737 46461 13771 46495
rect 13771 46461 13780 46495
rect 13728 46452 13780 46461
rect 14648 46495 14700 46504
rect 14648 46461 14657 46495
rect 14657 46461 14691 46495
rect 14691 46461 14700 46495
rect 14648 46452 14700 46461
rect 16396 46452 16448 46504
rect 8484 46427 8536 46436
rect 8484 46393 8493 46427
rect 8493 46393 8527 46427
rect 8527 46393 8536 46427
rect 8484 46384 8536 46393
rect 10416 46359 10468 46368
rect 10416 46325 10425 46359
rect 10425 46325 10459 46359
rect 10459 46325 10468 46359
rect 10416 46316 10468 46325
rect 26056 46316 26108 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 14648 46112 14700 46164
rect 17684 45976 17736 46028
rect 10600 45908 10652 45960
rect 12808 45908 12860 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 17500 45883 17552 45892
rect 17500 45849 17509 45883
rect 17509 45849 17543 45883
rect 17543 45849 17552 45883
rect 17500 45840 17552 45849
rect 25780 45772 25832 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 10508 45500 10560 45552
rect 12808 45500 12860 45552
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 9404 45024 9456 45076
rect 9128 44931 9180 44940
rect 9128 44897 9137 44931
rect 9137 44897 9171 44931
rect 9171 44897 9180 44931
rect 9128 44888 9180 44897
rect 9404 44888 9456 44940
rect 9956 44888 10008 44940
rect 9680 44752 9732 44804
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 10784 44752 10836 44804
rect 10416 44684 10468 44736
rect 24952 44684 25004 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 9220 44344 9272 44396
rect 10232 44344 10284 44396
rect 24768 44344 24820 44396
rect 8944 44319 8996 44328
rect 8944 44285 8953 44319
rect 8953 44285 8987 44319
rect 8987 44285 8996 44319
rect 8944 44276 8996 44285
rect 10508 44208 10560 44260
rect 17684 44208 17736 44260
rect 25228 44208 25280 44260
rect 25504 44208 25556 44260
rect 10692 44183 10744 44192
rect 10692 44149 10701 44183
rect 10701 44149 10735 44183
rect 10735 44149 10744 44183
rect 10692 44140 10744 44149
rect 10968 44140 11020 44192
rect 17224 44140 17276 44192
rect 23940 44140 23992 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 24124 43800 24176 43852
rect 19524 43732 19576 43784
rect 20812 43664 20864 43716
rect 22192 43639 22244 43648
rect 22192 43605 22201 43639
rect 22201 43605 22235 43639
rect 22235 43605 22244 43639
rect 22192 43596 22244 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25136 43299 25188 43308
rect 25136 43265 25145 43299
rect 25145 43265 25179 43299
rect 25179 43265 25188 43299
rect 25136 43256 25188 43265
rect 25228 43095 25280 43104
rect 25228 43061 25237 43095
rect 25237 43061 25271 43095
rect 25271 43061 25280 43095
rect 25228 43052 25280 43061
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 9772 42755 9824 42764
rect 9772 42721 9781 42755
rect 9781 42721 9815 42755
rect 9815 42721 9824 42755
rect 9772 42712 9824 42721
rect 10140 42712 10192 42764
rect 8852 42644 8904 42696
rect 25136 42619 25188 42628
rect 25136 42585 25145 42619
rect 25145 42585 25179 42619
rect 25179 42585 25188 42619
rect 25136 42576 25188 42585
rect 26700 42576 26752 42628
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 9680 42304 9732 42356
rect 10784 42168 10836 42220
rect 9404 42143 9456 42152
rect 9404 42109 9413 42143
rect 9413 42109 9447 42143
rect 9447 42109 9456 42143
rect 9404 42100 9456 42109
rect 9680 42143 9732 42152
rect 9680 42109 9689 42143
rect 9689 42109 9723 42143
rect 9723 42109 9732 42143
rect 9680 42100 9732 42109
rect 10692 42100 10744 42152
rect 16304 42032 16356 42084
rect 19984 42032 20036 42084
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 10876 41760 10928 41812
rect 10968 41624 11020 41676
rect 9220 41556 9272 41608
rect 25136 41531 25188 41540
rect 25136 41497 25145 41531
rect 25145 41497 25179 41531
rect 25179 41497 25188 41531
rect 25136 41488 25188 41497
rect 25228 41463 25280 41472
rect 25228 41429 25237 41463
rect 25237 41429 25271 41463
rect 25271 41429 25280 41463
rect 25228 41420 25280 41429
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 26424 40876 26476 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 22836 40128 22888 40180
rect 25320 40035 25372 40044
rect 25320 40001 25329 40035
rect 25329 40001 25363 40035
rect 25363 40001 25372 40035
rect 25320 39992 25372 40001
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 23756 39244 23808 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 24860 38292 24912 38344
rect 25228 38292 25280 38344
rect 25320 38335 25372 38344
rect 25320 38301 25329 38335
rect 25329 38301 25363 38335
rect 25363 38301 25372 38335
rect 25320 38292 25372 38301
rect 24860 38156 24912 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 7840 37952 7892 38004
rect 9496 37816 9548 37868
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 25596 37680 25648 37732
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 15660 37272 15712 37324
rect 18604 37272 18656 37324
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 25228 36320 25280 36372
rect 25964 36252 26016 36304
rect 26056 36252 26108 36304
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 25228 35980 25280 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 9680 35776 9732 35828
rect 20260 35776 20312 35828
rect 25688 35776 25740 35828
rect 21088 35751 21140 35760
rect 21088 35717 21097 35751
rect 21097 35717 21131 35751
rect 21131 35717 21140 35751
rect 21088 35708 21140 35717
rect 26332 35708 26384 35760
rect 10784 35640 10836 35692
rect 16396 35640 16448 35692
rect 22744 35640 22796 35692
rect 9404 35615 9456 35624
rect 9404 35581 9413 35615
rect 9413 35581 9447 35615
rect 9447 35581 9456 35615
rect 9404 35572 9456 35581
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 21180 35572 21232 35624
rect 22652 35615 22704 35624
rect 22652 35581 22661 35615
rect 22661 35581 22695 35615
rect 22695 35581 22704 35615
rect 22652 35572 22704 35581
rect 19892 35436 19944 35488
rect 21088 35436 21140 35488
rect 23388 35436 23440 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 23296 35139 23348 35148
rect 23296 35105 23305 35139
rect 23305 35105 23339 35139
rect 23339 35105 23348 35139
rect 23296 35096 23348 35105
rect 17500 35028 17552 35080
rect 20536 35028 20588 35080
rect 24952 35028 25004 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 22468 34892 22520 34944
rect 25688 34892 25740 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 23480 34688 23532 34740
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 8944 34144 8996 34196
rect 21732 34144 21784 34196
rect 9404 34008 9456 34060
rect 19708 34008 19760 34060
rect 22284 34008 22336 34060
rect 9036 33940 9088 33992
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 20812 33940 20864 33992
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 14648 33915 14700 33924
rect 14648 33881 14657 33915
rect 14657 33881 14691 33915
rect 14691 33881 14700 33915
rect 14648 33872 14700 33881
rect 19984 33872 20036 33924
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 22928 33872 22980 33924
rect 22560 33804 22612 33856
rect 23204 33804 23256 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 22652 33600 22704 33652
rect 23204 33600 23256 33652
rect 20812 33532 20864 33584
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 22284 33532 22336 33584
rect 22928 33532 22980 33584
rect 25412 33464 25464 33516
rect 22376 33396 22428 33448
rect 22652 33396 22704 33448
rect 19984 33260 20036 33312
rect 20444 33260 20496 33312
rect 22928 33260 22980 33312
rect 23664 33260 23716 33312
rect 25872 33260 25924 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 16672 33056 16724 33108
rect 20904 33056 20956 33108
rect 22376 33056 22428 33108
rect 23296 33056 23348 33108
rect 25228 33056 25280 33108
rect 25688 33056 25740 33108
rect 23572 32988 23624 33040
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 23848 32920 23900 32972
rect 24768 32920 24820 32972
rect 26424 32988 26476 33040
rect 25136 32963 25188 32972
rect 25136 32929 25145 32963
rect 25145 32929 25179 32963
rect 25179 32929 25188 32963
rect 25136 32920 25188 32929
rect 19432 32852 19484 32904
rect 23664 32852 23716 32904
rect 14648 32784 14700 32836
rect 20352 32784 20404 32836
rect 25228 32784 25280 32836
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 14280 32444 14332 32496
rect 14648 32444 14700 32496
rect 18328 32444 18380 32496
rect 21180 32512 21232 32564
rect 20812 32444 20864 32496
rect 22284 32444 22336 32496
rect 19432 32376 19484 32428
rect 23664 32444 23716 32496
rect 24492 32512 24544 32564
rect 24768 32512 24820 32564
rect 12808 32308 12860 32360
rect 16764 32308 16816 32360
rect 18236 32308 18288 32360
rect 20352 32308 20404 32360
rect 25136 32308 25188 32360
rect 19064 32215 19116 32224
rect 19064 32181 19073 32215
rect 19073 32181 19107 32215
rect 19107 32181 19116 32215
rect 19064 32172 19116 32181
rect 20812 32172 20864 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 18236 31968 18288 32020
rect 18604 31968 18656 32020
rect 19708 31968 19760 32020
rect 14096 31900 14148 31952
rect 19064 31900 19116 31952
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 16764 31875 16816 31884
rect 16764 31841 16773 31875
rect 16773 31841 16807 31875
rect 16807 31841 16816 31875
rect 16764 31832 16816 31841
rect 18420 31832 18472 31884
rect 19432 31875 19484 31884
rect 19432 31841 19441 31875
rect 19441 31841 19475 31875
rect 19475 31841 19484 31875
rect 19432 31832 19484 31841
rect 16672 31764 16724 31816
rect 23756 31968 23808 32020
rect 23388 31900 23440 31952
rect 25044 31900 25096 31952
rect 22560 31832 22612 31884
rect 22652 31832 22704 31884
rect 22836 31764 22888 31816
rect 22928 31764 22980 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 18328 31696 18380 31748
rect 21088 31696 21140 31748
rect 21272 31696 21324 31748
rect 22744 31696 22796 31748
rect 17132 31628 17184 31680
rect 20996 31628 21048 31680
rect 22376 31628 22428 31680
rect 23296 31628 23348 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 24860 31424 24912 31476
rect 14924 31356 14976 31408
rect 16120 31356 16172 31408
rect 15844 31288 15896 31340
rect 16028 31331 16080 31340
rect 16028 31297 16037 31331
rect 16037 31297 16071 31331
rect 16071 31297 16080 31331
rect 16028 31288 16080 31297
rect 17224 31331 17276 31340
rect 17224 31297 17233 31331
rect 17233 31297 17267 31331
rect 17267 31297 17276 31331
rect 17224 31288 17276 31297
rect 20536 31399 20588 31408
rect 20536 31365 20545 31399
rect 20545 31365 20579 31399
rect 20579 31365 20588 31399
rect 20536 31356 20588 31365
rect 22100 31356 22152 31408
rect 22652 31399 22704 31408
rect 22652 31365 22661 31399
rect 22661 31365 22695 31399
rect 22695 31365 22704 31399
rect 22652 31356 22704 31365
rect 24492 31356 24544 31408
rect 12808 31220 12860 31272
rect 16212 31263 16264 31272
rect 16212 31229 16221 31263
rect 16221 31229 16255 31263
rect 16255 31229 16264 31263
rect 16212 31220 16264 31229
rect 17316 31263 17368 31272
rect 17316 31229 17325 31263
rect 17325 31229 17359 31263
rect 17359 31229 17368 31263
rect 17316 31220 17368 31229
rect 22192 31288 22244 31340
rect 22284 31288 22336 31340
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 18420 31220 18472 31272
rect 18696 31220 18748 31272
rect 14556 31152 14608 31204
rect 17132 31152 17184 31204
rect 24676 31220 24728 31272
rect 15016 31127 15068 31136
rect 15016 31093 15025 31127
rect 15025 31093 15059 31127
rect 15059 31093 15068 31127
rect 15016 31084 15068 31093
rect 15936 31084 15988 31136
rect 18512 31084 18564 31136
rect 23664 31084 23716 31136
rect 24952 31084 25004 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 9220 30880 9272 30932
rect 17408 30880 17460 30932
rect 18696 30880 18748 30932
rect 22652 30880 22704 30932
rect 26240 30812 26292 30864
rect 19432 30744 19484 30796
rect 20996 30744 21048 30796
rect 26516 30744 26568 30796
rect 8760 30676 8812 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 20168 30719 20220 30728
rect 20168 30685 20177 30719
rect 20177 30685 20211 30719
rect 20211 30685 20220 30719
rect 20168 30676 20220 30685
rect 25412 30676 25464 30728
rect 13912 30608 13964 30660
rect 18328 30608 18380 30660
rect 18696 30608 18748 30660
rect 20904 30651 20956 30660
rect 20904 30617 20913 30651
rect 20913 30617 20947 30651
rect 20947 30617 20956 30651
rect 20904 30608 20956 30617
rect 18788 30540 18840 30592
rect 21272 30540 21324 30592
rect 22744 30540 22796 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 12808 30336 12860 30388
rect 16028 30336 16080 30388
rect 20996 30336 21048 30388
rect 7656 30200 7708 30252
rect 14280 30311 14332 30320
rect 14280 30277 14289 30311
rect 14289 30277 14323 30311
rect 14323 30277 14332 30311
rect 14280 30268 14332 30277
rect 20168 30311 20220 30320
rect 20168 30277 20177 30311
rect 20177 30277 20211 30311
rect 20211 30277 20220 30311
rect 20168 30268 20220 30277
rect 20260 30311 20312 30320
rect 20260 30277 20269 30311
rect 20269 30277 20303 30311
rect 20303 30277 20312 30311
rect 20260 30268 20312 30277
rect 22468 30311 22520 30320
rect 22468 30277 22477 30311
rect 22477 30277 22511 30311
rect 22511 30277 22520 30311
rect 22468 30268 22520 30277
rect 24584 30268 24636 30320
rect 12716 30132 12768 30184
rect 8852 30107 8904 30116
rect 8852 30073 8861 30107
rect 8861 30073 8895 30107
rect 8895 30073 8904 30107
rect 8852 30064 8904 30073
rect 10784 29996 10836 30048
rect 12532 29996 12584 30048
rect 14924 30200 14976 30252
rect 13728 30132 13780 30184
rect 20628 30200 20680 30252
rect 15108 30175 15160 30184
rect 15108 30141 15117 30175
rect 15117 30141 15151 30175
rect 15151 30141 15160 30175
rect 15108 30132 15160 30141
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 22836 30132 22888 30184
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 23664 30132 23716 30184
rect 25136 30132 25188 30184
rect 15568 30064 15620 30116
rect 13452 30039 13504 30048
rect 13452 30005 13461 30039
rect 13461 30005 13495 30039
rect 13495 30005 13504 30039
rect 13452 29996 13504 30005
rect 16120 29996 16172 30048
rect 19248 29996 19300 30048
rect 21916 29996 21968 30048
rect 25964 29996 26016 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 11612 29792 11664 29844
rect 13452 29792 13504 29844
rect 18788 29835 18840 29844
rect 18788 29801 18797 29835
rect 18797 29801 18831 29835
rect 18831 29801 18840 29835
rect 18788 29792 18840 29801
rect 12716 29724 12768 29776
rect 11428 29656 11480 29708
rect 13912 29656 13964 29708
rect 18328 29724 18380 29776
rect 16212 29656 16264 29708
rect 17868 29656 17920 29708
rect 12532 29588 12584 29640
rect 15568 29631 15620 29640
rect 15568 29597 15577 29631
rect 15577 29597 15611 29631
rect 15611 29597 15620 29631
rect 15568 29588 15620 29597
rect 18696 29656 18748 29708
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 20812 29656 20864 29708
rect 11060 29520 11112 29572
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 15384 29452 15436 29504
rect 18880 29588 18932 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 20628 29520 20680 29572
rect 19432 29495 19484 29504
rect 19432 29461 19441 29495
rect 19441 29461 19475 29495
rect 19475 29461 19484 29495
rect 19432 29452 19484 29461
rect 19524 29452 19576 29504
rect 23480 29520 23532 29572
rect 23940 29452 23992 29504
rect 25136 29495 25188 29504
rect 25136 29461 25145 29495
rect 25145 29461 25179 29495
rect 25179 29461 25188 29495
rect 25136 29452 25188 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 9496 29291 9548 29300
rect 9496 29257 9505 29291
rect 9505 29257 9539 29291
rect 9539 29257 9548 29291
rect 9496 29248 9548 29257
rect 15200 29248 15252 29300
rect 16212 29248 16264 29300
rect 19432 29248 19484 29300
rect 19708 29291 19760 29300
rect 19708 29257 19717 29291
rect 19717 29257 19751 29291
rect 19751 29257 19760 29291
rect 19708 29248 19760 29257
rect 24860 29248 24912 29300
rect 10324 29180 10376 29232
rect 10232 29112 10284 29164
rect 13912 29180 13964 29232
rect 14924 29180 14976 29232
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 9680 29044 9732 29096
rect 10876 29044 10928 29096
rect 13636 29044 13688 29096
rect 16120 29087 16172 29096
rect 16120 29053 16129 29087
rect 16129 29053 16163 29087
rect 16163 29053 16172 29087
rect 16120 29044 16172 29053
rect 16672 29044 16724 29096
rect 14924 28976 14976 29028
rect 14188 28908 14240 28960
rect 15200 28976 15252 29028
rect 15752 28976 15804 29028
rect 17132 29044 17184 29096
rect 23940 29223 23992 29232
rect 23940 29189 23949 29223
rect 23949 29189 23983 29223
rect 23983 29189 23992 29223
rect 23940 29180 23992 29189
rect 25228 29180 25280 29232
rect 19524 29112 19576 29164
rect 19616 29155 19668 29164
rect 19616 29121 19625 29155
rect 19625 29121 19659 29155
rect 19659 29121 19668 29155
rect 19616 29112 19668 29121
rect 20352 29112 20404 29164
rect 23480 29112 23532 29164
rect 24584 29112 24636 29164
rect 24768 29112 24820 29164
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 20904 29044 20956 29096
rect 17776 28976 17828 29028
rect 19156 28976 19208 29028
rect 22192 28976 22244 29028
rect 23296 29044 23348 29096
rect 23756 29044 23808 29096
rect 24308 28976 24360 29028
rect 24860 28976 24912 29028
rect 18696 28908 18748 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 10876 28747 10928 28756
rect 10876 28713 10885 28747
rect 10885 28713 10919 28747
rect 10919 28713 10928 28747
rect 10876 28704 10928 28713
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 19616 28704 19668 28756
rect 21456 28704 21508 28756
rect 13820 28636 13872 28688
rect 10416 28568 10468 28620
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 12440 28568 12492 28620
rect 19064 28568 19116 28620
rect 19432 28568 19484 28620
rect 20536 28611 20588 28620
rect 20536 28577 20545 28611
rect 20545 28577 20579 28611
rect 20579 28577 20588 28611
rect 20536 28568 20588 28577
rect 20812 28611 20864 28620
rect 20812 28577 20821 28611
rect 20821 28577 20855 28611
rect 20855 28577 20864 28611
rect 20812 28568 20864 28577
rect 21272 28568 21324 28620
rect 23480 28636 23532 28688
rect 23572 28611 23624 28620
rect 23572 28577 23581 28611
rect 23581 28577 23615 28611
rect 23615 28577 23624 28611
rect 23572 28568 23624 28577
rect 23848 28568 23900 28620
rect 15108 28500 15160 28552
rect 9680 28432 9732 28484
rect 9956 28432 10008 28484
rect 11612 28432 11664 28484
rect 12716 28432 12768 28484
rect 18696 28432 18748 28484
rect 18880 28432 18932 28484
rect 20812 28432 20864 28484
rect 21272 28432 21324 28484
rect 14188 28364 14240 28416
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 14924 28364 14976 28416
rect 15660 28364 15712 28416
rect 15936 28364 15988 28416
rect 16304 28407 16356 28416
rect 16304 28373 16313 28407
rect 16313 28373 16347 28407
rect 16347 28373 16356 28407
rect 16304 28364 16356 28373
rect 16396 28407 16448 28416
rect 16396 28373 16405 28407
rect 16405 28373 16439 28407
rect 16439 28373 16448 28407
rect 26148 28432 26200 28484
rect 16396 28364 16448 28373
rect 23756 28364 23808 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 14096 28203 14148 28212
rect 14096 28169 14105 28203
rect 14105 28169 14139 28203
rect 14139 28169 14148 28203
rect 14096 28160 14148 28169
rect 18512 28203 18564 28212
rect 18512 28169 18521 28203
rect 18521 28169 18555 28203
rect 18555 28169 18564 28203
rect 18512 28160 18564 28169
rect 23296 28160 23348 28212
rect 14556 28092 14608 28144
rect 17684 28092 17736 28144
rect 20352 28135 20404 28144
rect 20352 28101 20361 28135
rect 20361 28101 20395 28135
rect 20395 28101 20404 28135
rect 20352 28092 20404 28101
rect 20536 28092 20588 28144
rect 16580 28024 16632 28076
rect 17224 28067 17276 28076
rect 17224 28033 17233 28067
rect 17233 28033 17267 28067
rect 17267 28033 17276 28067
rect 17224 28024 17276 28033
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 22192 28092 22244 28144
rect 23664 28092 23716 28144
rect 23388 28024 23440 28076
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 9404 27956 9456 28008
rect 15016 27956 15068 28008
rect 17316 27999 17368 28008
rect 17316 27965 17325 27999
rect 17325 27965 17359 27999
rect 17359 27965 17368 27999
rect 17316 27956 17368 27965
rect 17408 27999 17460 28008
rect 17408 27965 17417 27999
rect 17417 27965 17451 27999
rect 17451 27965 17460 27999
rect 17408 27956 17460 27965
rect 18604 27999 18656 28008
rect 18604 27965 18613 27999
rect 18613 27965 18647 27999
rect 18647 27965 18656 27999
rect 18604 27956 18656 27965
rect 22652 27956 22704 28008
rect 12164 27820 12216 27872
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 18788 27820 18840 27872
rect 22836 27820 22888 27872
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 18420 27616 18472 27668
rect 22836 27616 22888 27668
rect 24584 27616 24636 27668
rect 22100 27548 22152 27600
rect 9220 27480 9272 27532
rect 13084 27480 13136 27532
rect 13544 27523 13596 27532
rect 13544 27489 13553 27523
rect 13553 27489 13587 27523
rect 13587 27489 13596 27523
rect 13544 27480 13596 27489
rect 15016 27480 15068 27532
rect 14740 27412 14792 27464
rect 22836 27523 22888 27532
rect 22836 27489 22845 27523
rect 22845 27489 22879 27523
rect 22879 27489 22888 27523
rect 22836 27480 22888 27489
rect 22192 27412 22244 27464
rect 23296 27412 23348 27464
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 25228 27523 25280 27532
rect 25228 27489 25237 27523
rect 25237 27489 25271 27523
rect 25271 27489 25280 27523
rect 25228 27480 25280 27489
rect 10784 27387 10836 27396
rect 10784 27353 10793 27387
rect 10793 27353 10827 27387
rect 10827 27353 10836 27387
rect 10784 27344 10836 27353
rect 9956 27276 10008 27328
rect 13820 27344 13872 27396
rect 14280 27344 14332 27396
rect 14924 27344 14976 27396
rect 17500 27344 17552 27396
rect 20812 27344 20864 27396
rect 25872 27344 25924 27396
rect 12440 27276 12492 27328
rect 12532 27276 12584 27328
rect 15292 27276 15344 27328
rect 15936 27276 15988 27328
rect 19064 27276 19116 27328
rect 19708 27276 19760 27328
rect 20904 27276 20956 27328
rect 21824 27276 21876 27328
rect 22560 27319 22612 27328
rect 22560 27285 22569 27319
rect 22569 27285 22603 27319
rect 22603 27285 22612 27319
rect 22560 27276 22612 27285
rect 22836 27276 22888 27328
rect 23480 27276 23532 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 11060 27072 11112 27124
rect 13084 27072 13136 27124
rect 15108 27072 15160 27124
rect 16856 27072 16908 27124
rect 18880 27072 18932 27124
rect 9956 27004 10008 27056
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 12808 26936 12860 26988
rect 13636 27004 13688 27056
rect 13820 27004 13872 27056
rect 15752 27047 15804 27056
rect 15752 27013 15761 27047
rect 15761 27013 15795 27047
rect 15795 27013 15804 27047
rect 15752 27004 15804 27013
rect 19708 27115 19760 27124
rect 19708 27081 19717 27115
rect 19717 27081 19751 27115
rect 19751 27081 19760 27115
rect 19708 27072 19760 27081
rect 21732 27072 21784 27124
rect 20812 27004 20864 27056
rect 23572 27004 23624 27056
rect 24400 27072 24452 27124
rect 15108 26936 15160 26988
rect 16028 26936 16080 26988
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 21088 26979 21140 26988
rect 21088 26945 21097 26979
rect 21097 26945 21131 26979
rect 21131 26945 21140 26979
rect 21088 26936 21140 26945
rect 10048 26868 10100 26920
rect 10692 26800 10744 26852
rect 12440 26800 12492 26852
rect 11980 26732 12032 26784
rect 14924 26732 14976 26784
rect 18604 26732 18656 26784
rect 23296 26911 23348 26920
rect 23296 26877 23305 26911
rect 23305 26877 23339 26911
rect 23339 26877 23348 26911
rect 23296 26868 23348 26877
rect 25228 26868 25280 26920
rect 24584 26800 24636 26852
rect 25136 26800 25188 26852
rect 21180 26732 21232 26784
rect 22652 26732 22704 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 10048 26528 10100 26580
rect 13544 26528 13596 26580
rect 11796 26460 11848 26512
rect 10416 26435 10468 26444
rect 10416 26401 10425 26435
rect 10425 26401 10459 26435
rect 10459 26401 10468 26435
rect 10416 26392 10468 26401
rect 10692 26435 10744 26444
rect 10692 26401 10701 26435
rect 10701 26401 10735 26435
rect 10735 26401 10744 26435
rect 10692 26392 10744 26401
rect 12072 26392 12124 26444
rect 21088 26528 21140 26580
rect 21180 26571 21232 26580
rect 21180 26537 21189 26571
rect 21189 26537 21223 26571
rect 21223 26537 21232 26571
rect 21180 26528 21232 26537
rect 25044 26528 25096 26580
rect 14832 26435 14884 26444
rect 14832 26401 14841 26435
rect 14841 26401 14875 26435
rect 14875 26401 14884 26435
rect 14832 26392 14884 26401
rect 16396 26460 16448 26512
rect 14740 26324 14792 26376
rect 15016 26324 15068 26376
rect 17960 26392 18012 26444
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 20904 26392 20956 26444
rect 18420 26367 18472 26376
rect 18420 26333 18429 26367
rect 18429 26333 18463 26367
rect 18463 26333 18472 26367
rect 18420 26324 18472 26333
rect 20812 26324 20864 26376
rect 21640 26460 21692 26512
rect 22468 26460 22520 26512
rect 25412 26460 25464 26512
rect 22284 26392 22336 26444
rect 9864 26256 9916 26308
rect 15844 26256 15896 26308
rect 16856 26256 16908 26308
rect 22192 26367 22244 26376
rect 22192 26333 22201 26367
rect 22201 26333 22235 26367
rect 22235 26333 22244 26367
rect 22192 26324 22244 26333
rect 22376 26324 22428 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 24952 26392 25004 26444
rect 25136 26435 25188 26444
rect 25136 26401 25145 26435
rect 25145 26401 25179 26435
rect 25179 26401 25188 26435
rect 25136 26392 25188 26401
rect 22836 26256 22888 26308
rect 24584 26256 24636 26308
rect 12716 26188 12768 26240
rect 13820 26188 13872 26240
rect 15108 26188 15160 26240
rect 15568 26231 15620 26240
rect 15568 26197 15577 26231
rect 15577 26197 15611 26231
rect 15611 26197 15620 26231
rect 15568 26188 15620 26197
rect 16304 26188 16356 26240
rect 17224 26188 17276 26240
rect 25872 26256 25924 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 10784 25984 10836 26036
rect 8944 25916 8996 25968
rect 9404 25959 9456 25968
rect 9404 25925 9413 25959
rect 9413 25925 9447 25959
rect 9447 25925 9456 25959
rect 9404 25916 9456 25925
rect 9864 25916 9916 25968
rect 12532 26027 12584 26036
rect 12532 25993 12541 26027
rect 12541 25993 12575 26027
rect 12575 25993 12584 26027
rect 12532 25984 12584 25993
rect 15200 25984 15252 26036
rect 16764 25984 16816 26036
rect 17592 25984 17644 26036
rect 18420 25984 18472 26036
rect 22100 25984 22152 26036
rect 22376 26027 22428 26036
rect 22376 25993 22385 26027
rect 22385 25993 22419 26027
rect 22419 25993 22428 26027
rect 22376 25984 22428 25993
rect 22744 25984 22796 26036
rect 25228 25984 25280 26036
rect 9128 25891 9180 25900
rect 9128 25857 9137 25891
rect 9137 25857 9171 25891
rect 9171 25857 9180 25891
rect 9128 25848 9180 25857
rect 12440 25891 12492 25900
rect 12440 25857 12449 25891
rect 12449 25857 12483 25891
rect 12483 25857 12492 25891
rect 12440 25848 12492 25857
rect 11060 25780 11112 25832
rect 10968 25712 11020 25764
rect 13820 25848 13872 25900
rect 18328 25959 18380 25968
rect 18328 25925 18337 25959
rect 18337 25925 18371 25959
rect 18371 25925 18380 25959
rect 18328 25916 18380 25925
rect 24400 25916 24452 25968
rect 13636 25780 13688 25832
rect 14188 25823 14240 25832
rect 14188 25789 14197 25823
rect 14197 25789 14231 25823
rect 14231 25789 14240 25823
rect 14188 25780 14240 25789
rect 18696 25780 18748 25832
rect 22836 25780 22888 25832
rect 23296 25780 23348 25832
rect 23572 25823 23624 25832
rect 23572 25789 23581 25823
rect 23581 25789 23615 25823
rect 23615 25789 23624 25823
rect 23572 25780 23624 25789
rect 25228 25780 25280 25832
rect 20904 25712 20956 25764
rect 10416 25644 10468 25696
rect 13452 25644 13504 25696
rect 16764 25644 16816 25696
rect 16948 25644 17000 25696
rect 19892 25687 19944 25696
rect 19892 25653 19901 25687
rect 19901 25653 19935 25687
rect 19935 25653 19944 25687
rect 19892 25644 19944 25653
rect 20720 25644 20772 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 10324 25440 10376 25492
rect 11152 25440 11204 25492
rect 14832 25440 14884 25492
rect 13360 25372 13412 25424
rect 9680 25304 9732 25356
rect 12808 25304 12860 25356
rect 13452 25304 13504 25356
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 16764 25304 16816 25356
rect 10968 25279 11020 25288
rect 10968 25245 10977 25279
rect 10977 25245 11011 25279
rect 11011 25245 11020 25279
rect 10968 25236 11020 25245
rect 13728 25236 13780 25288
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 23940 25304 23992 25356
rect 10784 25168 10836 25220
rect 11980 25168 12032 25220
rect 12716 25168 12768 25220
rect 11704 25100 11756 25152
rect 14832 25168 14884 25220
rect 15476 25168 15528 25220
rect 16580 25168 16632 25220
rect 15200 25100 15252 25152
rect 15384 25100 15436 25152
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 15936 25100 15988 25152
rect 18512 25168 18564 25220
rect 19984 25211 20036 25220
rect 19984 25177 19993 25211
rect 19993 25177 20027 25211
rect 20027 25177 20036 25211
rect 19984 25168 20036 25177
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 19800 25100 19852 25152
rect 24952 25168 25004 25220
rect 21732 25100 21784 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 7472 24896 7524 24948
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 18696 24896 18748 24948
rect 9864 24828 9916 24880
rect 12716 24828 12768 24880
rect 15200 24828 15252 24880
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 12808 24760 12860 24812
rect 16580 24828 16632 24880
rect 20260 24828 20312 24880
rect 24124 24828 24176 24880
rect 24400 24828 24452 24880
rect 18512 24803 18564 24812
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 9312 24735 9364 24744
rect 9312 24701 9321 24735
rect 9321 24701 9355 24735
rect 9355 24701 9364 24735
rect 9312 24692 9364 24701
rect 9680 24692 9732 24744
rect 10876 24624 10928 24676
rect 13360 24692 13412 24744
rect 14832 24692 14884 24744
rect 18420 24692 18472 24744
rect 19432 24760 19484 24812
rect 21088 24760 21140 24812
rect 23480 24760 23532 24812
rect 17040 24624 17092 24676
rect 19616 24692 19668 24744
rect 20444 24692 20496 24744
rect 22284 24692 22336 24744
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 23296 24692 23348 24744
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 25136 24692 25188 24744
rect 25228 24692 25280 24744
rect 11152 24556 11204 24608
rect 13728 24556 13780 24608
rect 14740 24599 14792 24608
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 15476 24556 15528 24608
rect 17224 24556 17276 24608
rect 17776 24556 17828 24608
rect 17868 24556 17920 24608
rect 19708 24556 19760 24608
rect 20628 24556 20680 24608
rect 22192 24556 22244 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 14740 24352 14792 24404
rect 21088 24352 21140 24404
rect 23296 24284 23348 24336
rect 9312 24216 9364 24268
rect 12348 24216 12400 24268
rect 18604 24259 18656 24268
rect 18604 24225 18613 24259
rect 18613 24225 18647 24259
rect 18647 24225 18656 24259
rect 18604 24216 18656 24225
rect 19064 24216 19116 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 20444 24216 20496 24268
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 18880 24148 18932 24200
rect 21088 24148 21140 24200
rect 9864 24080 9916 24132
rect 9128 24012 9180 24064
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 18328 24012 18380 24064
rect 19984 24080 20036 24132
rect 22100 24080 22152 24132
rect 22284 24080 22336 24132
rect 24124 24352 24176 24404
rect 24952 24148 25004 24200
rect 25412 24148 25464 24200
rect 23572 24080 23624 24132
rect 24400 24080 24452 24132
rect 23480 24012 23532 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 8668 23740 8720 23792
rect 9128 23740 9180 23792
rect 9864 23808 9916 23860
rect 9496 23740 9548 23792
rect 12624 23740 12676 23792
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 15108 23808 15160 23860
rect 15568 23740 15620 23792
rect 15936 23740 15988 23792
rect 7840 23604 7892 23656
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 13912 23672 13964 23724
rect 13360 23536 13412 23588
rect 17224 23604 17276 23656
rect 19892 23808 19944 23860
rect 20904 23851 20956 23860
rect 20904 23817 20913 23851
rect 20913 23817 20947 23851
rect 20947 23817 20956 23851
rect 20904 23808 20956 23817
rect 21824 23808 21876 23860
rect 25136 23808 25188 23860
rect 19524 23740 19576 23792
rect 19800 23740 19852 23792
rect 9680 23468 9732 23520
rect 10508 23511 10560 23520
rect 10508 23477 10517 23511
rect 10517 23477 10551 23511
rect 10551 23477 10560 23511
rect 10508 23468 10560 23477
rect 12256 23468 12308 23520
rect 13728 23468 13780 23520
rect 15292 23468 15344 23520
rect 15844 23511 15896 23520
rect 15844 23477 15853 23511
rect 15853 23477 15887 23511
rect 15887 23477 15896 23511
rect 15844 23468 15896 23477
rect 16304 23468 16356 23520
rect 22008 23672 22060 23724
rect 24492 23740 24544 23792
rect 19432 23604 19484 23656
rect 19708 23604 19760 23656
rect 19984 23647 20036 23656
rect 19984 23613 19993 23647
rect 19993 23613 20027 23647
rect 20027 23613 20036 23647
rect 19984 23604 20036 23613
rect 20996 23604 21048 23656
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 23480 23647 23532 23656
rect 23480 23613 23489 23647
rect 23489 23613 23523 23647
rect 23523 23613 23532 23647
rect 23480 23604 23532 23613
rect 22836 23536 22888 23588
rect 19892 23468 19944 23520
rect 20536 23511 20588 23520
rect 20536 23477 20545 23511
rect 20545 23477 20579 23511
rect 20579 23477 20588 23511
rect 20536 23468 20588 23477
rect 22652 23468 22704 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 9036 23264 9088 23316
rect 14740 23307 14792 23316
rect 14740 23273 14749 23307
rect 14749 23273 14783 23307
rect 14783 23273 14792 23307
rect 14740 23264 14792 23273
rect 16396 23264 16448 23316
rect 17316 23264 17368 23316
rect 18236 23264 18288 23316
rect 18420 23264 18472 23316
rect 20812 23264 20864 23316
rect 20904 23307 20956 23316
rect 20904 23273 20913 23307
rect 20913 23273 20947 23307
rect 20947 23273 20956 23307
rect 20904 23264 20956 23273
rect 9220 23196 9272 23248
rect 8576 23128 8628 23180
rect 11060 23128 11112 23180
rect 13360 23196 13412 23248
rect 15108 23196 15160 23248
rect 16580 23196 16632 23248
rect 17592 23196 17644 23248
rect 21364 23196 21416 23248
rect 8392 23060 8444 23112
rect 9496 23060 9548 23112
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 12808 23060 12860 23112
rect 18236 23171 18288 23180
rect 18236 23137 18245 23171
rect 18245 23137 18279 23171
rect 18279 23137 18288 23171
rect 18236 23128 18288 23137
rect 18604 23128 18656 23180
rect 20444 23128 20496 23180
rect 23388 23128 23440 23180
rect 24860 23128 24912 23180
rect 25320 23128 25372 23180
rect 15844 23060 15896 23112
rect 8852 22992 8904 23044
rect 11796 22992 11848 23044
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 10324 22924 10376 22976
rect 12532 22924 12584 22976
rect 13360 22967 13412 22976
rect 13360 22933 13369 22967
rect 13369 22933 13403 22967
rect 13403 22933 13412 22967
rect 13360 22924 13412 22933
rect 17224 22992 17276 23044
rect 16580 22924 16632 22976
rect 18420 22992 18472 23044
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 20720 23060 20772 23112
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22652 23103 22704 23112
rect 22652 23069 22661 23103
rect 22661 23069 22695 23103
rect 22695 23069 22704 23103
rect 22652 23060 22704 23069
rect 25872 23060 25924 23112
rect 18696 22992 18748 23044
rect 20996 22992 21048 23044
rect 18512 22924 18564 22976
rect 22652 22924 22704 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 3424 22720 3476 22772
rect 12072 22720 12124 22772
rect 13452 22720 13504 22772
rect 21824 22720 21876 22772
rect 8392 22652 8444 22704
rect 12624 22695 12676 22704
rect 12624 22661 12633 22695
rect 12633 22661 12667 22695
rect 12667 22661 12676 22695
rect 12624 22652 12676 22661
rect 12716 22652 12768 22704
rect 17224 22652 17276 22704
rect 19892 22652 19944 22704
rect 21732 22652 21784 22704
rect 7840 22584 7892 22636
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 10968 22516 11020 22568
rect 12716 22516 12768 22568
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 22376 22652 22428 22704
rect 24860 22652 24912 22704
rect 21088 22584 21140 22593
rect 23756 22584 23808 22636
rect 23940 22627 23992 22636
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 10416 22448 10468 22500
rect 20076 22448 20128 22500
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 20168 22423 20220 22432
rect 20168 22389 20177 22423
rect 20177 22389 20211 22423
rect 20211 22389 20220 22423
rect 20168 22380 20220 22389
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 20812 22380 20864 22432
rect 21088 22380 21140 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 10508 22176 10560 22228
rect 10600 22108 10652 22160
rect 11612 22108 11664 22160
rect 12256 22040 12308 22092
rect 15752 22108 15804 22160
rect 22836 22108 22888 22160
rect 9864 21972 9916 22024
rect 10140 21972 10192 22024
rect 11060 21972 11112 22024
rect 13820 21972 13872 22024
rect 14096 21972 14148 22024
rect 17040 22040 17092 22092
rect 19616 22040 19668 22092
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 23204 22040 23256 22092
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 20260 21972 20312 22024
rect 22928 21972 22980 22024
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 25228 22108 25280 22160
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 12716 21904 12768 21956
rect 16580 21904 16632 21956
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 17132 21836 17184 21888
rect 20628 21904 20680 21956
rect 21824 21947 21876 21956
rect 21824 21913 21833 21947
rect 21833 21913 21867 21947
rect 21867 21913 21876 21947
rect 21824 21904 21876 21913
rect 22008 21836 22060 21888
rect 23388 21836 23440 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 7380 21632 7432 21684
rect 10140 21632 10192 21684
rect 10232 21632 10284 21684
rect 8392 21564 8444 21616
rect 7840 21496 7892 21548
rect 9312 21428 9364 21480
rect 12256 21632 12308 21684
rect 11612 21564 11664 21616
rect 11796 21564 11848 21616
rect 13452 21564 13504 21616
rect 11060 21496 11112 21548
rect 12348 21496 12400 21548
rect 12716 21496 12768 21548
rect 14832 21564 14884 21616
rect 20168 21632 20220 21684
rect 21824 21632 21876 21684
rect 22836 21632 22888 21684
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 14096 21428 14148 21480
rect 12164 21360 12216 21412
rect 11152 21292 11204 21344
rect 13360 21292 13412 21344
rect 14924 21428 14976 21480
rect 16212 21496 16264 21548
rect 22560 21564 22612 21616
rect 19432 21496 19484 21548
rect 21824 21496 21876 21548
rect 22192 21496 22244 21548
rect 20076 21428 20128 21480
rect 22008 21428 22060 21480
rect 23480 21564 23532 21616
rect 23572 21564 23624 21616
rect 23204 21496 23256 21548
rect 14648 21360 14700 21412
rect 19616 21360 19668 21412
rect 20444 21292 20496 21344
rect 22376 21292 22428 21344
rect 25320 21428 25372 21480
rect 22928 21292 22980 21344
rect 23572 21292 23624 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 12440 21088 12492 21140
rect 16212 21088 16264 21140
rect 17040 21088 17092 21140
rect 22100 21088 22152 21140
rect 23940 21088 23992 21140
rect 21272 21020 21324 21072
rect 22192 21063 22244 21072
rect 22192 21029 22201 21063
rect 22201 21029 22235 21063
rect 22235 21029 22244 21063
rect 22192 21020 22244 21029
rect 22744 21020 22796 21072
rect 23388 21020 23440 21072
rect 9588 20952 9640 21004
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 12624 20952 12676 21004
rect 16028 20952 16080 21004
rect 16488 20952 16540 21004
rect 19524 20952 19576 21004
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 22376 20952 22428 21004
rect 23848 20952 23900 21004
rect 6552 20884 6604 20936
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 16580 20884 16632 20936
rect 19708 20884 19760 20936
rect 19892 20927 19944 20936
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21824 20884 21876 20936
rect 22100 20884 22152 20936
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 24952 20884 25004 20936
rect 8484 20816 8536 20868
rect 10876 20816 10928 20868
rect 11428 20816 11480 20868
rect 15752 20816 15804 20868
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 13452 20748 13504 20800
rect 14372 20748 14424 20800
rect 19984 20816 20036 20868
rect 25136 20816 25188 20868
rect 24860 20748 24912 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 9496 20544 9548 20596
rect 14740 20544 14792 20596
rect 15476 20587 15528 20596
rect 15476 20553 15485 20587
rect 15485 20553 15519 20587
rect 15519 20553 15528 20587
rect 15476 20544 15528 20553
rect 8484 20476 8536 20528
rect 9772 20476 9824 20528
rect 11428 20476 11480 20528
rect 13452 20476 13504 20528
rect 14372 20476 14424 20528
rect 16580 20476 16632 20528
rect 6552 20408 6604 20460
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 9588 20408 9640 20460
rect 8576 20340 8628 20392
rect 9680 20340 9732 20392
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 19340 20544 19392 20596
rect 22100 20587 22152 20596
rect 22100 20553 22109 20587
rect 22109 20553 22143 20587
rect 22143 20553 22152 20587
rect 22100 20544 22152 20553
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 17132 20519 17184 20528
rect 17132 20485 17141 20519
rect 17141 20485 17175 20519
rect 17175 20485 17184 20519
rect 17132 20476 17184 20485
rect 17408 20476 17460 20528
rect 23572 20476 23624 20528
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 13360 20340 13412 20392
rect 17500 20340 17552 20392
rect 18144 20340 18196 20392
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 18604 20340 18656 20349
rect 20168 20408 20220 20460
rect 22560 20408 22612 20460
rect 21180 20340 21232 20392
rect 22100 20340 22152 20392
rect 22744 20340 22796 20392
rect 25136 20340 25188 20392
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 17776 20204 17828 20256
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 22652 20204 22704 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 8392 20000 8444 20052
rect 9220 20000 9272 20052
rect 13912 20000 13964 20052
rect 15752 20000 15804 20052
rect 16120 20000 16172 20052
rect 19340 20000 19392 20052
rect 20168 20000 20220 20052
rect 20812 20000 20864 20052
rect 7840 19864 7892 19916
rect 10692 19864 10744 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12716 19864 12768 19916
rect 14924 19864 14976 19916
rect 17132 19864 17184 19916
rect 18144 19864 18196 19916
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 17868 19796 17920 19848
rect 19156 19796 19208 19848
rect 8484 19728 8536 19780
rect 11428 19728 11480 19780
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 11888 19660 11940 19712
rect 16580 19728 16632 19780
rect 17040 19728 17092 19780
rect 17408 19728 17460 19780
rect 15936 19660 15988 19712
rect 19248 19728 19300 19780
rect 17868 19703 17920 19712
rect 17868 19669 17877 19703
rect 17877 19669 17911 19703
rect 17911 19669 17920 19703
rect 17868 19660 17920 19669
rect 19156 19660 19208 19712
rect 20260 19864 20312 19916
rect 22744 19864 22796 19916
rect 23572 20000 23624 20052
rect 23848 20043 23900 20052
rect 23848 20009 23857 20043
rect 23857 20009 23891 20043
rect 23891 20009 23900 20043
rect 23848 20000 23900 20009
rect 24032 19796 24084 19848
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 20812 19660 20864 19712
rect 20904 19660 20956 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 11428 19456 11480 19508
rect 8484 19388 8536 19440
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 10048 19320 10100 19372
rect 11704 19320 11756 19372
rect 12716 19388 12768 19440
rect 13728 19456 13780 19508
rect 14096 19456 14148 19508
rect 14924 19499 14976 19508
rect 14924 19465 14933 19499
rect 14933 19465 14967 19499
rect 14967 19465 14976 19499
rect 14924 19456 14976 19465
rect 16304 19388 16356 19440
rect 15108 19363 15160 19372
rect 15108 19329 15117 19363
rect 15117 19329 15151 19363
rect 15151 19329 15160 19363
rect 15108 19320 15160 19329
rect 16764 19456 16816 19508
rect 17316 19456 17368 19508
rect 16856 19388 16908 19440
rect 18696 19388 18748 19440
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 20720 19456 20772 19508
rect 20812 19456 20864 19508
rect 24584 19456 24636 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 23572 19388 23624 19440
rect 23756 19388 23808 19440
rect 24124 19388 24176 19440
rect 17776 19320 17828 19372
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6920 19252 6972 19304
rect 7380 19252 7432 19304
rect 8576 19184 8628 19236
rect 14464 19252 14516 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 17316 19184 17368 19236
rect 20904 19252 20956 19304
rect 22836 19320 22888 19372
rect 22928 19252 22980 19304
rect 22284 19184 22336 19236
rect 23296 19184 23348 19236
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 9220 19116 9272 19168
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 21088 19116 21140 19168
rect 23388 19116 23440 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8392 18955 8444 18964
rect 8392 18921 8401 18955
rect 8401 18921 8435 18955
rect 8435 18921 8444 18955
rect 8392 18912 8444 18921
rect 10784 18912 10836 18964
rect 16672 18912 16724 18964
rect 10416 18844 10468 18896
rect 8300 18776 8352 18828
rect 11612 18844 11664 18896
rect 10876 18776 10928 18828
rect 6552 18708 6604 18760
rect 8484 18708 8536 18760
rect 9956 18708 10008 18760
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 12440 18708 12492 18760
rect 18788 18844 18840 18896
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17776 18776 17828 18828
rect 16856 18708 16908 18760
rect 17500 18708 17552 18760
rect 7564 18572 7616 18624
rect 12532 18640 12584 18692
rect 21088 18912 21140 18964
rect 21180 18912 21232 18964
rect 22560 18844 22612 18896
rect 19340 18776 19392 18828
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 21456 18708 21508 18760
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 23572 18708 23624 18760
rect 10508 18615 10560 18624
rect 10508 18581 10517 18615
rect 10517 18581 10551 18615
rect 10551 18581 10560 18615
rect 10508 18572 10560 18581
rect 10876 18572 10928 18624
rect 21916 18640 21968 18692
rect 22008 18640 22060 18692
rect 25504 18640 25556 18692
rect 15660 18572 15712 18624
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 18788 18572 18840 18624
rect 20720 18572 20772 18624
rect 24124 18572 24176 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 9588 18368 9640 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10508 18368 10560 18420
rect 8484 18300 8536 18352
rect 9220 18300 9272 18352
rect 10140 18232 10192 18284
rect 6552 18164 6604 18216
rect 10784 18300 10836 18352
rect 12808 18300 12860 18352
rect 17224 18368 17276 18420
rect 22008 18368 22060 18420
rect 17040 18300 17092 18352
rect 25688 18368 25740 18420
rect 23664 18300 23716 18352
rect 24032 18300 24084 18352
rect 12532 18232 12584 18284
rect 9588 18096 9640 18148
rect 14188 18207 14240 18216
rect 14188 18173 14197 18207
rect 14197 18173 14231 18207
rect 14231 18173 14240 18207
rect 14188 18164 14240 18173
rect 16488 18232 16540 18284
rect 19248 18232 19300 18284
rect 16396 18164 16448 18216
rect 18604 18164 18656 18216
rect 22744 18232 22796 18284
rect 24216 18164 24268 18216
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 15108 18096 15160 18148
rect 23296 18096 23348 18148
rect 10784 18028 10836 18080
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 20904 18028 20956 18080
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 7656 17824 7708 17876
rect 7748 17688 7800 17740
rect 9680 17688 9732 17740
rect 12532 17824 12584 17876
rect 12624 17824 12676 17876
rect 12900 17824 12952 17876
rect 13544 17824 13596 17876
rect 14280 17824 14332 17876
rect 20168 17824 20220 17876
rect 7380 17663 7432 17672
rect 7380 17629 7389 17663
rect 7389 17629 7423 17663
rect 7423 17629 7432 17663
rect 7380 17620 7432 17629
rect 9404 17620 9456 17672
rect 9588 17620 9640 17672
rect 12808 17756 12860 17808
rect 11612 17688 11664 17740
rect 12256 17688 12308 17740
rect 12716 17688 12768 17740
rect 18420 17731 18472 17740
rect 18420 17697 18429 17731
rect 18429 17697 18463 17731
rect 18463 17697 18472 17731
rect 18420 17688 18472 17697
rect 18604 17731 18656 17740
rect 18604 17697 18613 17731
rect 18613 17697 18647 17731
rect 18647 17697 18656 17731
rect 18604 17688 18656 17697
rect 9220 17552 9272 17604
rect 9956 17484 10008 17536
rect 10232 17484 10284 17536
rect 10968 17484 11020 17536
rect 13636 17663 13688 17672
rect 13636 17629 13645 17663
rect 13645 17629 13679 17663
rect 13679 17629 13688 17663
rect 13636 17620 13688 17629
rect 16120 17620 16172 17672
rect 16948 17620 17000 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 25780 17756 25832 17808
rect 24860 17688 24912 17740
rect 24952 17688 25004 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 22560 17620 22612 17672
rect 17224 17552 17276 17604
rect 17684 17552 17736 17604
rect 18880 17552 18932 17604
rect 18972 17552 19024 17604
rect 20996 17552 21048 17604
rect 12624 17484 12676 17536
rect 15200 17484 15252 17536
rect 16856 17484 16908 17536
rect 21824 17552 21876 17604
rect 22652 17484 22704 17536
rect 22836 17484 22888 17536
rect 24676 17484 24728 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7380 17280 7432 17332
rect 9312 17280 9364 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11796 17280 11848 17332
rect 12440 17280 12492 17332
rect 13636 17280 13688 17332
rect 3516 17144 3568 17196
rect 9588 17212 9640 17264
rect 8668 17144 8720 17196
rect 3332 17076 3384 17128
rect 8944 17076 8996 17128
rect 9404 17076 9456 17128
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 11612 17144 11664 17196
rect 14188 17212 14240 17264
rect 13636 17144 13688 17196
rect 16488 17280 16540 17332
rect 16580 17280 16632 17332
rect 20444 17280 20496 17332
rect 24308 17280 24360 17332
rect 16948 17255 17000 17264
rect 16948 17221 16957 17255
rect 16957 17221 16991 17255
rect 16991 17221 17000 17255
rect 16948 17212 17000 17221
rect 18512 17212 18564 17264
rect 18696 17212 18748 17264
rect 17040 17144 17092 17196
rect 12900 17076 12952 17128
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 15476 17076 15528 17128
rect 16028 17076 16080 17128
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 24860 17212 24912 17264
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 24124 17187 24176 17196
rect 24124 17153 24133 17187
rect 24133 17153 24167 17187
rect 24167 17153 24176 17187
rect 24124 17144 24176 17153
rect 7472 17008 7524 17060
rect 12624 17008 12676 17060
rect 15936 17008 15988 17060
rect 17132 17051 17184 17060
rect 17132 17017 17141 17051
rect 17141 17017 17175 17051
rect 17175 17017 17184 17051
rect 17132 17008 17184 17017
rect 25320 17144 25372 17196
rect 24768 17119 24820 17128
rect 24768 17085 24777 17119
rect 24777 17085 24811 17119
rect 24811 17085 24820 17119
rect 24768 17076 24820 17085
rect 15384 16940 15436 16992
rect 16396 16940 16448 16992
rect 22008 17008 22060 17060
rect 22468 17008 22520 17060
rect 22652 17008 22704 17060
rect 17960 16940 18012 16992
rect 20444 16940 20496 16992
rect 24032 16940 24084 16992
rect 24768 16940 24820 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 8484 16736 8536 16788
rect 9036 16736 9088 16788
rect 9496 16600 9548 16652
rect 12716 16736 12768 16788
rect 14096 16736 14148 16788
rect 15108 16736 15160 16788
rect 17040 16736 17092 16788
rect 17500 16736 17552 16788
rect 21088 16736 21140 16788
rect 14740 16668 14792 16720
rect 17960 16668 18012 16720
rect 7472 16532 7524 16584
rect 9036 16532 9088 16584
rect 11428 16464 11480 16516
rect 12808 16464 12860 16516
rect 8852 16396 8904 16448
rect 11152 16396 11204 16448
rect 13452 16396 13504 16448
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16212 16600 16264 16609
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 16580 16600 16632 16652
rect 19432 16600 19484 16652
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 16028 16532 16080 16584
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 14832 16464 14884 16516
rect 15660 16396 15712 16448
rect 17868 16532 17920 16584
rect 19800 16532 19852 16584
rect 20444 16532 20496 16584
rect 17224 16464 17276 16516
rect 20168 16464 20220 16516
rect 21088 16532 21140 16584
rect 21456 16532 21508 16584
rect 22284 16532 22336 16584
rect 22376 16532 22428 16584
rect 17776 16396 17828 16448
rect 19340 16396 19392 16448
rect 20536 16396 20588 16448
rect 22100 16464 22152 16516
rect 24860 16464 24912 16516
rect 21548 16396 21600 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 9772 16192 9824 16244
rect 10508 16192 10560 16244
rect 11888 16192 11940 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 14372 16192 14424 16244
rect 14832 16192 14884 16244
rect 17408 16192 17460 16244
rect 7472 16124 7524 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 7840 15988 7892 16040
rect 9588 15988 9640 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 11888 15988 11940 16040
rect 12256 15988 12308 16040
rect 13544 16124 13596 16176
rect 5172 15852 5224 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8576 15852 8628 15904
rect 13636 15988 13688 16040
rect 17592 16124 17644 16176
rect 17868 16192 17920 16244
rect 20168 16192 20220 16244
rect 21364 16192 21416 16244
rect 22652 16192 22704 16244
rect 23296 16192 23348 16244
rect 21456 16124 21508 16176
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 15660 16056 15712 16108
rect 18328 16056 18380 16108
rect 19340 16056 19392 16108
rect 19432 16056 19484 16108
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 20076 15988 20128 16040
rect 20352 15988 20404 16040
rect 18144 15920 18196 15972
rect 11612 15852 11664 15904
rect 16304 15852 16356 15904
rect 17408 15852 17460 15904
rect 18420 15852 18472 15904
rect 20536 15852 20588 15904
rect 22652 15988 22704 16040
rect 24676 16056 24728 16108
rect 23664 15988 23716 16040
rect 24768 15988 24820 16040
rect 22652 15852 22704 15904
rect 24032 15852 24084 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 12624 15648 12676 15700
rect 14188 15648 14240 15700
rect 18604 15648 18656 15700
rect 22008 15648 22060 15700
rect 11336 15580 11388 15632
rect 13636 15580 13688 15632
rect 17684 15580 17736 15632
rect 9588 15512 9640 15564
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 12808 15512 12860 15564
rect 15200 15512 15252 15564
rect 16580 15512 16632 15564
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 17592 15444 17644 15496
rect 12624 15376 12676 15428
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 9588 15351 9640 15360
rect 9588 15317 9597 15351
rect 9597 15317 9631 15351
rect 9631 15317 9640 15351
rect 9588 15308 9640 15317
rect 10232 15308 10284 15360
rect 10600 15308 10652 15360
rect 12808 15308 12860 15360
rect 17500 15308 17552 15360
rect 20260 15512 20312 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 22652 15512 22704 15564
rect 23296 15512 23348 15564
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 23664 15444 23716 15496
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 21456 15376 21508 15428
rect 22100 15376 22152 15428
rect 22560 15376 22612 15428
rect 19524 15308 19576 15360
rect 20076 15308 20128 15360
rect 23480 15308 23532 15360
rect 24584 15351 24636 15360
rect 24584 15317 24593 15351
rect 24593 15317 24627 15351
rect 24627 15317 24636 15351
rect 24584 15308 24636 15317
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 13728 15104 13780 15156
rect 14464 15104 14516 15156
rect 15844 15104 15896 15156
rect 19984 15147 20036 15156
rect 19984 15113 19993 15147
rect 19993 15113 20027 15147
rect 20027 15113 20036 15147
rect 19984 15104 20036 15113
rect 20628 15104 20680 15156
rect 22192 15104 22244 15156
rect 22560 15104 22612 15156
rect 23296 15104 23348 15156
rect 7472 15036 7524 15088
rect 9680 15036 9732 15088
rect 11980 15036 12032 15088
rect 20168 15036 20220 15088
rect 6368 14900 6420 14952
rect 8300 14900 8352 14952
rect 11612 14968 11664 15020
rect 19340 14968 19392 15020
rect 20996 14968 21048 15020
rect 22008 14968 22060 15020
rect 22560 14968 22612 15020
rect 9036 14832 9088 14884
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 14096 14900 14148 14909
rect 15752 14900 15804 14952
rect 16028 14943 16080 14952
rect 16028 14909 16037 14943
rect 16037 14909 16071 14943
rect 16071 14909 16080 14943
rect 16028 14900 16080 14909
rect 16488 14900 16540 14952
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 22652 14900 22704 14952
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 13636 14832 13688 14884
rect 18880 14832 18932 14884
rect 21916 14832 21968 14884
rect 9956 14764 10008 14816
rect 12256 14764 12308 14816
rect 16396 14764 16448 14816
rect 18696 14764 18748 14816
rect 23572 14764 23624 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7748 14560 7800 14612
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 9312 14424 9364 14476
rect 11888 14424 11940 14476
rect 12072 14424 12124 14476
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 19524 14560 19576 14612
rect 26700 14560 26752 14612
rect 16488 14492 16540 14544
rect 17868 14492 17920 14544
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 15384 14424 15436 14476
rect 15476 14424 15528 14476
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 19616 14356 19668 14408
rect 23664 14356 23716 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 7380 14288 7432 14340
rect 9772 14220 9824 14272
rect 11244 14288 11296 14340
rect 13544 14288 13596 14340
rect 12716 14220 12768 14272
rect 13268 14220 13320 14272
rect 14924 14220 14976 14272
rect 20352 14288 20404 14340
rect 22284 14288 22336 14340
rect 16672 14220 16724 14272
rect 19984 14220 20036 14272
rect 23296 14220 23348 14272
rect 24124 14220 24176 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 7472 14016 7524 14068
rect 7748 13948 7800 14000
rect 8852 14016 8904 14068
rect 8484 13948 8536 14000
rect 9772 13991 9824 14000
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 9956 13948 10008 14000
rect 13268 13948 13320 14000
rect 11888 13880 11940 13932
rect 15200 13880 15252 13932
rect 16120 13880 16172 13932
rect 17592 13948 17644 14000
rect 18972 14016 19024 14068
rect 24768 14016 24820 14068
rect 19248 13948 19300 14000
rect 21640 13948 21692 14000
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 20812 13880 20864 13932
rect 24584 13948 24636 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 7288 13812 7340 13864
rect 8484 13812 8536 13864
rect 10968 13812 11020 13864
rect 12532 13812 12584 13864
rect 11244 13744 11296 13796
rect 11520 13744 11572 13796
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 15476 13812 15528 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17592 13812 17644 13864
rect 19064 13812 19116 13864
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 24860 13812 24912 13864
rect 11060 13676 11112 13728
rect 12440 13676 12492 13728
rect 13636 13676 13688 13728
rect 13912 13676 13964 13728
rect 14280 13676 14332 13728
rect 17316 13676 17368 13728
rect 18328 13676 18380 13728
rect 20168 13676 20220 13728
rect 21824 13744 21876 13796
rect 21088 13676 21140 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 7840 13472 7892 13524
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 9312 13472 9364 13524
rect 6368 13336 6420 13388
rect 7288 13336 7340 13388
rect 9864 13404 9916 13456
rect 11152 13472 11204 13524
rect 13912 13472 13964 13524
rect 14924 13472 14976 13524
rect 15476 13472 15528 13524
rect 13820 13404 13872 13456
rect 9128 13268 9180 13320
rect 12072 13336 12124 13388
rect 13636 13336 13688 13388
rect 15660 13404 15712 13456
rect 16212 13404 16264 13456
rect 19892 13404 19944 13456
rect 20168 13404 20220 13456
rect 26056 13404 26108 13456
rect 15384 13336 15436 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 7472 13200 7524 13252
rect 10600 13200 10652 13252
rect 9772 13132 9824 13184
rect 11244 13200 11296 13252
rect 13452 13268 13504 13320
rect 14464 13268 14516 13320
rect 14556 13200 14608 13252
rect 17316 13268 17368 13320
rect 17776 13268 17828 13320
rect 21364 13336 21416 13388
rect 23388 13336 23440 13388
rect 23480 13336 23532 13388
rect 17868 13243 17920 13252
rect 17868 13209 17877 13243
rect 17877 13209 17911 13243
rect 17911 13209 17920 13243
rect 17868 13200 17920 13209
rect 18512 13200 18564 13252
rect 18604 13243 18656 13252
rect 18604 13209 18613 13243
rect 18613 13209 18647 13243
rect 18647 13209 18656 13243
rect 18604 13200 18656 13209
rect 20260 13243 20312 13252
rect 20260 13209 20269 13243
rect 20269 13209 20303 13243
rect 20303 13209 20312 13243
rect 20260 13200 20312 13209
rect 20352 13200 20404 13252
rect 24032 13268 24084 13320
rect 24952 13200 25004 13252
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 13636 13132 13688 13184
rect 14004 13132 14056 13184
rect 14648 13132 14700 13184
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 15660 13175 15712 13184
rect 15660 13141 15669 13175
rect 15669 13141 15703 13175
rect 15703 13141 15712 13175
rect 15660 13132 15712 13141
rect 16580 13132 16632 13184
rect 21180 13132 21232 13184
rect 24584 13175 24636 13184
rect 24584 13141 24593 13175
rect 24593 13141 24627 13175
rect 24627 13141 24636 13175
rect 24584 13132 24636 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 6920 12860 6972 12912
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 4160 12724 4212 12776
rect 7564 12928 7616 12980
rect 9588 12928 9640 12980
rect 8300 12860 8352 12912
rect 9496 12860 9548 12912
rect 11060 12928 11112 12980
rect 11888 12903 11940 12912
rect 11888 12869 11897 12903
rect 11897 12869 11931 12903
rect 11931 12869 11940 12903
rect 11888 12860 11940 12869
rect 4252 12656 4304 12708
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 12440 12792 12492 12844
rect 9772 12724 9824 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 11704 12724 11756 12776
rect 15016 12928 15068 12980
rect 13820 12860 13872 12912
rect 13912 12860 13964 12912
rect 13728 12792 13780 12844
rect 15108 12860 15160 12912
rect 15660 12928 15712 12980
rect 16672 12928 16724 12980
rect 16764 12928 16816 12980
rect 18328 12860 18380 12912
rect 17408 12792 17460 12844
rect 20352 12928 20404 12980
rect 21272 12928 21324 12980
rect 22560 12928 22612 12980
rect 20996 12860 21048 12912
rect 23296 12903 23348 12912
rect 10324 12656 10376 12708
rect 10600 12656 10652 12708
rect 12348 12656 12400 12708
rect 13820 12724 13872 12776
rect 14004 12724 14056 12776
rect 13912 12656 13964 12708
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 14924 12724 14976 12776
rect 16028 12724 16080 12776
rect 12440 12588 12492 12640
rect 16764 12656 16816 12708
rect 18972 12724 19024 12776
rect 18880 12588 18932 12640
rect 19800 12792 19852 12844
rect 20720 12792 20772 12844
rect 20536 12724 20588 12776
rect 23296 12869 23305 12903
rect 23305 12869 23339 12903
rect 23339 12869 23348 12903
rect 23296 12860 23348 12869
rect 23756 12860 23808 12912
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22836 12724 22888 12776
rect 19892 12699 19944 12708
rect 19892 12665 19901 12699
rect 19901 12665 19935 12699
rect 19935 12665 19944 12699
rect 19892 12656 19944 12665
rect 24676 12724 24728 12776
rect 22100 12588 22152 12640
rect 23388 12588 23440 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 7012 12384 7064 12436
rect 8300 12384 8352 12436
rect 10048 12384 10100 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 14832 12384 14884 12436
rect 18604 12384 18656 12436
rect 20996 12384 21048 12436
rect 10140 12316 10192 12368
rect 10508 12316 10560 12368
rect 11796 12316 11848 12368
rect 12532 12316 12584 12368
rect 14556 12316 14608 12368
rect 15108 12316 15160 12368
rect 16672 12316 16724 12368
rect 17040 12316 17092 12368
rect 17224 12316 17276 12368
rect 17316 12316 17368 12368
rect 17684 12316 17736 12368
rect 9220 12248 9272 12300
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 13360 12248 13412 12300
rect 17040 12180 17092 12232
rect 19156 12248 19208 12300
rect 20260 12248 20312 12300
rect 17776 12180 17828 12232
rect 19248 12180 19300 12232
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 22100 12180 22152 12232
rect 22284 12180 22336 12232
rect 24584 12248 24636 12300
rect 23572 12180 23624 12232
rect 12532 12112 12584 12164
rect 12900 12112 12952 12164
rect 13728 12112 13780 12164
rect 14464 12112 14516 12164
rect 16856 12112 16908 12164
rect 19156 12112 19208 12164
rect 20720 12112 20772 12164
rect 23664 12112 23716 12164
rect 24952 12112 25004 12164
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 12624 12044 12676 12096
rect 14648 12044 14700 12096
rect 15016 12044 15068 12096
rect 17500 12044 17552 12096
rect 18512 12044 18564 12096
rect 19708 12044 19760 12096
rect 23480 12044 23532 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 9220 11840 9272 11892
rect 9864 11840 9916 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 12440 11840 12492 11892
rect 12808 11840 12860 11892
rect 13268 11840 13320 11892
rect 14188 11840 14240 11892
rect 14832 11840 14884 11892
rect 12716 11772 12768 11824
rect 13360 11772 13412 11824
rect 13728 11772 13780 11824
rect 16672 11840 16724 11892
rect 16948 11840 17000 11892
rect 19340 11840 19392 11892
rect 20628 11840 20680 11892
rect 8576 11704 8628 11756
rect 9864 11704 9916 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 11060 11636 11112 11688
rect 10968 11568 11020 11620
rect 12072 11568 12124 11620
rect 12440 11500 12492 11552
rect 13268 11568 13320 11620
rect 15292 11772 15344 11824
rect 14096 11704 14148 11756
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 14556 11568 14608 11620
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 12808 11500 12860 11552
rect 13452 11500 13504 11552
rect 13728 11500 13780 11552
rect 17408 11772 17460 11824
rect 22192 11840 22244 11892
rect 21088 11772 21140 11824
rect 22376 11815 22428 11824
rect 22376 11781 22385 11815
rect 22385 11781 22419 11815
rect 22419 11781 22428 11815
rect 22376 11772 22428 11781
rect 23388 11815 23440 11824
rect 23388 11781 23397 11815
rect 23397 11781 23431 11815
rect 23431 11781 23440 11815
rect 23388 11772 23440 11781
rect 23664 11772 23716 11824
rect 16304 11636 16356 11688
rect 19616 11704 19668 11756
rect 21640 11704 21692 11756
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22284 11704 22336 11756
rect 22836 11704 22888 11756
rect 19432 11636 19484 11688
rect 19524 11568 19576 11620
rect 17776 11500 17828 11552
rect 19800 11500 19852 11552
rect 21548 11568 21600 11620
rect 22652 11568 22704 11620
rect 22100 11500 22152 11552
rect 24860 11543 24912 11552
rect 24860 11509 24869 11543
rect 24869 11509 24903 11543
rect 24903 11509 24912 11543
rect 24860 11500 24912 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 10600 11296 10652 11348
rect 12992 11296 13044 11348
rect 13728 11296 13780 11348
rect 12164 11160 12216 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 10508 11092 10560 11144
rect 11060 11092 11112 11144
rect 13544 11160 13596 11212
rect 15200 11296 15252 11348
rect 17408 11296 17460 11348
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 22376 11296 22428 11348
rect 23296 11296 23348 11348
rect 16304 11228 16356 11280
rect 16856 11160 16908 11212
rect 18328 11203 18380 11212
rect 18328 11169 18337 11203
rect 18337 11169 18371 11203
rect 18371 11169 18380 11203
rect 18328 11160 18380 11169
rect 19616 11160 19668 11212
rect 23848 11228 23900 11280
rect 21180 11160 21232 11212
rect 21272 11160 21324 11212
rect 16120 11092 16172 11144
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 12808 11024 12860 11076
rect 9680 10956 9732 11008
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 12624 10956 12676 11008
rect 13728 10956 13780 11008
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 17408 11135 17460 11144
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 18604 11092 18656 11144
rect 20168 11135 20220 11144
rect 20168 11101 20177 11135
rect 20177 11101 20211 11135
rect 20211 11101 20220 11135
rect 20168 11092 20220 11101
rect 17960 11024 18012 11076
rect 15200 10956 15252 11008
rect 15660 10956 15712 11008
rect 19524 11024 19576 11076
rect 22744 11092 22796 11144
rect 20444 11024 20496 11076
rect 21916 11024 21968 11076
rect 24676 11092 24728 11144
rect 22008 10956 22060 11008
rect 22744 10999 22796 11008
rect 22744 10965 22753 10999
rect 22753 10965 22787 10999
rect 22787 10965 22796 10999
rect 22744 10956 22796 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 9772 10752 9824 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 15108 10752 15160 10804
rect 7104 10684 7156 10736
rect 9864 10684 9916 10736
rect 10600 10684 10652 10736
rect 7288 10548 7340 10600
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 8944 10548 8996 10600
rect 14004 10684 14056 10736
rect 17684 10752 17736 10804
rect 15936 10727 15988 10736
rect 15936 10693 15945 10727
rect 15945 10693 15979 10727
rect 15979 10693 15988 10727
rect 15936 10684 15988 10693
rect 15568 10616 15620 10668
rect 24032 10752 24084 10804
rect 19616 10684 19668 10736
rect 21364 10684 21416 10736
rect 13912 10548 13964 10600
rect 13452 10480 13504 10532
rect 14832 10548 14884 10600
rect 15844 10548 15896 10600
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11980 10412 12032 10464
rect 13360 10412 13412 10464
rect 17316 10548 17368 10600
rect 18052 10548 18104 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 21088 10616 21140 10668
rect 18788 10548 18840 10600
rect 16856 10480 16908 10532
rect 20720 10548 20772 10600
rect 21456 10591 21508 10600
rect 21456 10557 21465 10591
rect 21465 10557 21499 10591
rect 21499 10557 21508 10591
rect 21456 10548 21508 10557
rect 22560 10616 22612 10668
rect 24584 10616 24636 10668
rect 22652 10548 22704 10600
rect 24860 10616 24912 10668
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 16396 10412 16448 10464
rect 19340 10412 19392 10464
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 22100 10412 22152 10464
rect 23480 10480 23532 10532
rect 23572 10412 23624 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 13360 10208 13412 10260
rect 13452 10208 13504 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 17960 10208 18012 10260
rect 22560 10208 22612 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 10876 10140 10928 10192
rect 8208 10072 8260 10124
rect 9588 10072 9640 10124
rect 11428 10072 11480 10124
rect 12348 10140 12400 10192
rect 15476 10140 15528 10192
rect 13544 10072 13596 10124
rect 14924 10072 14976 10124
rect 17316 10072 17368 10124
rect 17868 10072 17920 10124
rect 18236 10140 18288 10192
rect 18420 10140 18472 10192
rect 22100 10140 22152 10192
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 13728 10004 13780 10056
rect 9036 9936 9088 9988
rect 10600 9936 10652 9988
rect 11152 9936 11204 9988
rect 15292 9936 15344 9988
rect 17592 9936 17644 9988
rect 20076 10072 20128 10124
rect 21180 10072 21232 10124
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 22284 10115 22336 10124
rect 22284 10081 22293 10115
rect 22293 10081 22327 10115
rect 22327 10081 22336 10115
rect 22284 10072 22336 10081
rect 22652 10072 22704 10124
rect 20812 10004 20864 10056
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 23664 10004 23716 10056
rect 23848 10004 23900 10056
rect 19432 9936 19484 9988
rect 20536 9936 20588 9988
rect 7104 9868 7156 9920
rect 14832 9868 14884 9920
rect 15108 9868 15160 9920
rect 16488 9868 16540 9920
rect 16764 9868 16816 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 18052 9868 18104 9920
rect 18788 9868 18840 9920
rect 19708 9868 19760 9920
rect 22652 9936 22704 9988
rect 22836 9868 22888 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 9772 9664 9824 9716
rect 15292 9664 15344 9716
rect 10600 9596 10652 9648
rect 14556 9596 14608 9648
rect 10784 9460 10836 9512
rect 12532 9460 12584 9512
rect 14280 9460 14332 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14924 9460 14976 9512
rect 17316 9664 17368 9716
rect 17500 9664 17552 9716
rect 22192 9664 22244 9716
rect 22652 9664 22704 9716
rect 24400 9664 24452 9716
rect 17868 9596 17920 9648
rect 18604 9596 18656 9648
rect 19984 9596 20036 9648
rect 20352 9596 20404 9648
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 19248 9528 19300 9580
rect 23388 9528 23440 9580
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 17500 9460 17552 9512
rect 12348 9324 12400 9376
rect 15200 9435 15252 9444
rect 15200 9401 15209 9435
rect 15209 9401 15243 9435
rect 15243 9401 15252 9435
rect 15200 9392 15252 9401
rect 17316 9392 17368 9444
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 14740 9324 14792 9376
rect 17132 9324 17184 9376
rect 17500 9324 17552 9376
rect 20168 9460 20220 9512
rect 20260 9392 20312 9444
rect 22560 9460 22612 9512
rect 22836 9460 22888 9512
rect 23572 9460 23624 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 20628 9392 20680 9444
rect 22192 9392 22244 9444
rect 22376 9392 22428 9444
rect 19064 9324 19116 9376
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 19984 9324 20036 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 11612 9163 11664 9172
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 10692 9052 10744 9104
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 10784 8984 10836 9036
rect 12072 8984 12124 9036
rect 16488 9120 16540 9172
rect 16672 9120 16724 9172
rect 19248 9120 19300 9172
rect 19892 9120 19944 9172
rect 21732 9120 21784 9172
rect 13360 9052 13412 9104
rect 17316 9052 17368 9104
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 13636 8984 13688 9036
rect 14004 8916 14056 8968
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 16120 8984 16172 9036
rect 17500 8984 17552 9036
rect 24676 9052 24728 9104
rect 19432 8984 19484 9036
rect 20168 9027 20220 9036
rect 20168 8993 20177 9027
rect 20177 8993 20211 9027
rect 20211 8993 20220 9027
rect 20168 8984 20220 8993
rect 15936 8916 15988 8968
rect 17132 8916 17184 8968
rect 18880 8955 18932 8968
rect 18880 8921 18889 8955
rect 18889 8921 18923 8955
rect 18923 8921 18932 8955
rect 18880 8916 18932 8921
rect 19248 8916 19300 8968
rect 9680 8848 9732 8900
rect 10692 8848 10744 8900
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 14464 8848 14516 8900
rect 19064 8848 19116 8900
rect 19524 8848 19576 8900
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 16672 8780 16724 8832
rect 19248 8780 19300 8832
rect 19432 8780 19484 8832
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 20812 8959 20864 8968
rect 20812 8925 20821 8959
rect 20821 8925 20855 8959
rect 20855 8925 20864 8959
rect 20812 8916 20864 8925
rect 20904 8916 20956 8968
rect 22744 8916 22796 8968
rect 21824 8891 21876 8900
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 24952 8848 25004 8900
rect 22008 8780 22060 8832
rect 24584 8823 24636 8832
rect 24584 8789 24593 8823
rect 24593 8789 24627 8823
rect 24627 8789 24636 8823
rect 24584 8780 24636 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12164 8576 12216 8628
rect 14096 8576 14148 8628
rect 14464 8576 14516 8628
rect 20168 8576 20220 8628
rect 7656 8508 7708 8560
rect 11520 8508 11572 8560
rect 13820 8508 13872 8560
rect 2228 8372 2280 8424
rect 14740 8440 14792 8492
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 17132 8440 17184 8492
rect 17500 8440 17552 8492
rect 17684 8440 17736 8492
rect 11152 8304 11204 8356
rect 16672 8372 16724 8424
rect 16948 8372 17000 8424
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 14648 8304 14700 8356
rect 17132 8304 17184 8356
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 19892 8508 19944 8560
rect 20260 8508 20312 8560
rect 21088 8440 21140 8492
rect 22468 8440 22520 8492
rect 23480 8440 23532 8492
rect 20720 8372 20772 8424
rect 21272 8372 21324 8424
rect 22376 8372 22428 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 13452 8236 13504 8288
rect 19340 8304 19392 8356
rect 19984 8279 20036 8288
rect 19984 8245 20014 8279
rect 20014 8245 20036 8279
rect 19984 8236 20036 8245
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 13728 8032 13780 8084
rect 12072 7964 12124 8016
rect 12532 7964 12584 8016
rect 16488 8032 16540 8084
rect 18328 8032 18380 8084
rect 18880 8032 18932 8084
rect 10876 7939 10928 7948
rect 10876 7905 10885 7939
rect 10885 7905 10919 7939
rect 10919 7905 10928 7939
rect 10876 7896 10928 7905
rect 10968 7896 11020 7948
rect 17408 7964 17460 8016
rect 20996 7964 21048 8016
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14464 7828 14516 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 16212 7896 16264 7948
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 19524 7896 19576 7948
rect 22192 8032 22244 8084
rect 24124 8032 24176 8084
rect 24216 7964 24268 8016
rect 15016 7828 15068 7880
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 22284 7939 22336 7948
rect 22284 7905 22293 7939
rect 22293 7905 22327 7939
rect 22327 7905 22336 7939
rect 22284 7896 22336 7905
rect 22560 7939 22612 7948
rect 22560 7905 22569 7939
rect 22569 7905 22603 7939
rect 22603 7905 22612 7939
rect 22560 7896 22612 7905
rect 23848 7896 23900 7948
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 5264 7760 5316 7812
rect 11336 7760 11388 7812
rect 10048 7692 10100 7744
rect 10324 7692 10376 7744
rect 10508 7692 10560 7744
rect 12072 7692 12124 7744
rect 12716 7760 12768 7812
rect 14280 7760 14332 7812
rect 16948 7760 17000 7812
rect 18880 7760 18932 7812
rect 20168 7760 20220 7812
rect 12808 7692 12860 7744
rect 12900 7692 12952 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 17316 7692 17368 7744
rect 17500 7692 17552 7744
rect 19340 7692 19392 7744
rect 21640 7803 21692 7812
rect 21640 7769 21649 7803
rect 21649 7769 21683 7803
rect 21683 7769 21692 7803
rect 21640 7760 21692 7769
rect 23664 7828 23716 7880
rect 24032 7735 24084 7744
rect 24032 7701 24041 7735
rect 24041 7701 24075 7735
rect 24075 7701 24084 7735
rect 24032 7692 24084 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 6736 7488 6788 7540
rect 10968 7488 11020 7540
rect 14740 7488 14792 7540
rect 15752 7488 15804 7540
rect 14280 7420 14332 7472
rect 15016 7420 15068 7472
rect 15568 7420 15620 7472
rect 17040 7463 17092 7472
rect 17040 7429 17049 7463
rect 17049 7429 17083 7463
rect 17083 7429 17092 7463
rect 17040 7420 17092 7429
rect 18420 7420 18472 7472
rect 10692 7352 10744 7404
rect 13452 7352 13504 7404
rect 15752 7352 15804 7404
rect 17500 7352 17552 7404
rect 19248 7352 19300 7404
rect 20720 7352 20772 7404
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 10876 7284 10928 7336
rect 11060 7284 11112 7336
rect 11704 7284 11756 7336
rect 9588 7148 9640 7200
rect 16304 7284 16356 7336
rect 16856 7284 16908 7336
rect 18604 7284 18656 7336
rect 18972 7284 19024 7336
rect 19616 7284 19668 7336
rect 21916 7284 21968 7336
rect 23296 7327 23348 7336
rect 23296 7293 23305 7327
rect 23305 7293 23339 7327
rect 23339 7293 23348 7327
rect 23296 7284 23348 7293
rect 17224 7259 17276 7268
rect 17224 7225 17233 7259
rect 17233 7225 17267 7259
rect 17267 7225 17276 7259
rect 17224 7216 17276 7225
rect 20628 7216 20680 7268
rect 24860 7216 24912 7268
rect 15108 7148 15160 7200
rect 16488 7148 16540 7200
rect 18328 7148 18380 7200
rect 18696 7148 18748 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 13820 6944 13872 6996
rect 19248 6944 19300 6996
rect 21456 6944 21508 6996
rect 22100 6944 22152 6996
rect 24032 6944 24084 6996
rect 5448 6808 5500 6860
rect 8852 6808 8904 6860
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 13360 6808 13412 6860
rect 15108 6876 15160 6928
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 13728 6740 13780 6792
rect 10692 6672 10744 6724
rect 9680 6604 9732 6656
rect 13268 6604 13320 6656
rect 15292 6740 15344 6792
rect 15476 6808 15528 6860
rect 17040 6808 17092 6860
rect 18696 6808 18748 6860
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 19340 6740 19392 6792
rect 21272 6740 21324 6792
rect 23664 6740 23716 6792
rect 20444 6672 20496 6724
rect 15200 6604 15252 6656
rect 15568 6604 15620 6656
rect 16028 6604 16080 6656
rect 19248 6604 19300 6656
rect 19984 6604 20036 6656
rect 21732 6604 21784 6656
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 24032 6604 24084 6656
rect 24952 6647 25004 6656
rect 24952 6613 24961 6647
rect 24961 6613 24995 6647
rect 24995 6613 25004 6647
rect 24952 6604 25004 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 12440 6400 12492 6452
rect 13728 6400 13780 6452
rect 15200 6400 15252 6452
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 17408 6400 17460 6452
rect 13268 6332 13320 6384
rect 18420 6332 18472 6384
rect 12808 6264 12860 6316
rect 13820 6264 13872 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 19524 6400 19576 6452
rect 23848 6400 23900 6452
rect 22560 6332 22612 6384
rect 25136 6375 25188 6384
rect 25136 6341 25145 6375
rect 25145 6341 25179 6375
rect 25179 6341 25188 6375
rect 25136 6332 25188 6341
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 21732 6264 21784 6316
rect 24584 6264 24636 6316
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 14832 6196 14884 6248
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 22100 6196 22152 6248
rect 14464 6060 14516 6112
rect 24032 6128 24084 6180
rect 20352 6060 20404 6112
rect 20444 6060 20496 6112
rect 22836 6060 22888 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 21732 5856 21784 5908
rect 10968 5720 11020 5772
rect 14924 5720 14976 5772
rect 20076 5788 20128 5840
rect 9588 5652 9640 5704
rect 13544 5652 13596 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 16120 5652 16172 5704
rect 10692 5584 10744 5636
rect 20444 5720 20496 5772
rect 22284 5720 22336 5772
rect 18604 5652 18656 5704
rect 19616 5652 19668 5704
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 25044 5652 25096 5704
rect 17592 5584 17644 5636
rect 20628 5584 20680 5636
rect 14188 5516 14240 5568
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 15016 5516 15068 5568
rect 20352 5516 20404 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 3884 5244 3936 5296
rect 10416 5244 10468 5296
rect 13360 5287 13412 5296
rect 13360 5253 13369 5287
rect 13369 5253 13403 5287
rect 13403 5253 13412 5287
rect 13360 5244 13412 5253
rect 15016 5244 15068 5296
rect 22744 5312 22796 5364
rect 17040 5244 17092 5296
rect 18420 5244 18472 5296
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 19892 5244 19944 5296
rect 21272 5244 21324 5296
rect 10784 5108 10836 5160
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 17132 5108 17184 5160
rect 19524 5108 19576 5160
rect 20628 5108 20680 5160
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 13912 4972 13964 5024
rect 14464 4972 14516 5024
rect 15936 4972 15988 5024
rect 21456 5083 21508 5092
rect 21456 5049 21465 5083
rect 21465 5049 21499 5083
rect 21499 5049 21508 5083
rect 21456 5040 21508 5049
rect 20628 4972 20680 5024
rect 21272 4972 21324 5024
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 15660 4768 15712 4820
rect 16212 4768 16264 4820
rect 17040 4768 17092 4820
rect 23388 4768 23440 4820
rect 24860 4743 24912 4752
rect 24860 4709 24869 4743
rect 24869 4709 24903 4743
rect 24903 4709 24912 4743
rect 24860 4700 24912 4709
rect 9588 4632 9640 4684
rect 13636 4632 13688 4684
rect 16856 4632 16908 4684
rect 17500 4632 17552 4684
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 20904 4632 20956 4684
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 5356 4539 5408 4548
rect 5356 4505 5365 4539
rect 5365 4505 5399 4539
rect 5399 4505 5408 4539
rect 5356 4496 5408 4505
rect 10692 4496 10744 4548
rect 18788 4564 18840 4616
rect 19800 4564 19852 4616
rect 21548 4564 21600 4616
rect 24400 4632 24452 4684
rect 24216 4564 24268 4616
rect 15384 4496 15436 4548
rect 15476 4539 15528 4548
rect 15476 4505 15485 4539
rect 15485 4505 15519 4539
rect 15519 4505 15528 4539
rect 15476 4496 15528 4505
rect 15016 4428 15068 4480
rect 18420 4496 18472 4548
rect 21088 4496 21140 4548
rect 19432 4428 19484 4480
rect 22468 4428 22520 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 15476 4224 15528 4276
rect 20168 4224 20220 4276
rect 14924 4156 14976 4208
rect 20904 4199 20956 4208
rect 20904 4165 20913 4199
rect 20913 4165 20947 4199
rect 20947 4165 20956 4199
rect 20904 4156 20956 4165
rect 1492 4088 1544 4140
rect 1860 4088 1912 4140
rect 4068 4088 4120 4140
rect 5908 4088 5960 4140
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16580 4088 16632 4140
rect 17224 4088 17276 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 22652 4156 22704 4208
rect 2228 3995 2280 4004
rect 2228 3961 2237 3995
rect 2237 3961 2271 3995
rect 2271 3961 2280 3995
rect 2228 3952 2280 3961
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 11796 3952 11848 4004
rect 5356 3884 5408 3936
rect 14832 4020 14884 4072
rect 16212 4020 16264 4072
rect 18328 4020 18380 4072
rect 21456 4020 21508 4072
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 16856 3952 16908 4004
rect 17684 3952 17736 4004
rect 19984 3952 20036 4004
rect 18052 3884 18104 3936
rect 18144 3884 18196 3936
rect 20996 3884 21048 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 3332 3680 3384 3732
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 7748 3680 7800 3732
rect 13820 3680 13872 3732
rect 16304 3680 16356 3732
rect 18052 3680 18104 3732
rect 25136 3680 25188 3732
rect 9404 3612 9456 3664
rect 15844 3612 15896 3664
rect 18788 3612 18840 3664
rect 19892 3612 19944 3664
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 12532 3544 12584 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 2228 3476 2280 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4804 3476 4856 3528
rect 6644 3476 6696 3528
rect 7840 3476 7892 3528
rect 9588 3476 9640 3528
rect 10692 3476 10744 3528
rect 12164 3476 12216 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 16396 3476 16448 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19708 3476 19760 3528
rect 20720 3476 20772 3528
rect 3608 3408 3660 3460
rect 3240 3340 3292 3392
rect 10048 3408 10100 3460
rect 14556 3408 14608 3460
rect 19156 3408 19208 3460
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 24860 3451 24912 3460
rect 24860 3417 24869 3451
rect 24869 3417 24903 3451
rect 24903 3417 24912 3451
rect 24860 3408 24912 3417
rect 9128 3340 9180 3392
rect 13728 3340 13780 3392
rect 19524 3340 19576 3392
rect 21088 3340 21140 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 9680 3136 9732 3188
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 12624 3136 12676 3188
rect 16028 3136 16080 3188
rect 2596 3000 2648 3052
rect 3240 2932 3292 2984
rect 3332 2932 3384 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 5264 2932 5316 2984
rect 7012 3000 7064 3052
rect 8484 3000 8536 3052
rect 8852 3000 8904 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 10324 3000 10376 3052
rect 11060 3000 11112 3052
rect 11796 3000 11848 3052
rect 14372 3068 14424 3120
rect 16580 3068 16632 3120
rect 20260 3136 20312 3188
rect 23204 3136 23256 3188
rect 23664 3136 23716 3188
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 14096 3000 14148 3052
rect 18420 3000 18472 3052
rect 18512 3000 18564 3052
rect 10140 2932 10192 2984
rect 9128 2796 9180 2848
rect 9772 2796 9824 2848
rect 11428 2932 11480 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 20720 3000 20772 3052
rect 22008 3068 22060 3120
rect 22284 3111 22336 3120
rect 22284 3077 22293 3111
rect 22293 3077 22327 3111
rect 22327 3077 22336 3111
rect 22284 3068 22336 3077
rect 22468 3000 22520 3052
rect 24308 3000 24360 3052
rect 16856 2864 16908 2916
rect 16948 2864 17000 2916
rect 19892 2864 19944 2916
rect 20628 2864 20680 2916
rect 21272 2864 21324 2916
rect 21364 2864 21416 2916
rect 22192 2864 22244 2916
rect 22284 2864 22336 2916
rect 22652 2864 22704 2916
rect 22744 2907 22796 2916
rect 22744 2873 22753 2907
rect 22753 2873 22787 2907
rect 22787 2873 22796 2907
rect 22744 2864 22796 2873
rect 12716 2796 12768 2848
rect 15108 2796 15160 2848
rect 17316 2796 17368 2848
rect 18420 2796 18472 2848
rect 22100 2796 22152 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 9036 2592 9088 2644
rect 10232 2524 10284 2576
rect 17132 2592 17184 2644
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 20904 2592 20956 2644
rect 21640 2592 21692 2644
rect 23204 2592 23256 2644
rect 24952 2592 25004 2644
rect 12348 2524 12400 2576
rect 16488 2524 16540 2576
rect 2964 2456 3016 2508
rect 5540 2456 5592 2508
rect 7656 2456 7708 2508
rect 14372 2456 14424 2508
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 7380 2388 7432 2440
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 6276 2320 6328 2372
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 12164 2388 12216 2440
rect 12900 2388 12952 2440
rect 14188 2388 14240 2440
rect 16764 2388 16816 2440
rect 9956 2320 10008 2372
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 14280 2320 14332 2372
rect 19064 2388 19116 2440
rect 22100 2456 22152 2508
rect 23756 2388 23808 2440
rect 10508 2252 10560 2304
rect 13452 2252 13504 2304
rect 19616 2320 19668 2372
rect 22836 2320 22888 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 9864 1980 9916 2032
rect 24860 1980 24912 2032
rect 10968 1912 11020 1964
rect 22100 1912 22152 1964
rect 3424 1844 3476 1896
rect 8760 1844 8812 1896
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3804 53650 3832 56200
rect 4068 54188 4120 54194
rect 4068 54130 4120 54136
rect 4804 54188 4856 54194
rect 4804 54130 4856 54136
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 4080 53242 4108 54130
rect 4068 53236 4120 53242
rect 4068 53178 4120 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 4816 51406 4844 54130
rect 5184 54126 5212 56200
rect 5172 54120 5224 54126
rect 5172 54062 5224 54068
rect 6564 53650 6592 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7380 54188 7432 54194
rect 7380 54130 7432 54136
rect 6552 53644 6604 53650
rect 6552 53586 6604 53592
rect 6644 53576 6696 53582
rect 6644 53518 6696 53524
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 4804 51400 4856 51406
rect 4804 51342 4856 51348
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 5552 50522 5580 53450
rect 6656 52154 6684 53518
rect 6644 52148 6696 52154
rect 6644 52090 6696 52096
rect 7392 51610 7420 54130
rect 7852 54126 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8576 54256 8628 54262
rect 8576 54198 8628 54204
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 7840 53576 7892 53582
rect 7840 53518 7892 53524
rect 7748 53100 7800 53106
rect 7748 53042 7800 53048
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 7760 50454 7788 53042
rect 7852 51542 7880 53518
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7840 51536 7892 51542
rect 7840 51478 7892 51484
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8392 50516 8444 50522
rect 8392 50458 8444 50464
rect 7748 50448 7800 50454
rect 7748 50390 7800 50396
rect 8300 50448 8352 50454
rect 8300 50390 8352 50396
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 8312 48142 8340 50390
rect 8404 48890 8432 50458
rect 8392 48884 8444 48890
rect 8392 48826 8444 48832
rect 8300 48136 8352 48142
rect 8300 48078 8352 48084
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8312 46578 8340 48078
rect 8300 46572 8352 46578
rect 8300 46514 8352 46520
rect 7840 46504 7892 46510
rect 7840 46446 7892 46452
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7852 38010 7880 46446
rect 8496 46442 8524 51342
rect 8588 50318 8616 54198
rect 9324 54126 9352 56200
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 9312 54120 9364 54126
rect 9312 54062 9364 54068
rect 9404 52012 9456 52018
rect 9404 51954 9456 51960
rect 8576 50312 8628 50318
rect 8576 50254 8628 50260
rect 8588 47666 8616 50254
rect 9128 48612 9180 48618
rect 9128 48554 9180 48560
rect 8576 47660 8628 47666
rect 8576 47602 8628 47608
rect 8484 46436 8536 46442
rect 8484 46378 8536 46384
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 9140 44946 9168 48554
rect 9416 47802 9444 51954
rect 9600 50522 9628 54130
rect 10704 53718 10732 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53712 10744 53718
rect 10692 53654 10744 53660
rect 10692 53576 10744 53582
rect 10692 53518 10744 53524
rect 10508 51400 10560 51406
rect 10508 51342 10560 51348
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 9588 50312 9640 50318
rect 9588 50254 9640 50260
rect 9496 48680 9548 48686
rect 9496 48622 9548 48628
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9404 47796 9456 47802
rect 9404 47738 9456 47744
rect 9232 47054 9260 47738
rect 9508 47462 9536 48622
rect 9496 47456 9548 47462
rect 9496 47398 9548 47404
rect 9220 47048 9272 47054
rect 9220 46990 9272 46996
rect 9128 44940 9180 44946
rect 9128 44882 9180 44888
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 9232 44402 9260 46990
rect 9508 45554 9536 47398
rect 9416 45526 9536 45554
rect 9416 45082 9444 45526
rect 9404 45076 9456 45082
rect 9404 45018 9456 45024
rect 9404 44940 9456 44946
rect 9404 44882 9456 44888
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 8944 44328 8996 44334
rect 8944 44270 8996 44276
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8852 42696 8904 42702
rect 8852 42638 8904 42644
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1504 800 1532 4082
rect 1872 800 1900 4082
rect 2240 4010 2268 8366
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3344 3738 3372 17070
rect 3436 6497 3464 22714
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6564 20466 6592 20878
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 19310 6592 20402
rect 7392 19310 7420 21626
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 6564 18766 6592 19246
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6564 18222 6592 18702
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3528 8809 3556 17138
rect 6564 16114 6592 18158
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3514 8800 3570 8809
rect 3514 8735 3570 8744
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3896 4185 3924 5238
rect 3882 4176 3938 4185
rect 3882 4111 3938 4120
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 800 2268 3470
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 800 2636 2994
rect 3252 2990 3280 3334
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 800 3004 2450
rect 3344 800 3372 2926
rect 3424 1896 3476 1902
rect 3422 1864 3424 1873
rect 3476 1864 3478 1873
rect 3620 1850 3648 3402
rect 3620 1822 3740 1850
rect 3422 1799 3478 1808
rect 3712 800 3740 1822
rect 4080 800 4108 4082
rect 4172 4010 4200 12718
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4264 3738 4292 12650
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 5184 3602 5212 15846
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6380 14482 6408 14894
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6380 13394 6408 14418
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6932 12918 6960 19246
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17338 7420 17614
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7484 17066 7512 24890
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 16182 7512 16526
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7484 15094 7512 16118
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 14362 7512 15030
rect 7392 14346 7512 14362
rect 7380 14340 7512 14346
rect 7432 14334 7512 14340
rect 7380 14282 7432 14288
rect 7484 14074 7512 14334
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13394 7328 13806
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12442 7052 12786
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7300 11694 7328 13330
rect 7484 13258 7512 14010
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7576 12986 7604 18566
rect 7668 17882 7696 30194
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8668 23792 8720 23798
rect 8668 23734 8720 23740
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7852 22642 7880 23598
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8404 22710 8432 23054
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 21554 7880 22578
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8404 21622 8432 22646
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7748 20460 7800 20466
rect 7852 20448 7880 21490
rect 8404 21434 8432 21558
rect 8404 21406 8524 21434
rect 8496 20874 8524 21406
rect 8588 21146 8616 23122
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8496 20534 8524 20810
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 7800 20420 7880 20448
rect 7748 20402 7800 20408
rect 7852 19922 7880 20420
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18834 8340 19110
rect 8404 18970 8432 19994
rect 8496 19786 8524 20470
rect 8588 20398 8616 21082
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8496 19446 8524 19722
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 14618 7788 17682
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7760 14006 7788 14554
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7852 13530 7880 15982
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8312 14958 8340 15846
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 8300 12912 8352 12918
rect 7746 12880 7802 12889
rect 8300 12854 8352 12860
rect 7746 12815 7802 12824
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7116 9926 7144 10678
rect 7300 10606 7328 11630
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4448 800 4476 3470
rect 4816 800 4844 3470
rect 5276 2990 5304 7754
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 3942 5396 4490
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5184 800 5212 2926
rect 5460 2446 5488 6802
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5552 800 5580 2450
rect 5920 800 5948 4082
rect 6748 3738 6776 7482
rect 7116 4622 7144 9862
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6276 2372 6328 2378
rect 6276 2314 6328 2320
rect 6288 800 6316 2314
rect 6656 800 6684 3470
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7024 800 7052 2994
rect 7668 2514 7696 8502
rect 7760 3738 7788 12815
rect 8312 12442 8340 12854
rect 8404 12782 8432 18906
rect 8496 18766 8524 19382
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 18358 8524 18702
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8496 16794 8524 18294
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8588 15910 8616 19178
rect 8680 17202 8708 23734
rect 8772 19514 8800 30670
rect 8864 30122 8892 42638
rect 8956 34202 8984 44270
rect 9416 42158 9444 44882
rect 9600 44538 9628 50254
rect 10140 49156 10192 49162
rect 10140 49098 10192 49104
rect 9956 48816 10008 48822
rect 9956 48758 10008 48764
rect 9772 46708 9824 46714
rect 9772 46650 9824 46656
rect 9680 44804 9732 44810
rect 9680 44746 9732 44752
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 9692 42362 9720 44746
rect 9784 42770 9812 46650
rect 9968 44946 9996 48758
rect 9956 44940 10008 44946
rect 9956 44882 10008 44888
rect 10152 42770 10180 49098
rect 10232 47660 10284 47666
rect 10232 47602 10284 47608
rect 10244 46578 10272 47602
rect 10232 46572 10284 46578
rect 10232 46514 10284 46520
rect 10244 44402 10272 46514
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 44742 10456 46310
rect 10520 45558 10548 51342
rect 10600 51332 10652 51338
rect 10600 51274 10652 51280
rect 10612 46714 10640 51274
rect 10704 49366 10732 53518
rect 11716 49366 11744 54130
rect 12360 54126 12388 56222
rect 13450 56200 13506 57000
rect 13556 56222 13768 56250
rect 13464 56114 13492 56200
rect 13556 56114 13584 56222
rect 13464 56086 13584 56114
rect 13740 54194 13768 56222
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 13728 54188 13780 54194
rect 13728 54130 13780 54136
rect 14832 54188 14884 54194
rect 16500 54176 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 20456 56222 20668 56250
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18604 54324 18656 54330
rect 18604 54266 18656 54272
rect 16580 54188 16632 54194
rect 16500 54148 16580 54176
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 17592 54130 17644 54136
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 15844 54052 15896 54058
rect 15844 53994 15896 54000
rect 12440 53984 12492 53990
rect 12440 53926 12492 53932
rect 14924 53984 14976 53990
rect 14924 53926 14976 53932
rect 10692 49360 10744 49366
rect 10692 49302 10744 49308
rect 11704 49360 11756 49366
rect 11704 49302 11756 49308
rect 10876 49156 10928 49162
rect 10876 49098 10928 49104
rect 10600 46708 10652 46714
rect 10600 46650 10652 46656
rect 10612 45966 10640 46650
rect 10600 45960 10652 45966
rect 10600 45902 10652 45908
rect 10508 45552 10560 45558
rect 10508 45494 10560 45500
rect 10416 44736 10468 44742
rect 10416 44678 10468 44684
rect 10232 44396 10284 44402
rect 10232 44338 10284 44344
rect 10520 44266 10548 45494
rect 10784 44804 10836 44810
rect 10784 44746 10836 44752
rect 10508 44260 10560 44266
rect 10508 44202 10560 44208
rect 10692 44192 10744 44198
rect 10692 44134 10744 44140
rect 9772 42764 9824 42770
rect 9772 42706 9824 42712
rect 10140 42764 10192 42770
rect 10140 42706 10192 42712
rect 9680 42356 9732 42362
rect 9680 42298 9732 42304
rect 10704 42158 10732 44134
rect 10796 42226 10824 44746
rect 10784 42220 10836 42226
rect 10784 42162 10836 42168
rect 9404 42152 9456 42158
rect 9404 42094 9456 42100
rect 9680 42152 9732 42158
rect 9680 42094 9732 42100
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 9220 41608 9272 41614
rect 9220 41550 9272 41556
rect 8944 34196 8996 34202
rect 8944 34138 8996 34144
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 8852 30116 8904 30122
rect 8852 30058 8904 30064
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8864 16454 8892 22986
rect 8956 17134 8984 25910
rect 9048 23322 9076 33934
rect 9232 30938 9260 41550
rect 9416 35630 9444 42094
rect 9496 37868 9548 37874
rect 9496 37810 9548 37816
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9416 34066 9444 35566
rect 9404 34060 9456 34066
rect 9404 34002 9456 34008
rect 9220 30932 9272 30938
rect 9220 30874 9272 30880
rect 9508 29306 9536 37810
rect 9692 35834 9720 42094
rect 9680 35828 9732 35834
rect 9680 35770 9732 35776
rect 10796 35698 10824 42162
rect 10888 41818 10916 49098
rect 12348 48000 12400 48006
rect 12348 47942 12400 47948
rect 12360 46646 12388 47942
rect 12348 46640 12400 46646
rect 12348 46582 12400 46588
rect 12452 46510 12480 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 14936 47122 14964 53926
rect 14924 47116 14976 47122
rect 14924 47058 14976 47064
rect 12440 46504 12492 46510
rect 12440 46446 12492 46452
rect 13728 46504 13780 46510
rect 13728 46446 13780 46452
rect 14648 46504 14700 46510
rect 14648 46446 14700 46452
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12808 45960 12860 45966
rect 12808 45902 12860 45908
rect 12820 45558 12848 45902
rect 12808 45552 12860 45558
rect 12808 45494 12860 45500
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10980 41682 11008 44134
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9692 29102 9720 35566
rect 10796 30054 10824 35634
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12808 32360 12860 32366
rect 12808 32302 12860 32308
rect 12820 31278 12848 32302
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12820 30394 12848 31214
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 13740 30190 13768 46446
rect 14660 46170 14688 46446
rect 14648 46164 14700 46170
rect 14648 46106 14700 46112
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 14648 33924 14700 33930
rect 14648 33866 14700 33872
rect 14660 32842 14688 33866
rect 14648 32836 14700 32842
rect 14648 32778 14700 32784
rect 14660 32502 14688 32778
rect 14280 32496 14332 32502
rect 14280 32438 14332 32444
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14096 31952 14148 31958
rect 14096 31894 14148 31900
rect 13912 30660 13964 30666
rect 13912 30602 13964 30608
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 10784 30048 10836 30054
rect 10784 29990 10836 29996
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 11612 29844 11664 29850
rect 11612 29786 11664 29792
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9956 28484 10008 28490
rect 9956 28426 10008 28432
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9220 27532 9272 27538
rect 9220 27474 9272 27480
rect 9232 26994 9260 27474
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9128 25900 9180 25906
rect 9232 25888 9260 26930
rect 9416 25974 9444 27950
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9180 25860 9260 25888
rect 9128 25842 9180 25848
rect 9692 25362 9720 28426
rect 9968 27334 9996 28426
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 9968 27062 9996 27270
rect 9956 27056 10008 27062
rect 9956 26998 10008 27004
rect 9968 26738 9996 26998
rect 10048 26920 10100 26926
rect 10048 26862 10100 26868
rect 9876 26710 9996 26738
rect 9876 26314 9904 26710
rect 10060 26586 10088 26862
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9876 25974 9904 26250
rect 9864 25968 9916 25974
rect 9864 25910 9916 25916
rect 9680 25356 9732 25362
rect 9732 25316 9812 25344
rect 9680 25298 9732 25304
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9324 24274 9352 24686
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23798 9168 24006
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9220 23248 9272 23254
rect 9220 23190 9272 23196
rect 9232 20058 9260 23190
rect 9508 23118 9536 23734
rect 9692 23526 9720 24686
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9034 18184 9090 18193
rect 9034 18119 9090 18128
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 9048 16946 9076 18119
rect 8956 16918 9076 16946
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8956 14226 8984 16918
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9048 16590 9076 16730
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9140 15706 9168 19314
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18358 9260 19110
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8772 14198 8984 14226
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8496 13870 8524 13942
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12436 8352 12442
rect 8496 12434 8524 13806
rect 8496 12406 8616 12434
rect 8300 12378 8352 12384
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8588 11762 8616 12406
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 10130 8248 10542
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7392 800 7420 2382
rect 7760 800 7788 2382
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 2994
rect 8772 1902 8800 14198
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8864 6866 8892 14010
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8864 800 8892 2994
rect 8956 2774 8984 10542
rect 9048 9994 9076 14826
rect 9232 13530 9260 17546
rect 9324 17338 9352 21422
rect 9508 20602 9536 22918
rect 9784 22574 9812 25316
rect 9876 24886 9904 25910
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9876 24138 9904 24822
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23866 9904 24074
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9600 20466 9628 20946
rect 9876 20942 9904 21966
rect 10060 21010 10088 26522
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10152 21690 10180 21966
rect 10244 21690 10272 29106
rect 10336 25498 10364 29174
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10888 28762 10916 29038
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 10428 26450 10456 28562
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10692 26852 10744 26858
rect 10692 26794 10744 26800
rect 10704 26450 10732 26794
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10796 26042 10824 27338
rect 11072 27130 11100 29514
rect 11440 28626 11468 29650
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11624 28490 11652 29786
rect 12544 29646 12572 29990
rect 12728 29782 12756 30126
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13464 29850 13492 29990
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 12716 29776 12768 29782
rect 12716 29718 12768 29724
rect 13924 29714 13952 30602
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 13924 29238 13952 29650
rect 13912 29232 13964 29238
rect 13912 29174 13964 29180
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10784 26036 10836 26042
rect 10836 25996 10916 26024
rect 10784 25978 10836 25984
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9600 18426 9628 20402
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9600 18306 9628 18362
rect 9508 18278 9628 18306
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9416 17338 9444 17614
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 13530 9352 14418
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9140 11150 9168 13262
rect 9324 12434 9352 13466
rect 9416 12850 9444 17070
rect 9508 16658 9536 18278
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9600 17678 9628 18090
rect 9692 17746 9720 20334
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 17270 9628 17614
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9784 16250 9812 20470
rect 9968 18766 9996 20742
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9968 16574 9996 17478
rect 10060 16946 10088 19314
rect 10336 18426 10364 22918
rect 10428 22506 10456 25638
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10428 18902 10456 22442
rect 10520 22234 10548 23462
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10152 17082 10180 18226
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17202 10272 17478
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10152 17054 10272 17082
rect 10060 16918 10180 16946
rect 9968 16546 10088 16574
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15570 9628 15982
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15450 9628 15506
rect 9600 15422 9720 15450
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9508 12918 9536 15302
rect 9600 12986 9628 15302
rect 9692 15094 9720 15422
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14414 9996 14758
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 14006 9812 14214
rect 9968 14006 9996 14350
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9232 12406 9352 12434
rect 9232 12306 9260 12406
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9232 11898 9260 12242
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 9140 9042 9168 11086
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9416 3670 9444 12786
rect 9784 12782 9812 13126
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9600 7206 9628 10066
rect 9692 8906 9720 10950
rect 9784 10810 9812 12718
rect 9876 11898 9904 13398
rect 10060 12442 10088 16546
rect 10152 15162 10180 16918
rect 10244 16574 10272 17054
rect 10244 16546 10364 16574
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10152 11762 10180 12310
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9876 10742 9904 11698
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 5710 9628 7142
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 4690 9628 5646
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 2854 9168 3334
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8956 2746 9076 2774
rect 9048 2650 9076 2746
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9232 800 9260 2994
rect 9600 800 9628 3470
rect 9692 3194 9720 6598
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9784 2854 9812 9658
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 3466 10088 7686
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10152 2990 10180 11698
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 10244 2582 10272 15302
rect 10336 12714 10364 16546
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10428 12434 10456 18702
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 18426 10548 18566
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10336 12406 10456 12434
rect 10336 7750 10364 12406
rect 10520 12374 10548 16186
rect 10612 16114 10640 22102
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10704 19922 10732 20878
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10796 18970 10824 25162
rect 10888 24682 10916 25996
rect 11072 25838 11100 27066
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 10980 25294 11008 25706
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 11164 24614 11192 25434
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 21486 11008 22510
rect 11072 22030 11100 23122
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21554 11100 21830
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 11164 21350 11192 24550
rect 11624 22166 11652 28426
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11796 26512 11848 26518
rect 11796 26454 11848 26460
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11716 23118 11744 25094
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11808 23050 11836 26454
rect 11992 25226 12020 26726
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 10888 19718 10916 20810
rect 11440 20534 11468 20810
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11440 19786 11468 20470
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10888 18834 10916 19654
rect 11440 19514 11468 19722
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11624 19122 11652 21558
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19378 11744 19654
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11624 19094 11744 19122
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10796 18086 10824 18294
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15366 10640 16050
rect 10796 16046 10824 18022
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12714 10640 13194
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10888 12434 10916 18566
rect 11624 17746 11652 18838
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 13870 11008 17478
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 12986 11100 13670
rect 11164 13530 11192 16390
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11256 13802 11284 14282
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11256 13258 11284 13738
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10704 12406 10916 12434
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10704 12186 10732 12406
rect 10428 12158 10732 12186
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10428 5302 10456 12158
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10612 11354 10640 12038
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11144 10560 11150
rect 10560 11092 10640 11098
rect 10508 11086 10640 11092
rect 10520 11070 10640 11086
rect 10612 10742 10640 11070
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10612 9994 10640 10678
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10612 9654 10640 9930
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10612 8922 10640 9590
rect 10704 9110 10732 12038
rect 10980 11626 11008 12718
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 11072 11150 11100 11630
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10198 10916 10950
rect 11072 10266 11100 11086
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 11164 9994 11192 10406
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10612 8906 10732 8922
rect 10612 8900 10744 8906
rect 10612 8894 10692 8900
rect 10692 8842 10744 8848
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9876 2038 9904 2382
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9864 2032 9916 2038
rect 9864 1974 9916 1980
rect 9968 800 9996 2314
rect 10336 800 10364 2994
rect 10520 2310 10548 7686
rect 10704 7410 10732 8842
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 6730 10732 7346
rect 10796 6798 10824 8978
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 7954 10916 8774
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10888 7342 10916 7890
rect 10980 7546 11008 7890
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 5642 10732 6666
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10704 4554 10732 5578
rect 10796 5166 10824 6734
rect 10980 5778 11008 7482
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11072 6866 11100 7278
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10704 800 10732 3470
rect 10968 3188 11020 3194
rect 11164 3176 11192 8298
rect 11348 7818 11376 15574
rect 11440 12442 11468 16458
rect 11624 15910 11652 17138
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11716 15706 11744 19094
rect 11808 17338 11836 21558
rect 11992 19922 12020 25162
rect 12084 22778 12112 26386
rect 12176 24818 12204 27814
rect 12452 27334 12480 28562
rect 12716 28484 12768 28490
rect 12716 28426 12768 28432
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12452 26858 12480 27270
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12544 26042 12572 27270
rect 12728 26246 12756 28426
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 13096 27130 13124 27474
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12268 22098 12296 23462
rect 12360 22642 12388 24210
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21690 12296 21830
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12360 21554 12388 22578
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11900 16250 11928 19654
rect 12176 16250 12204 21354
rect 12452 21146 12480 25842
rect 12728 25226 12756 26182
rect 12820 25362 12848 26930
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13556 26586 13584 27474
rect 13648 27062 13676 29038
rect 13820 28688 13872 28694
rect 13820 28630 13872 28636
rect 13832 27402 13860 28630
rect 14108 28218 14136 31894
rect 14292 30734 14320 32438
rect 15672 31754 15700 37266
rect 15396 31726 15700 31754
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14292 30326 14320 30670
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14200 28422 14228 28902
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13832 26246 13860 26998
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13636 25832 13688 25838
rect 13464 25780 13636 25786
rect 13464 25774 13688 25780
rect 13464 25758 13676 25774
rect 13464 25702 13492 25758
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13360 25424 13412 25430
rect 13360 25366 13412 25372
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12728 24886 12756 25162
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 23798 12664 24006
rect 12624 23792 12676 23798
rect 12624 23734 12676 23740
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12268 16046 12296 17682
rect 12452 17338 12480 18702
rect 12544 18698 12572 22918
rect 12728 22710 12756 24822
rect 12820 24818 12848 25298
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 13372 24750 13400 25366
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13372 23594 13400 24686
rect 13360 23588 13412 23594
rect 13360 23530 13412 23536
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13360 23248 13412 23254
rect 13360 23190 13412 23196
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12636 21010 12664 22646
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 21962 12756 22510
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 17882 12572 18226
rect 12636 17882 12664 20946
rect 12728 20466 12756 21490
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 19922 12756 20402
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19446 12756 19858
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 16574 12572 17818
rect 12728 17746 12756 19382
rect 12820 18358 12848 23054
rect 13372 22982 13400 23190
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13464 22778 13492 25298
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13740 24614 13768 25230
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13740 23526 13768 23598
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13832 22030 13860 25842
rect 14200 25838 14228 28358
rect 14568 28150 14596 31146
rect 14936 30258 14964 31350
rect 15016 31136 15068 31142
rect 15016 31078 15068 31084
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14936 29238 14964 30194
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 14936 29034 14964 29174
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14924 28416 14976 28422
rect 14924 28358 14976 28364
rect 14556 28144 14608 28150
rect 14556 28086 14608 28092
rect 14752 27470 14780 28358
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14936 27402 14964 28358
rect 15028 28014 15056 31078
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 15120 28558 15148 30126
rect 15396 29510 15424 31726
rect 15856 31498 15884 53994
rect 16120 53984 16172 53990
rect 16120 53926 16172 53932
rect 17684 53984 17736 53990
rect 17684 53926 17736 53932
rect 15936 47592 15988 47598
rect 15936 47534 15988 47540
rect 15672 31470 15884 31498
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15580 29646 15608 30058
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 15212 29306 15240 29446
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 14280 27396 14332 27402
rect 14280 27338 14332 27344
rect 14924 27396 14976 27402
rect 14924 27338 14976 27344
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 20398 13400 21286
rect 13464 20806 13492 21558
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13464 20534 13492 20742
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17066 12664 17478
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12728 16794 12756 17682
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12544 16546 12756 16574
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10130 11468 10950
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11532 8566 11560 13738
rect 11624 9178 11652 14962
rect 11900 14482 11928 15982
rect 12268 15570 12296 15982
rect 12636 15706 12664 16050
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12728 15450 12756 16546
rect 12820 16522 12848 17750
rect 12912 17134 12940 17818
rect 13372 17134 13400 20334
rect 13924 20058 13952 23666
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22030 14136 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21486 14136 21966
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13556 16574 13584 17818
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 17338 13676 17614
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13372 16546 13584 16574
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12820 15570 12848 16458
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15609 13400 16546
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13358 15600 13414 15609
rect 12808 15564 12860 15570
rect 13358 15535 13414 15544
rect 12808 15506 12860 15512
rect 12624 15428 12676 15434
rect 12728 15422 13400 15450
rect 12624 15370 12676 15376
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 12918 11928 13874
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11716 8634 11744 12718
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11808 11082 11836 12310
rect 11992 11898 12020 15030
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13394 12112 14418
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12306 12112 13330
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11716 5914 11744 7278
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11808 4010 11836 11018
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 10062 12020 10406
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12084 9042 12112 11562
rect 12176 11218 12204 13126
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 12084 7750 12112 7958
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 12176 3534 12204 8570
rect 12268 4146 12296 14758
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 12850 12480 13670
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12360 10198 12388 12650
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 11898 12480 12582
rect 12544 12374 12572 13806
rect 12636 12442 12664 15370
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11020 3148 11192 3176
rect 10968 3130 11020 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10980 1970 11008 2314
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 11072 800 11100 2994
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11440 800 11468 2926
rect 11808 800 11836 2994
rect 12360 2582 12388 9318
rect 12452 6458 12480 11494
rect 12544 10810 12572 12106
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11014 12664 12038
rect 12728 11830 12756 14214
rect 12820 11898 12848 15302
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 14006 13308 14214
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12306 13400 15422
rect 13464 13326 13492 16390
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13556 14346 13584 16118
rect 13648 16046 13676 17138
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13648 15638 13676 15982
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13634 15464 13690 15473
rect 13634 15399 13690 15408
rect 13648 15042 13676 15399
rect 13740 15162 13768 19450
rect 14108 16794 14136 19450
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14200 17270 14228 18158
rect 14292 17882 14320 27338
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14832 26444 14884 26450
rect 14832 26386 14884 26392
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14752 24614 14780 26318
rect 14844 25498 14872 26386
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14844 25362 14872 25434
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14844 25129 14872 25162
rect 14830 25120 14886 25129
rect 14830 25055 14886 25064
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14752 24410 14780 24550
rect 14740 24404 14792 24410
rect 14740 24346 14792 24352
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14384 20534 14412 20742
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19310 14504 20198
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13648 15014 13768 15042
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14482 13676 14826
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13450 13016 13506 13025
rect 13450 12951 13506 12960
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12912 11676 12940 12106
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 12728 11648 12940 11676
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12728 10826 12756 11648
rect 13280 11626 13308 11834
rect 13372 11830 13400 12242
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13464 11558 13492 12951
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 12820 11082 12848 11494
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12992 11348 13044 11354
rect 13556 11336 13584 14282
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13394 13676 13670
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 12992 11290 13044 11296
rect 13464 11308 13584 11336
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10798 12756 10826
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 8022 12572 9454
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 6866 12572 7958
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12452 3534 12480 4111
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12176 800 12204 2382
rect 12544 800 12572 3538
rect 12636 3194 12664 10798
rect 12820 10656 12848 11018
rect 12728 10628 12848 10656
rect 12728 8401 12756 10628
rect 13004 10452 13032 11290
rect 13464 10538 13492 11308
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 12820 10424 13032 10452
rect 13360 10464 13412 10470
rect 12714 8392 12770 8401
rect 12714 8327 12770 8336
rect 12820 8004 12848 10424
rect 13360 10406 13412 10412
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 10266 13400 10406
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13372 8838 13400 9046
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13464 8378 13492 10202
rect 13556 10130 13584 11154
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9042 13584 10066
rect 13648 9042 13676 13126
rect 13740 13025 13768 15014
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13462 13860 13806
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13726 13016 13782 13025
rect 13726 12951 13782 12960
rect 13832 12918 13860 13398
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12170 13768 12786
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 11694 13768 11766
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11354 13768 11494
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10810 13768 10950
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13634 8936 13690 8945
rect 13634 8871 13690 8880
rect 13464 8350 13584 8378
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12820 7976 12940 8004
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 2854 12756 7754
rect 12912 7750 12940 7976
rect 13372 7886 13400 8230
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12820 6322 12848 7686
rect 13464 7410 13492 8230
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6390 13308 6598
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13372 5302 13400 6802
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12820 1714 12848 3538
rect 13174 3088 13230 3097
rect 13174 3023 13176 3032
rect 13228 3023 13230 3032
rect 13176 2994 13228 3000
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12898 2544 12954 2553
rect 12898 2479 12954 2488
rect 12912 2446 12940 2479
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13464 2310 13492 6190
rect 13556 5710 13584 8350
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13648 4690 13676 8871
rect 13740 8090 13768 9998
rect 13832 8566 13860 12718
rect 13924 12714 13952 12854
rect 14016 12782 14044 13126
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 14108 12434 14136 14894
rect 14016 12406 14136 12434
rect 14016 10742 14044 12406
rect 14200 11898 14228 15642
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 12782 14320 13670
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 8560 13872 8566
rect 13924 8537 13952 10542
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8974 14044 9318
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14108 8634 14136 11698
rect 14292 9518 14320 12718
rect 14384 12442 14412 16186
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14476 15162 14504 15438
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14476 12170 14504 13262
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 12374 14596 13194
rect 14660 13190 14688 21354
rect 14752 20602 14780 23258
rect 14844 21978 14872 24686
rect 14936 23866 14964 26726
rect 15028 26382 15056 27474
rect 15120 27130 15148 28494
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 15120 26246 15148 26930
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 23866 15148 26182
rect 15212 26042 15240 28970
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24886 15240 25094
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15120 23254 15148 23802
rect 15304 23526 15332 27270
rect 15396 25158 15424 29446
rect 15580 26364 15608 29582
rect 15672 28422 15700 31470
rect 15844 31340 15896 31346
rect 15948 31328 15976 47534
rect 16132 46646 16160 53926
rect 17592 50720 17644 50726
rect 17592 50662 17644 50668
rect 16120 46640 16172 46646
rect 16120 46582 16172 46588
rect 16396 46504 16448 46510
rect 16396 46446 16448 46452
rect 16304 42084 16356 42090
rect 16304 42026 16356 42032
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31414 16160 31826
rect 16120 31408 16172 31414
rect 16120 31350 16172 31356
rect 15896 31300 15976 31328
rect 16028 31340 16080 31346
rect 15844 31282 15896 31288
rect 16028 31282 16080 31288
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15660 28416 15712 28422
rect 15660 28358 15712 28364
rect 15764 27062 15792 28970
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15488 26336 15608 26364
rect 15488 25226 15516 26336
rect 15856 26314 15884 31282
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15948 29238 15976 31078
rect 16040 30394 16068 31282
rect 16212 31272 16264 31278
rect 16212 31214 16264 31220
rect 16028 30388 16080 30394
rect 16028 30330 16080 30336
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15948 27334 15976 28358
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 14844 21950 14964 21978
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21622 14872 21830
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14936 21486 14964 21950
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 14936 19514 14964 19858
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15120 18154 15148 19314
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15212 17542 15240 21830
rect 15488 20602 15516 24550
rect 15580 23798 15608 26182
rect 15948 25158 15976 27270
rect 16040 26994 16068 30330
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16132 29102 16160 29990
rect 16224 29714 16252 31214
rect 16212 29708 16264 29714
rect 16212 29650 16264 29656
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16120 29096 16172 29102
rect 16120 29038 16172 29044
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15764 22166 15792 25094
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15856 23118 15884 23462
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15396 16998 15424 20402
rect 15764 20058 15792 20810
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15948 19718 15976 23734
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16040 21010 16068 21966
rect 16224 21554 16252 29242
rect 16316 28422 16344 42026
rect 16408 35698 16436 46446
rect 17500 45892 17552 45898
rect 17500 45834 17552 45840
rect 17224 44192 17276 44198
rect 17224 44134 17276 44140
rect 16396 35692 16448 35698
rect 16396 35634 16448 35640
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16684 31822 16712 33050
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16776 31890 16804 32302
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16684 29102 16712 31758
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17144 31210 17172 31622
rect 17236 31346 17264 44134
rect 17512 35086 17540 45834
rect 17500 35080 17552 35086
rect 17500 35022 17552 35028
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17132 31204 17184 31210
rect 17132 31146 17184 31152
rect 17144 29102 17172 31146
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 16304 28416 16356 28422
rect 16304 28358 16356 28364
rect 16396 28416 16448 28422
rect 16396 28358 16448 28364
rect 16316 26246 16344 28358
rect 16408 26518 16436 28358
rect 16580 28076 16632 28082
rect 16580 28018 16632 28024
rect 16396 26512 16448 26518
rect 16396 26454 16448 26460
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14752 12434 14780 16662
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16250 14872 16458
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 14278 14964 16050
rect 15120 16046 15148 16730
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 15212 13938 15240 15506
rect 15488 14482 15516 17070
rect 15672 16574 15700 18566
rect 15948 17066 15976 19654
rect 16132 19310 16160 19994
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16224 18850 16252 21082
rect 16316 19446 16344 23462
rect 16408 23322 16436 26454
rect 16592 25226 16620 28018
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27130 16896 27814
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16776 25945 16804 25978
rect 16762 25936 16818 25945
rect 16762 25871 16818 25880
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 16776 25362 16804 25638
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16592 24886 16620 25162
rect 16580 24880 16632 24886
rect 16580 24822 16632 24828
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16592 22982 16620 23190
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16224 18822 16344 18850
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15948 16946 15976 17002
rect 15580 16546 15700 16574
rect 15764 16918 15976 16946
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14936 12782 14964 13466
rect 15396 13394 15424 14418
rect 15488 13870 15516 14418
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15014 13016 15070 13025
rect 15014 12951 15016 12960
rect 15068 12951 15070 12960
rect 15016 12922 15068 12928
rect 15108 12912 15160 12918
rect 15106 12880 15108 12889
rect 15160 12880 15162 12889
rect 15106 12815 15162 12824
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14660 12406 14780 12434
rect 14832 12436 14884 12442
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14476 9518 14504 12106
rect 14660 12102 14688 12406
rect 14832 12378 14884 12384
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 10266 14596 11562
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14660 10146 14688 12038
rect 14844 11898 14872 12378
rect 14832 11892 14884 11898
rect 14568 10118 14688 10146
rect 14752 11852 14832 11880
rect 14568 9654 14596 10118
rect 14752 10044 14780 11852
rect 14832 11834 14884 11840
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 10606 14872 11630
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14936 10130 14964 12718
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11082 15056 12038
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14660 10016 14780 10044
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9330 14504 9454
rect 14384 9302 14504 9330
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13820 8502 13872 8508
rect 13910 8528 13966 8537
rect 13910 8463 13966 8472
rect 13818 8392 13874 8401
rect 13818 8327 13874 8336
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13832 7970 13860 8327
rect 13740 7942 13860 7970
rect 13740 6798 13768 7942
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13740 3398 13768 6394
rect 13832 6322 13860 6938
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13924 6202 13952 8463
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13832 6174 13952 6202
rect 13832 3738 13860 6174
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13924 4146 13952 4966
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13648 800 13676 2926
rect 14016 800 14044 3538
rect 14108 3058 14136 8298
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7478 14320 7754
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2446 14228 5510
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14292 2378 14320 5510
rect 14384 3126 14412 9302
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8634 14504 8842
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14464 7880 14516 7886
rect 14462 7848 14464 7857
rect 14516 7848 14518 7857
rect 14462 7783 14518 7792
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5710 14504 6054
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 3534 14504 4966
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14568 3466 14596 9590
rect 14660 8838 14688 10016
rect 14832 9920 14884 9926
rect 14936 9874 14964 10066
rect 14884 9868 14964 9874
rect 14832 9862 14964 9868
rect 14844 9846 14964 9862
rect 14936 9518 14964 9846
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14752 8498 14780 9318
rect 14936 9042 14964 9454
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 7886 14688 8298
rect 14844 8265 14872 8434
rect 14830 8256 14886 8265
rect 14830 8191 14886 8200
rect 15028 7886 15056 11018
rect 15120 10810 15148 12310
rect 15212 11354 15240 13126
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7546 14780 7686
rect 15120 7562 15148 9862
rect 15212 9450 15240 10950
rect 15304 9994 15332 11766
rect 15488 10198 15516 13466
rect 15580 10674 15608 16546
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 16114 15700 16390
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15764 14958 15792 16918
rect 16040 16590 16068 17070
rect 16132 16590 16160 17614
rect 16316 16658 16344 18822
rect 16500 18290 16528 20946
rect 16592 20942 16620 21898
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16592 20534 16620 20878
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16592 19786 16620 20470
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16684 18970 16712 19790
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16776 18714 16804 19450
rect 16868 19446 16896 26250
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 16856 19440 16908 19446
rect 16856 19382 16908 19388
rect 16868 18766 16896 19382
rect 16684 18686 16804 18714
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 17218 16436 18158
rect 16500 17338 16528 18226
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16408 17190 16528 17218
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 15162 15884 15438
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15672 13190 15700 13398
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15658 13016 15714 13025
rect 15658 12951 15660 12960
rect 15712 12951 15714 12960
rect 15660 12922 15712 12928
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9722 15332 9930
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14936 7534 15148 7562
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5370 14872 6190
rect 14936 5778 14964 7534
rect 15580 7478 15608 10610
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15028 5574 15056 7414
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6934 15148 7142
rect 15672 7018 15700 10950
rect 15764 9518 15792 13330
rect 16040 12889 16068 14894
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16026 12880 16082 12889
rect 16026 12815 16082 12824
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16040 12434 16068 12718
rect 15856 12406 16068 12434
rect 15856 10606 15884 12406
rect 16132 11150 16160 13874
rect 16224 13462 16252 16594
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16316 12434 16344 15846
rect 16408 14822 16436 16934
rect 16500 14958 16528 17190
rect 16592 16658 16620 17274
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 15570 16620 16594
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16224 12406 16344 12434
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15936 10736 15988 10742
rect 15934 10704 15936 10713
rect 15988 10704 15990 10713
rect 16224 10690 16252 12406
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16316 11286 16344 11630
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 15934 10639 15990 10648
rect 16040 10662 16252 10690
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7546 15792 7822
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15396 6990 15700 7018
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15212 6458 15240 6598
rect 15304 6458 15332 6734
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14844 4078 14872 5306
rect 15028 5302 15056 5510
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 15028 4486 15056 5238
rect 15396 4554 15424 6990
rect 15566 6896 15622 6905
rect 15476 6860 15528 6866
rect 15764 6882 15792 7346
rect 15622 6854 15792 6882
rect 15566 6831 15622 6840
rect 15476 6802 15528 6808
rect 15488 4554 15516 6802
rect 15580 6662 15608 6831
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 4826 15700 6258
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15016 4480 15068 4486
rect 14936 4428 15016 4434
rect 14936 4422 15068 4428
rect 14936 4406 15056 4422
rect 14936 4214 14964 4406
rect 15488 4282 15516 4490
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 15856 3670 15884 10542
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8838 15976 8910
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16040 6746 16068 10662
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 9042 16160 10542
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 15948 6718 16068 6746
rect 15948 5030 15976 6718
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 800 15148 2790
rect 15488 800 15516 3538
rect 16040 3194 16068 6598
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 4010 16160 5646
rect 16224 4826 16252 7890
rect 16316 7342 16344 11222
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15856 800 15884 2926
rect 16224 800 16252 4014
rect 16316 3738 16344 4082
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16408 3534 16436 10406
rect 16500 9926 16528 14486
rect 16684 14362 16712 18686
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 14498 16804 18566
rect 16960 17678 16988 25638
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 17052 22098 17080 24618
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21146 17080 22034
rect 17144 21978 17172 29038
rect 17236 28082 17264 31282
rect 17316 31272 17368 31278
rect 17316 31214 17368 31220
rect 17328 30954 17356 31214
rect 17328 30938 17448 30954
rect 17328 30932 17460 30938
rect 17328 30926 17408 30932
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17328 28014 17356 30926
rect 17408 30874 17460 30880
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17420 28014 17448 29038
rect 17604 28370 17632 50662
rect 17696 46034 17724 53926
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17684 46028 17736 46034
rect 17684 45970 17736 45976
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17684 44260 17736 44266
rect 17684 44202 17736 44208
rect 17512 28342 17632 28370
rect 17316 28008 17368 28014
rect 17314 27976 17316 27985
rect 17408 28008 17460 28014
rect 17368 27976 17370 27985
rect 17408 27950 17460 27956
rect 17314 27911 17370 27920
rect 17512 27402 17540 28342
rect 17696 28234 17724 44202
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 18616 37330 18644 54266
rect 18984 54194 19012 56200
rect 20364 56114 20392 56200
rect 20456 56114 20484 56222
rect 20364 56086 20484 56114
rect 20640 54194 20668 56222
rect 21730 56200 21786 57000
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 21744 54194 21772 56200
rect 23124 54194 23152 56200
rect 23294 56128 23350 56137
rect 23294 56063 23350 56072
rect 18972 54188 19024 54194
rect 18972 54130 19024 54136
rect 20628 54188 20680 54194
rect 20628 54130 20680 54136
rect 21732 54188 21784 54194
rect 21732 54130 21784 54136
rect 23112 54188 23164 54194
rect 23112 54130 23164 54136
rect 20904 53984 20956 53990
rect 20904 53926 20956 53932
rect 19984 52896 20036 52902
rect 19984 52838 20036 52844
rect 19800 49768 19852 49774
rect 19800 49710 19852 49716
rect 19524 43784 19576 43790
rect 19524 43726 19576 43732
rect 18604 37324 18656 37330
rect 18604 37266 18656 37272
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 19536 34048 19564 43726
rect 19708 34060 19760 34066
rect 19536 34020 19708 34048
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 19444 32910 19472 33934
rect 19536 33522 19564 34020
rect 19708 34002 19760 34008
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18328 32496 18380 32502
rect 18328 32438 18380 32444
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 18248 32026 18276 32302
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18340 31754 18368 32438
rect 19444 32434 19472 32846
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18340 30666 18368 31690
rect 18432 31278 18460 31826
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18328 30660 18380 30666
rect 18328 30602 18380 30608
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 17868 29708 17920 29714
rect 17868 29650 17920 29656
rect 17776 29028 17828 29034
rect 17776 28970 17828 28976
rect 17604 28206 17724 28234
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17236 24954 17264 26182
rect 17604 26042 17632 28206
rect 17684 28144 17736 28150
rect 17684 28086 17736 28092
rect 17592 26036 17644 26042
rect 17592 25978 17644 25984
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17236 23662 17264 24550
rect 17696 24206 17724 28086
rect 17788 24614 17816 28970
rect 17880 26976 17908 29650
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17960 26988 18012 26994
rect 17880 26948 17960 26976
rect 17960 26930 18012 26936
rect 17972 26450 18000 26930
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 25974 18368 29718
rect 18524 28218 18552 31078
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18432 27674 18460 28018
rect 18616 28014 18644 31962
rect 19076 31958 19104 32166
rect 19064 31952 19116 31958
rect 19064 31894 19116 31900
rect 19444 31890 19472 32370
rect 19708 32020 19760 32026
rect 19708 31962 19760 31968
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 19444 30802 19472 31826
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 18696 30660 18748 30666
rect 18696 30602 18748 30608
rect 18708 29714 18736 30602
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18800 29850 18828 30534
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18708 28966 18736 29650
rect 18696 28960 18748 28966
rect 18696 28902 18748 28908
rect 18708 28490 18736 28902
rect 18696 28484 18748 28490
rect 18696 28426 18748 28432
rect 18604 28008 18656 28014
rect 18800 27962 18828 29786
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18892 28762 18920 29582
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18604 27950 18656 27956
rect 18708 27934 18828 27962
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18604 26784 18656 26790
rect 18604 26726 18656 26732
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18432 26042 18460 26318
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18524 24818 18552 25162
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17236 23050 17264 23598
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17236 22710 17264 22986
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17144 21950 17264 21978
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17144 20534 17172 21830
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17144 19922 17172 20470
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 18358 17080 19722
rect 17236 18834 17264 21950
rect 17328 19514 17356 23258
rect 17592 23248 17644 23254
rect 17592 23190 17644 23196
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 17420 20346 17448 20470
rect 17500 20392 17552 20398
rect 17420 20340 17500 20346
rect 17420 20334 17552 20340
rect 17420 20318 17540 20334
rect 17420 19786 17448 20318
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17328 19417 17356 19450
rect 17314 19408 17370 19417
rect 17314 19343 17370 19352
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17040 18352 17092 18358
rect 17236 18329 17264 18362
rect 17040 18294 17092 18300
rect 17222 18320 17278 18329
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16946 17504 17002 17513
rect 16868 16574 16896 17478
rect 16946 17439 17002 17448
rect 16960 17270 16988 17439
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 17052 17202 17080 18294
rect 17222 18255 17278 18264
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16794 17080 17138
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17144 16697 17172 17002
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 16868 16546 17080 16574
rect 16776 14470 16988 14498
rect 16684 14334 16804 14362
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16500 8090 16528 9114
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16500 2582 16528 7142
rect 16592 4146 16620 13126
rect 16684 12986 16712 14214
rect 16776 12986 16804 14334
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16762 12744 16818 12753
rect 16762 12679 16764 12688
rect 16816 12679 16818 12688
rect 16764 12650 16816 12656
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16684 11898 16712 12310
rect 16868 12170 16896 13806
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16868 11218 16896 12106
rect 16960 11898 16988 14470
rect 17052 12374 17080 16546
rect 17236 16522 17264 17546
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17328 15994 17356 19178
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 17082 17540 18702
rect 17420 17054 17540 17082
rect 17420 16250 17448 17054
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17144 15966 17356 15994
rect 17144 13870 17172 15966
rect 17408 15904 17460 15910
rect 17236 15864 17408 15892
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16868 10538 16896 11154
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16684 8838 16712 9114
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 8430 16712 8774
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16592 800 16620 3062
rect 16776 2446 16804 9862
rect 16868 7342 16896 10474
rect 16946 10160 17002 10169
rect 16946 10095 17002 10104
rect 16960 8430 16988 10095
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 7818 16988 8366
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 17052 7478 17080 12174
rect 17144 9382 17172 13806
rect 17236 12434 17264 15864
rect 17408 15846 17460 15852
rect 17512 15586 17540 16730
rect 17604 16182 17632 23190
rect 17696 17610 17724 24142
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 19378 17816 20198
rect 17880 19854 17908 24550
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18248 23186 18276 23258
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 19922 18184 20334
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17788 16574 17816 18770
rect 17880 16590 17908 19654
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17972 16726 18000 16934
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17696 16546 17816 16574
rect 17868 16584 17920 16590
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17696 15638 17724 16546
rect 17868 16526 17920 16532
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17684 15632 17736 15638
rect 17512 15558 17632 15586
rect 17684 15574 17736 15580
rect 17604 15502 17632 15558
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13326 17356 13670
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17236 12406 17356 12434
rect 17328 12374 17356 12406
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17130 9072 17186 9081
rect 17130 9007 17186 9016
rect 17144 8974 17172 9007
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17130 8528 17186 8537
rect 17130 8463 17132 8472
rect 17184 8463 17186 8472
rect 17132 8434 17184 8440
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6254 16896 7278
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16868 5166 16896 6190
rect 17052 5302 17080 6802
rect 17144 6254 17172 8298
rect 17236 7834 17264 12310
rect 17420 12220 17448 12786
rect 17328 12192 17448 12220
rect 17328 10606 17356 12192
rect 17512 12102 17540 15302
rect 17604 14006 17632 15438
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17420 11354 17448 11766
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17328 9110 17356 9386
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17328 7954 17356 9046
rect 17420 8022 17448 11086
rect 17604 9994 17632 13806
rect 17788 13326 17816 16390
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17880 14550 17908 16186
rect 18340 16114 18368 24006
rect 18432 23322 18460 24686
rect 18616 24274 18644 26726
rect 18708 25838 18736 27934
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18432 17746 18460 22986
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18524 17270 18552 22918
rect 18616 20398 18644 23122
rect 18708 23050 18736 24890
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18616 18222 18644 20334
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17746 18644 18022
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18142 16008 18198 16017
rect 18142 15943 18144 15952
rect 18196 15943 18198 15952
rect 18144 15914 18196 15920
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18328 13728 18380 13734
rect 17866 13696 17922 13705
rect 18328 13670 18380 13676
rect 17866 13631 17922 13640
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17696 10810 17724 12310
rect 17788 12238 17816 13262
rect 17880 13258 17908 13631
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12918 18368 13670
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18326 12744 18382 12753
rect 18326 12679 18382 12688
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17512 9722 17540 9862
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17500 9512 17552 9518
rect 17498 9480 17500 9489
rect 17552 9480 17554 9489
rect 17498 9415 17554 9424
rect 17500 9376 17552 9382
rect 17498 9344 17500 9353
rect 17696 9364 17724 10746
rect 17788 9466 17816 11494
rect 18340 11218 18368 12679
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 17880 11082 18000 11098
rect 17880 11076 18012 11082
rect 17880 11070 17960 11076
rect 17880 10130 17908 11070
rect 17960 11018 18012 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18432 10690 18460 15846
rect 18616 15706 18644 17682
rect 18708 17270 18736 19382
rect 18800 18902 18828 27814
rect 18892 27130 18920 28426
rect 19076 27334 19104 28562
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 18880 27124 18932 27130
rect 18880 27066 18932 27072
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18892 24206 18920 25230
rect 19076 24274 19104 27270
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18694 16008 18750 16017
rect 18694 15943 18750 15952
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18708 15314 18736 15943
rect 18616 15286 18736 15314
rect 18616 13258 18644 15286
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18524 12186 18552 13194
rect 18708 13138 18736 14758
rect 18616 13110 18736 13138
rect 18616 12442 18644 13110
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18524 12158 18736 12186
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18156 10662 18460 10690
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17972 10010 18000 10202
rect 17880 9982 18000 10010
rect 17880 9654 17908 9982
rect 18064 9926 18092 10542
rect 18156 10044 18184 10662
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 10198 18460 10542
rect 18236 10192 18288 10198
rect 18234 10160 18236 10169
rect 18420 10192 18472 10198
rect 18288 10160 18290 10169
rect 18420 10134 18472 10140
rect 18234 10095 18290 10104
rect 18156 10016 18368 10044
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 18340 9489 18368 10016
rect 18326 9480 18382 9489
rect 17788 9438 17908 9466
rect 17552 9344 17554 9353
rect 17498 9279 17554 9288
rect 17604 9336 17724 9364
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17512 8498 17540 8978
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17236 7806 17448 7834
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4690 16896 5102
rect 17052 4826 17080 5238
rect 17144 5166 17172 6190
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 17236 4146 17264 7210
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 4026 17356 7686
rect 17420 6458 17448 7806
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17512 7410 17540 7686
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17604 5642 17632 9336
rect 17880 8922 17908 9438
rect 18326 9415 18382 9424
rect 17696 8894 17908 8922
rect 17696 8498 17724 8894
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 17144 3998 17356 4026
rect 16868 2922 16896 3946
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16960 800 16988 2858
rect 17144 2650 17172 3998
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17328 2514 17356 2790
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17512 2258 17540 4626
rect 17696 4010 17724 8434
rect 18340 8090 18368 9415
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4162 18368 7142
rect 18432 6390 18460 7414
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18432 5302 18460 6326
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18432 4554 18460 5238
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18340 4134 18460 4162
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18064 3738 18092 3878
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17328 2230 17540 2258
rect 17328 800 17356 2230
rect 17696 800 17724 3538
rect 18156 3534 18184 3878
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 4014
rect 18432 3058 18460 4134
rect 18524 3058 18552 12038
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 9654 18644 11086
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18616 6458 18644 7278
rect 18708 7206 18736 12158
rect 18800 10606 18828 18566
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18892 14890 18920 17546
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18984 14074 19012 17546
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18984 12782 19012 14010
rect 19076 13870 19104 20198
rect 19168 19854 19196 28970
rect 19260 20466 19288 29990
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 19444 29306 19472 29446
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19536 29170 19564 29446
rect 19720 29306 19748 31962
rect 19708 29300 19760 29306
rect 19708 29242 19760 29248
rect 19524 29164 19576 29170
rect 19524 29106 19576 29112
rect 19616 29164 19668 29170
rect 19616 29106 19668 29112
rect 19628 28762 19656 29106
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19444 26450 19472 28562
rect 19708 27328 19760 27334
rect 19708 27270 19760 27276
rect 19720 27130 19748 27270
rect 19708 27124 19760 27130
rect 19708 27066 19760 27072
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19444 24818 19472 26386
rect 19812 25294 19840 49710
rect 19996 42090 20024 52838
rect 20812 43716 20864 43722
rect 20812 43658 20864 43664
rect 19984 42084 20036 42090
rect 19984 42026 20036 42032
rect 20260 35828 20312 35834
rect 20260 35770 20312 35776
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 19904 29714 19932 35430
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19996 33318 20024 33866
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 20168 30728 20220 30734
rect 20168 30670 20220 30676
rect 20180 30326 20208 30670
rect 20272 30326 20300 35770
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20352 32836 20404 32842
rect 20352 32778 20404 32784
rect 20364 32366 20392 32778
rect 20352 32360 20404 32366
rect 20352 32302 20404 32308
rect 20168 30320 20220 30326
rect 20168 30262 20220 30268
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 20364 29170 20392 32302
rect 20456 30190 20484 33254
rect 20548 31414 20576 35022
rect 20824 33998 20852 43658
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20824 33590 20852 33934
rect 20812 33584 20864 33590
rect 20812 33526 20864 33532
rect 20824 32502 20852 33526
rect 20916 33114 20944 53926
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53582 23336 56063
rect 23386 55448 23442 55457
rect 23386 55383 23442 55392
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 22100 53440 22152 53446
rect 22100 53382 22152 53388
rect 21456 48000 21508 48006
rect 21456 47942 21508 47948
rect 21088 46980 21140 46986
rect 21088 46922 21140 46928
rect 21100 35766 21128 46922
rect 21088 35760 21140 35766
rect 21088 35702 21140 35708
rect 21100 35494 21128 35702
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 21192 33862 21220 35566
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 21192 32570 21220 33798
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 20812 32496 20864 32502
rect 20864 32456 21128 32484
rect 20812 32438 20864 32444
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20536 31408 20588 31414
rect 20536 31350 20588 31356
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20640 29578 20668 30194
rect 20824 29714 20852 32166
rect 21100 31754 21128 32456
rect 21468 31754 21496 47942
rect 22112 47598 22140 53382
rect 23400 53106 23428 55383
rect 23754 54632 23810 54641
rect 23754 54567 23810 54576
rect 23768 53582 23796 54567
rect 24504 54194 24532 56200
rect 24492 54188 24544 54194
rect 24492 54130 24544 54136
rect 24676 53984 24728 53990
rect 24676 53926 24728 53932
rect 23756 53576 23808 53582
rect 23756 53518 23808 53524
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 23388 53100 23440 53106
rect 23388 53042 23440 53048
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22100 47592 22152 47598
rect 22100 47534 22152 47540
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23952 44198 23980 53382
rect 24124 51808 24176 51814
rect 24124 51750 24176 51756
rect 23940 44192 23992 44198
rect 23940 44134 23992 44140
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 24136 43858 24164 51750
rect 24124 43852 24176 43858
rect 24124 43794 24176 43800
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21376 31726 21496 31754
rect 20996 31680 21048 31686
rect 20916 31640 20996 31668
rect 20916 30666 20944 31640
rect 20996 31622 21048 31628
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 20904 30660 20956 30666
rect 20904 30602 20956 30608
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20364 28150 20392 29106
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 20548 28150 20576 28562
rect 20352 28144 20404 28150
rect 20352 28086 20404 28092
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19800 25152 19852 25158
rect 19800 25094 19852 25100
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 24274 19472 24754
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19432 24268 19484 24274
rect 19352 24228 19432 24256
rect 19352 20602 19380 24228
rect 19432 24210 19484 24216
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19444 21554 19472 23598
rect 19536 21978 19564 23734
rect 19628 22098 19656 24686
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19720 23662 19748 24550
rect 19812 23798 19840 25094
rect 19904 23866 19932 25638
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 19996 24313 20024 25162
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 19982 24304 20038 24313
rect 19982 24239 20038 24248
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 19996 23662 20024 24074
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19904 23118 19932 23462
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19536 21950 19748 21978
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19616 21412 19668 21418
rect 19616 21354 19668 21360
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18616 3913 18644 5646
rect 18602 3904 18658 3913
rect 18602 3839 18658 3848
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18432 800 18460 2790
rect 18708 2650 18736 6802
rect 18800 4622 18828 9862
rect 18892 8974 18920 12582
rect 19168 12306 19196 19654
rect 19260 18290 19288 19722
rect 19352 18834 19380 19994
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19246 18184 19302 18193
rect 19246 18119 19302 18128
rect 19260 14006 19288 18119
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 16658 19472 17614
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16114 19380 16390
rect 19444 16114 19472 16594
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19536 15366 19564 20946
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19260 12238 19288 13942
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19064 9376 19116 9382
rect 19062 9344 19064 9353
rect 19116 9344 19118 9353
rect 19062 9279 19118 9288
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18892 7818 18920 8026
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18984 7342 19012 8366
rect 19076 8265 19104 8842
rect 19062 8256 19118 8265
rect 19062 8191 19118 8200
rect 18972 7336 19024 7342
rect 19168 7290 19196 12106
rect 19352 11898 19380 14962
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19536 12238 19564 14554
rect 19628 14414 19656 21354
rect 19720 20942 19748 21950
rect 19904 20942 19932 22646
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 20088 21486 20116 22442
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20180 21690 20208 22374
rect 20272 22030 20300 24822
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20456 24274 20484 24686
rect 20640 24614 20668 29514
rect 20824 28626 20852 29650
rect 20916 29102 20944 30602
rect 21008 30394 21036 30738
rect 21284 30598 21312 31690
rect 21272 30592 21324 30598
rect 21272 30534 21324 30540
rect 20996 30388 21048 30394
rect 20996 30330 21048 30336
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 21284 28626 21312 30534
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21284 28490 21312 28562
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 20824 27402 20852 28426
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20824 27062 20852 27338
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 20824 26382 20852 26998
rect 20916 26450 20944 27270
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26586 21128 26930
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21192 26586 21220 26726
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21180 26580 21232 26586
rect 21180 26522 21232 26528
rect 20904 26444 20956 26450
rect 20956 26404 21036 26432
rect 20904 26386 20956 26392
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 20456 23186 20484 24210
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19720 13954 19748 15370
rect 19628 13926 19748 13954
rect 19628 13682 19656 13926
rect 19708 13864 19760 13870
rect 19706 13832 19708 13841
rect 19760 13832 19762 13841
rect 19706 13767 19762 13776
rect 19628 13654 19748 13682
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19720 12102 19748 13654
rect 19812 12850 19840 16526
rect 19996 15162 20024 20810
rect 20088 19938 20116 21422
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20180 20058 20208 20402
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20088 19910 20208 19938
rect 20180 19786 20208 19910
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20088 16130 20116 19110
rect 20180 17882 20208 19722
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20272 16658 20300 19858
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 16250 20208 16458
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20088 16102 20208 16130
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20088 15366 20116 15982
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20088 14958 20116 15302
rect 20180 15094 20208 16102
rect 20272 15994 20300 16594
rect 20364 16266 20392 22034
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 19514 20484 21286
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 17338 20484 18702
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16590 20484 16934
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20548 16454 20576 23462
rect 20732 23118 20760 25638
rect 20916 25294 20944 25706
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 20916 23322 20944 23802
rect 21008 23662 21036 26404
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 24410 21128 24754
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 21100 24206 21128 24346
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20824 22438 20852 23258
rect 21376 23254 21404 31726
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20364 16238 20576 16266
rect 20352 16040 20404 16046
rect 20272 15988 20352 15994
rect 20272 15982 20404 15988
rect 20272 15966 20392 15982
rect 20272 15570 20300 15966
rect 20548 15910 20576 16238
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19904 12714 19932 13398
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19708 12096 19760 12102
rect 19444 12044 19708 12050
rect 19444 12038 19760 12044
rect 19444 12022 19748 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11694 19472 12022
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19536 11082 19564 11562
rect 19628 11354 19656 11698
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19628 10742 19656 11154
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19260 9178 19288 9522
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19260 8974 19288 9007
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19248 8832 19300 8838
rect 19246 8800 19248 8809
rect 19300 8800 19302 8809
rect 19246 8735 19302 8744
rect 19352 8362 19380 10406
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19444 9042 19472 9930
rect 19522 9072 19578 9081
rect 19432 9036 19484 9042
rect 19522 9007 19578 9016
rect 19432 8978 19484 8984
rect 19536 8906 19564 9007
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 18972 7278 19024 7284
rect 19076 7262 19196 7290
rect 18878 5400 18934 5409
rect 18878 5335 18934 5344
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18800 800 18828 3606
rect 18892 3534 18920 5335
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19076 2446 19104 7262
rect 19260 7002 19288 7346
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19352 6798 19380 7686
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 5234 19288 6598
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19444 4486 19472 8774
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 6458 19564 7890
rect 19628 7342 19656 10678
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19536 5166 19564 6394
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19168 800 19196 3402
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19536 800 19564 3334
rect 19628 2378 19656 5646
rect 19720 3534 19748 9862
rect 19812 4622 19840 11494
rect 19996 9654 20024 14214
rect 20364 13938 20392 14282
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13462 20208 13670
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20180 11150 20208 13398
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20272 12306 20300 13194
rect 20364 12986 20392 13194
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20548 12782 20576 15846
rect 20640 15162 20668 21898
rect 20732 19514 20760 22374
rect 21008 20942 21036 22986
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21100 22545 21128 22578
rect 21086 22536 21142 22545
rect 21086 22471 21142 22480
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 21010 21128 22374
rect 21272 21072 21324 21078
rect 21272 21014 21324 21020
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20824 19718 20852 19994
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20732 15042 20760 18566
rect 20640 15014 20760 15042
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20640 12434 20668 15014
rect 20824 13938 20852 19450
rect 20916 19310 20944 19654
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18970 21128 19110
rect 21192 18970 21220 20334
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20916 13274 20944 18022
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 21008 16674 21036 17546
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21100 16794 21128 17138
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21008 16646 21128 16674
rect 21100 16590 21128 16646
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20824 13246 20944 13274
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20548 12406 20668 12434
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19904 9178 19932 9318
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19996 8974 20024 9318
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19904 6866 19932 8502
rect 19984 8288 20036 8294
rect 20088 8276 20116 10066
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20180 9042 20208 9454
rect 20272 9450 20300 12242
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20180 8634 20208 8978
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20272 8566 20300 9386
rect 20364 8809 20392 9590
rect 20350 8800 20406 8809
rect 20350 8735 20406 8744
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20036 8248 20116 8276
rect 19984 8230 20036 8236
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19904 5302 19932 6802
rect 19996 6662 20024 8230
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19904 3670 19932 4626
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19904 2514 19932 2858
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19616 2372 19668 2378
rect 19616 2314 19668 2320
rect 19996 2122 20024 3946
rect 20088 3233 20116 5782
rect 20180 4282 20208 7754
rect 20456 6848 20484 11018
rect 20548 9994 20576 12406
rect 20732 12288 20760 12786
rect 20640 12260 20760 12288
rect 20640 11898 20668 12260
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 10606 20760 12106
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20824 10062 20852 13246
rect 21008 12918 21036 14962
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 21100 12753 21128 13670
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21086 12744 21142 12753
rect 21086 12679 21142 12688
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20640 8401 20668 9386
rect 20812 8968 20864 8974
rect 20904 8968 20956 8974
rect 20812 8910 20864 8916
rect 20902 8936 20904 8945
rect 20956 8936 20958 8945
rect 20720 8424 20772 8430
rect 20626 8392 20682 8401
rect 20720 8366 20772 8372
rect 20626 8327 20682 8336
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7274 20668 7822
rect 20732 7410 20760 8366
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20456 6820 20576 6848
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20074 3224 20130 3233
rect 20272 3194 20300 6258
rect 20456 6118 20484 6666
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20364 5710 20392 6054
rect 20442 5808 20498 5817
rect 20442 5743 20444 5752
rect 20496 5743 20498 5752
rect 20444 5714 20496 5720
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20074 3159 20130 3168
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20364 2774 20392 5510
rect 20548 3618 20576 6820
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20640 5166 20668 5578
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20628 5024 20680 5030
rect 20824 4978 20852 8910
rect 20902 8871 20958 8880
rect 21008 8786 21036 12378
rect 21100 11830 21128 12679
rect 21192 12434 21220 13126
rect 21284 12986 21312 21014
rect 21468 18766 21496 28698
rect 21744 27130 21772 34138
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 21916 30048 21968 30054
rect 21916 29990 21968 29996
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21732 27124 21784 27130
rect 21732 27066 21784 27072
rect 21640 26512 21692 26518
rect 21640 26454 21692 26460
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21376 13394 21404 16186
rect 21468 16182 21496 16526
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 21468 15434 21496 16118
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21560 15314 21588 16390
rect 21468 15286 21588 15314
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21192 12406 21404 12434
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20680 4972 20852 4978
rect 20628 4966 20852 4972
rect 20640 4950 20852 4966
rect 20916 8758 21036 8786
rect 20916 4690 20944 8758
rect 21100 8498 21128 10610
rect 21192 10130 21220 11154
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21284 10062 21312 11154
rect 21376 10742 21404 12406
rect 21364 10736 21416 10742
rect 21468 10713 21496 15286
rect 21652 14006 21680 26454
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21744 22710 21772 25094
rect 21836 23866 21864 27270
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21836 22778 21864 23054
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21690 21864 21898
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 20942 21864 21490
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21928 18698 21956 29990
rect 22112 27606 22140 31350
rect 22204 31346 22232 43590
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22836 40180 22888 40186
rect 22836 40122 22888 40128
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22296 32978 22324 33526
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22388 33114 22416 33390
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22296 31346 22324 32438
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 22204 28150 22232 28970
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22100 27600 22152 27606
rect 22100 27542 22152 27548
rect 22112 26042 22140 27542
rect 22204 27470 22232 28086
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22204 26081 22232 26318
rect 22190 26072 22246 26081
rect 22100 26036 22152 26042
rect 22190 26007 22246 26016
rect 22100 25978 22152 25984
rect 22296 24750 22324 26386
rect 22388 26382 22416 31622
rect 22480 30326 22508 34886
rect 22560 33856 22612 33862
rect 22560 33798 22612 33804
rect 22572 33538 22600 33798
rect 22664 33658 22692 35566
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22572 33510 22692 33538
rect 22572 31890 22600 33510
rect 22664 33454 22692 33510
rect 22652 33448 22704 33454
rect 22652 33390 22704 33396
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22664 31414 22692 31826
rect 22756 31754 22784 35634
rect 22848 31906 22876 40122
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22928 33924 22980 33930
rect 22928 33866 22980 33872
rect 22940 33590 22968 33866
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23216 33658 23244 33798
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 22928 33584 22980 33590
rect 22928 33526 22980 33532
rect 22940 33318 22968 33526
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 33114 23336 35090
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 23400 32994 23428 35430
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23308 32966 23428 32994
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22848 31878 22968 31906
rect 22940 31822 22968 31878
rect 22836 31816 22888 31822
rect 22836 31758 22888 31764
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 22744 31748 22796 31754
rect 22744 31690 22796 31696
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22664 30938 22692 31350
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22756 30682 22784 31690
rect 22572 30654 22784 30682
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22572 27334 22600 30654
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22664 26790 22692 27950
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22020 21894 22048 23666
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22008 21480 22060 21486
rect 22006 21448 22008 21457
rect 22060 21448 22062 21457
rect 22006 21383 22062 21392
rect 22112 21146 22140 24074
rect 22204 21706 22232 24550
rect 22296 24138 22324 24686
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22388 22710 22416 25978
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22204 21678 22324 21706
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22204 21078 22232 21490
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22112 20602 22140 20878
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22100 20392 22152 20398
rect 22098 20360 22100 20369
rect 22152 20360 22154 20369
rect 22098 20295 22154 20304
rect 22296 20210 22324 21678
rect 22480 21570 22508 26454
rect 22664 24750 22692 26726
rect 22756 26042 22784 30534
rect 22848 30190 22876 31758
rect 23308 31686 23336 32966
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23308 29102 23336 30126
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23400 28234 23428 31894
rect 23492 29578 23520 34682
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23492 28694 23520 29106
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 23308 28218 23428 28234
rect 23296 28212 23428 28218
rect 23348 28206 23428 28212
rect 23296 28154 23348 28160
rect 23492 28098 23520 28630
rect 23584 28626 23612 32982
rect 23676 32910 23704 33254
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23676 32502 23704 32846
rect 23664 32496 23716 32502
rect 23664 32438 23716 32444
rect 23768 32026 23796 39238
rect 23848 32972 23900 32978
rect 23848 32914 23900 32920
rect 23756 32020 23808 32026
rect 23756 31962 23808 31968
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23676 30190 23704 31078
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 23676 28150 23704 30126
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 28422 23796 29038
rect 23860 28626 23888 32914
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24504 31414 24532 32506
rect 24492 31408 24544 31414
rect 24492 31350 24544 31356
rect 24504 30410 24532 31350
rect 24688 31278 24716 53926
rect 25042 53816 25098 53825
rect 25042 53751 25098 53760
rect 25056 53582 25084 53751
rect 25044 53576 25096 53582
rect 25044 53518 25096 53524
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 25780 52896 25832 52902
rect 25780 52838 25832 52844
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24964 52193 24992 52362
rect 24950 52184 25006 52193
rect 24950 52119 25006 52128
rect 24950 51368 25006 51377
rect 24950 51303 24952 51312
rect 25004 51303 25006 51312
rect 24952 51274 25004 51280
rect 25044 51264 25096 51270
rect 25044 51206 25096 51212
rect 24952 50924 25004 50930
rect 24952 50866 25004 50872
rect 24964 50561 24992 50866
rect 24950 50552 25006 50561
rect 24950 50487 25006 50496
rect 24860 49836 24912 49842
rect 24860 49778 24912 49784
rect 24872 49745 24900 49778
rect 24858 49736 24914 49745
rect 24858 49671 24914 49680
rect 25056 45554 25084 51206
rect 25792 49178 25820 52838
rect 25884 52018 25912 56200
rect 26516 53440 26568 53446
rect 26516 53382 26568 53388
rect 25964 52488 26016 52494
rect 25964 52430 26016 52436
rect 25872 52012 25924 52018
rect 25872 51954 25924 51960
rect 25136 49156 25188 49162
rect 25792 49150 25912 49178
rect 25136 49098 25188 49104
rect 25148 48929 25176 49098
rect 25228 49088 25280 49094
rect 25228 49030 25280 49036
rect 25134 48920 25190 48929
rect 25134 48855 25190 48864
rect 25134 48104 25190 48113
rect 25134 48039 25136 48048
rect 25188 48039 25190 48048
rect 25136 48010 25188 48016
rect 24872 45526 25084 45554
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 44033 24808 44338
rect 24766 44024 24822 44033
rect 24766 43959 24822 43968
rect 24872 38350 24900 45526
rect 24952 44736 25004 44742
rect 24952 44678 25004 44684
rect 24860 38344 24912 38350
rect 24860 38286 24912 38292
rect 24860 38208 24912 38214
rect 24860 38150 24912 38156
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 24780 32570 24808 32914
rect 24872 32586 24900 38150
rect 24964 35086 24992 44678
rect 25240 44266 25268 49030
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 25332 47297 25360 47602
rect 25412 47456 25464 47462
rect 25412 47398 25464 47404
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25228 44260 25280 44266
rect 25228 44202 25280 44208
rect 25136 43308 25188 43314
rect 25136 43250 25188 43256
rect 25148 43217 25176 43250
rect 25134 43208 25190 43217
rect 25134 43143 25190 43152
rect 25228 43104 25280 43110
rect 25228 43046 25280 43052
rect 25136 42628 25188 42634
rect 25136 42570 25188 42576
rect 25148 42401 25176 42570
rect 25134 42392 25190 42401
rect 25134 42327 25190 42336
rect 25240 41721 25268 43046
rect 25226 41712 25282 41721
rect 25226 41647 25282 41656
rect 25134 41576 25190 41585
rect 25134 41511 25136 41520
rect 25188 41511 25190 41520
rect 25136 41482 25188 41488
rect 25228 41472 25280 41478
rect 25226 41440 25228 41449
rect 25280 41440 25282 41449
rect 25226 41375 25282 41384
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25320 40044 25372 40050
rect 25320 39986 25372 39992
rect 25332 39953 25360 39986
rect 25318 39944 25374 39953
rect 25318 39879 25374 39888
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25228 38344 25280 38350
rect 25320 38344 25372 38350
rect 25228 38286 25280 38292
rect 25318 38312 25320 38321
rect 25372 38312 25374 38321
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 37505 25176 37810
rect 25134 37496 25190 37505
rect 25134 37431 25190 37440
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 25148 36689 25176 36722
rect 25134 36680 25190 36689
rect 25134 36615 25190 36624
rect 25240 36378 25268 38286
rect 25318 38247 25374 38256
rect 25228 36372 25280 36378
rect 25228 36314 25280 36320
rect 25424 36258 25452 47398
rect 25780 45824 25832 45830
rect 25780 45766 25832 45772
rect 25504 44260 25556 44266
rect 25504 44202 25556 44208
rect 25148 36230 25452 36258
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 25148 33130 25176 36230
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 25056 33102 25176 33130
rect 25240 33114 25268 35974
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25374 34176
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 33425 25360 33934
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25228 33108 25280 33114
rect 24768 32564 24820 32570
rect 24872 32558 24992 32586
rect 24768 32506 24820 32512
rect 24964 32314 24992 32558
rect 24872 32286 24992 32314
rect 24872 31482 24900 32286
rect 25056 32178 25084 33102
rect 25228 33050 25280 33056
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25148 32366 25176 32914
rect 25228 32836 25280 32842
rect 25228 32778 25280 32784
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 24964 32150 25084 32178
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24676 31272 24728 31278
rect 24964 31226 24992 32150
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 24676 31214 24728 31220
rect 24872 31198 24992 31226
rect 24504 30382 24624 30410
rect 24596 30326 24624 30382
rect 24584 30320 24636 30326
rect 24584 30262 24636 30268
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23952 29238 23980 29446
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 24596 29170 24624 30262
rect 24872 29306 24900 31198
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 23848 28620 23900 28626
rect 23848 28562 23900 28568
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23664 28144 23716 28150
rect 23400 28082 23612 28098
rect 23664 28086 23716 28092
rect 23388 28076 23612 28082
rect 23440 28070 23612 28076
rect 23388 28018 23440 28024
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 22848 27674 22876 27814
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 22848 27538 22876 27610
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22848 26314 22876 27270
rect 23308 26926 23336 27406
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22848 25922 22876 26250
rect 22756 25894 22876 25922
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22664 23118 22692 23462
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22388 21542 22508 21570
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22388 21350 22416 21542
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22112 20182 22324 20210
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22020 18426 22048 18634
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21836 15502 21864 17546
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 22020 15706 22048 17002
rect 22112 16522 22140 20182
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22112 15042 22140 15370
rect 22204 15162 22232 17138
rect 22296 16590 22324 19178
rect 22388 17218 22416 20946
rect 22572 20466 22600 21558
rect 22664 20942 22692 22918
rect 22756 21078 22784 25894
rect 23308 25838 23336 26862
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 22848 23594 22876 25774
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23492 24818 23520 27270
rect 23584 27062 23612 28070
rect 23768 27962 23796 28358
rect 23676 27934 23796 27962
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23584 24750 23612 25774
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24342 23336 24686
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23204 23656 23256 23662
rect 23308 23610 23336 24278
rect 23572 24132 23624 24138
rect 23572 24074 23624 24080
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23662 23520 24006
rect 23480 23656 23532 23662
rect 23256 23604 23336 23610
rect 23204 23598 23336 23604
rect 22836 23588 22888 23594
rect 23216 23582 23336 23598
rect 22836 23530 22888 23536
rect 22848 22166 22876 23530
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22836 22160 22888 22166
rect 22836 22102 22888 22108
rect 23204 22094 23256 22098
rect 23308 22094 23336 23582
rect 23386 23624 23442 23633
rect 23480 23598 23532 23604
rect 23386 23559 23442 23568
rect 23400 23186 23428 23559
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23204 22092 23336 22094
rect 23256 22066 23336 22092
rect 23204 22034 23256 22040
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22744 21072 22796 21078
rect 22744 21014 22796 21020
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22572 17678 22600 18838
rect 22664 18766 22692 20198
rect 22756 19922 22784 20334
rect 22848 19938 22876 21626
rect 22940 21350 22968 21966
rect 23216 21554 23244 22034
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 23400 21434 23428 21830
rect 23492 21622 23520 23598
rect 23584 21622 23612 24074
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23308 21406 23428 21434
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22744 19916 22796 19922
rect 22848 19910 22968 19938
rect 22744 19858 22796 19864
rect 22756 19360 22784 19858
rect 22836 19372 22888 19378
rect 22756 19332 22836 19360
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22756 18290 22784 19332
rect 22836 19314 22888 19320
rect 22940 19310 22968 19910
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 23308 19242 23336 21406
rect 23584 21350 23612 21558
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23388 21072 23440 21078
rect 23388 21014 23440 21020
rect 23296 19236 23348 19242
rect 23296 19178 23348 19184
rect 23400 19174 23428 21014
rect 23584 20534 23612 21286
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23584 20058 23612 20470
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23584 18766 23612 19382
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23676 18358 23704 27934
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 24044 26382 24072 27639
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 23952 22642 23980 25298
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 24136 24410 24164 24822
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23768 22234 23796 22578
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 20058 23888 20946
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23860 19666 23888 19994
rect 23768 19638 23888 19666
rect 23768 19446 23796 19638
rect 23846 19544 23902 19553
rect 23846 19479 23902 19488
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 23860 18834 23888 19479
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22388 17190 22600 17218
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22008 15020 22060 15026
rect 22112 15014 22232 15042
rect 22008 14962 22060 14968
rect 22020 14906 22048 14962
rect 21916 14884 21968 14890
rect 22020 14878 22140 14906
rect 21916 14826 21968 14832
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21364 10678 21416 10684
rect 21454 10704 21510 10713
rect 21454 10639 21510 10648
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21468 10130 21496 10542
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20904 4208 20956 4214
rect 20904 4150 20956 4156
rect 20548 3590 20760 3618
rect 20732 3534 20760 3590
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20718 3360 20774 3369
rect 20718 3295 20774 3304
rect 20732 3058 20760 3295
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 19904 2094 20024 2122
rect 20272 2746 20392 2774
rect 19904 800 19932 2094
rect 20272 800 20300 2746
rect 20640 800 20668 2858
rect 20916 2650 20944 4150
rect 21008 4146 21036 7958
rect 21284 6798 21312 8366
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21272 6792 21324 6798
rect 21270 6760 21272 6769
rect 21324 6760 21326 6769
rect 21270 6695 21326 6704
rect 21284 5302 21312 6695
rect 21272 5296 21324 5302
rect 21272 5238 21324 5244
rect 21468 5098 21496 6938
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21008 800 21036 3878
rect 21100 3398 21128 4490
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21284 2922 21312 4966
rect 21468 4078 21496 5034
rect 21560 4622 21588 11562
rect 21652 11354 21680 11698
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21836 9674 21864 13738
rect 21928 11082 21956 14826
rect 22112 12646 22140 14878
rect 22204 14362 22232 15014
rect 22296 14482 22324 15506
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22204 14346 22324 14362
rect 22204 14340 22336 14346
rect 22204 14334 22284 14340
rect 22284 14282 22336 14288
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11558 22140 12174
rect 22204 11898 22232 12786
rect 22296 12238 22324 14282
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22388 11830 22416 16526
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10470 22048 10950
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10198 22140 10406
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22204 9722 22232 11698
rect 22296 10130 22324 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22192 9716 22244 9722
rect 21836 9646 22048 9674
rect 22192 9658 22244 9664
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21376 800 21404 2858
rect 21652 2650 21680 7754
rect 21744 6662 21772 9114
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21744 5914 21772 6258
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21836 2417 21864 8842
rect 22020 8838 22048 9646
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21928 5137 21956 7278
rect 21914 5128 21970 5137
rect 21914 5063 21970 5072
rect 22020 3126 22048 8774
rect 22204 8090 22232 9386
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22296 7954 22324 10066
rect 22388 9450 22416 11290
rect 22480 9602 22508 17002
rect 22572 15434 22600 17190
rect 22664 17066 22692 17478
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 16046 22692 16186
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22664 15570 22692 15846
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22572 15162 22600 15370
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 12986 22600 14962
rect 22664 14958 22692 15506
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22756 13920 22784 18022
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22664 13892 22784 13920
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22664 11626 22692 13892
rect 22848 13818 22876 17478
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16250 23336 18090
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23308 15162 23336 15506
rect 23676 15502 23704 15982
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 22756 13790 22876 13818
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22756 11150 22784 13790
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 12918 23336 14214
rect 23492 13394 23520 15302
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22848 11762 22876 12718
rect 23400 12646 23428 13330
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23400 11830 23428 12582
rect 23584 12238 23612 14758
rect 23676 14414 23704 15438
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23676 12730 23704 14350
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23768 12730 23796 12854
rect 23676 12702 23796 12730
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23676 12170 23704 12702
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22572 10266 22600 10610
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22664 10130 22692 10542
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22664 9722 22692 9930
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22480 9574 22692 9602
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22376 9444 22428 9450
rect 22376 9386 22428 9392
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22296 7834 22324 7890
rect 22112 7806 22324 7834
rect 22112 7002 22140 7806
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 22112 2938 22140 6190
rect 22190 5808 22246 5817
rect 22190 5743 22246 5752
rect 22284 5772 22336 5778
rect 22204 5710 22232 5743
rect 22284 5714 22336 5720
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22296 4026 22324 5714
rect 22020 2910 22140 2938
rect 22204 3998 22324 4026
rect 22204 2922 22232 3998
rect 22282 3904 22338 3913
rect 22282 3839 22338 3848
rect 22296 3126 22324 3839
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 22192 2916 22244 2922
rect 21822 2408 21878 2417
rect 21822 2343 21878 2352
rect 21744 870 21864 898
rect 21744 800 21772 870
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 21836 762 21864 870
rect 22020 762 22048 2910
rect 22192 2858 22244 2864
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 2514 22140 2790
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22100 1964 22152 1970
rect 22100 1906 22152 1912
rect 22112 1601 22140 1906
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 22296 1442 22324 2858
rect 22388 2774 22416 8366
rect 22480 5409 22508 8434
rect 22572 7954 22600 9454
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22466 5400 22522 5409
rect 22466 5335 22522 5344
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 3058 22508 4422
rect 22572 4026 22600 6326
rect 22664 4214 22692 9574
rect 22756 8974 22784 10950
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22848 9518 22876 9862
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23308 9081 23336 11290
rect 23492 10538 23520 12038
rect 23676 11830 23704 12106
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23584 9602 23612 10406
rect 23676 10062 23704 11766
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23860 10062 23888 11222
rect 23664 10056 23716 10062
rect 23848 10056 23900 10062
rect 23716 10004 23796 10010
rect 23664 9998 23796 10004
rect 23848 9998 23900 10004
rect 23676 9982 23796 9998
rect 23768 9738 23796 9982
rect 23768 9710 23888 9738
rect 23388 9580 23440 9586
rect 23584 9574 23796 9602
rect 23388 9522 23440 9528
rect 23294 9072 23350 9081
rect 23294 9007 23350 9016
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 22572 3998 22692 4026
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22664 2922 22692 3998
rect 22756 2922 22784 5306
rect 22848 4049 22876 6054
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5681 23336 7278
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4826 23428 9522
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 22834 4040 22890 4049
rect 22834 3975 22890 3984
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23492 3602 23520 8434
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23216 3194 23244 3470
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22388 2746 22508 2774
rect 22112 1414 22324 1442
rect 22112 800 22140 1414
rect 22480 800 22508 2746
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 22848 800 22876 2314
rect 23216 800 23244 2586
rect 23584 800 23612 9454
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23676 6798 23704 7822
rect 23664 6792 23716 6798
rect 23662 6760 23664 6769
rect 23716 6760 23718 6769
rect 23662 6695 23718 6704
rect 23676 3194 23704 6695
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23768 2446 23796 9574
rect 23860 7954 23888 9710
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23860 6458 23888 6598
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23952 800 23980 21082
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24044 19394 24072 19790
rect 24124 19440 24176 19446
rect 24044 19388 24124 19394
rect 24044 19382 24176 19388
rect 24044 19366 24164 19382
rect 24044 18358 24072 19366
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24044 16998 24072 18294
rect 24136 17202 24164 18566
rect 24228 18222 24256 27814
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24320 17338 24348 28970
rect 24780 28529 24808 29106
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24766 28520 24822 28529
rect 24766 28455 24822 28464
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24596 27674 24624 28018
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24412 25974 24440 27066
rect 24584 26852 24636 26858
rect 24584 26794 24636 26800
rect 24596 26314 24624 26794
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24400 25968 24452 25974
rect 24400 25910 24452 25916
rect 24412 24886 24440 25910
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 24412 24138 24440 24822
rect 24766 24440 24822 24449
rect 24766 24375 24822 24384
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24412 24018 24440 24074
rect 24412 23990 24532 24018
rect 24504 23798 24532 23990
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 19514 24624 22918
rect 24780 22574 24808 24375
rect 24872 23186 24900 28970
rect 24964 26450 24992 31078
rect 25056 27538 25084 31894
rect 25148 30190 25176 32302
rect 25136 30184 25188 30190
rect 25136 30126 25188 30132
rect 25136 29504 25188 29510
rect 25136 29446 25188 29452
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25148 26858 25176 29446
rect 25240 29238 25268 32778
rect 25424 32609 25452 33458
rect 25410 32600 25466 32609
rect 25410 32535 25466 32544
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25332 30977 25360 31282
rect 25318 30968 25374 30977
rect 25318 30903 25374 30912
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25424 29345 25452 30670
rect 25410 29336 25466 29345
rect 25410 29271 25466 29280
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 25228 27532 25280 27538
rect 25228 27474 25280 27480
rect 25240 26926 25268 27474
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 25318 26888 25374 26897
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24952 26444 25004 26450
rect 24952 26386 25004 26392
rect 24950 25256 25006 25265
rect 24950 25191 24952 25200
rect 25004 25191 25006 25200
rect 24952 25162 25004 25168
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24858 22808 24914 22817
rect 24858 22743 24914 22752
rect 24872 22710 24900 22743
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24964 20942 24992 24142
rect 25056 22098 25084 26522
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25148 24750 25176 26386
rect 25240 26042 25268 26862
rect 25318 26823 25374 26832
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 25240 24750 25268 25774
rect 25332 25294 25360 26823
rect 25412 26512 25464 26518
rect 25412 26454 25464 26460
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25148 23866 25176 24686
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25240 22166 25268 24686
rect 25424 24206 25452 26454
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25228 22160 25280 22166
rect 25228 22102 25280 22108
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25134 21992 25190 22001
rect 25134 21927 25190 21936
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 25148 20874 25176 21927
rect 25332 21486 25360 23122
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24766 18728 24822 18737
rect 24766 18663 24822 18672
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24688 16114 24716 17478
rect 24780 17134 24808 18663
rect 24872 18034 24900 20742
rect 25332 20602 25360 21422
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19514 25176 20334
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 24872 18006 24992 18034
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17746 24900 17847
rect 24964 17746 24992 18006
rect 25148 17746 25176 19450
rect 25516 18698 25544 44202
rect 25792 41414 25820 45766
rect 25700 41386 25820 41414
rect 25596 37732 25648 37738
rect 25596 37674 25648 37680
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24768 17128 24820 17134
rect 24872 17105 24900 17206
rect 25332 17202 25360 18158
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 24768 17070 24820 17076
rect 24858 17096 24914 17105
rect 24858 17031 24914 17040
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24780 16046 24808 16934
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24872 16289 24900 16458
rect 24858 16280 24914 16289
rect 24858 16215 24914 16224
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 13326 24072 15846
rect 24766 15464 24822 15473
rect 24766 15399 24822 15408
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13938 24164 14214
rect 24596 14006 24624 15302
rect 24780 14958 24808 15399
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24780 14074 24808 14350
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 25148 14006 25176 14583
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24860 13864 24912 13870
rect 24858 13832 24860 13841
rect 24912 13832 24914 13841
rect 24858 13767 24914 13776
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24596 12306 24624 13126
rect 24964 13025 24992 13194
rect 24950 13016 25006 13025
rect 24950 12951 25006 12960
rect 24676 12776 24728 12782
rect 25608 12753 25636 37674
rect 25700 35834 25728 41386
rect 25884 36394 25912 49150
rect 25976 36530 26004 52430
rect 26056 46368 26108 46374
rect 26056 46310 26108 46316
rect 26068 41414 26096 46310
rect 26068 41386 26372 41414
rect 25976 36502 26280 36530
rect 25884 36366 26188 36394
rect 25964 36304 26016 36310
rect 25964 36246 26016 36252
rect 26056 36304 26108 36310
rect 26056 36246 26108 36252
rect 25688 35828 25740 35834
rect 25688 35770 25740 35776
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25700 33402 25728 34886
rect 25700 33374 25820 33402
rect 25688 33108 25740 33114
rect 25688 33050 25740 33056
rect 25700 18426 25728 33050
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25792 17814 25820 33374
rect 25872 33312 25924 33318
rect 25872 33254 25924 33260
rect 25884 27402 25912 33254
rect 25976 30054 26004 36246
rect 25964 30048 26016 30054
rect 25964 29990 26016 29996
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25884 23118 25912 26250
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25780 17808 25832 17814
rect 25780 17750 25832 17756
rect 26068 13462 26096 36246
rect 26160 28490 26188 36366
rect 26252 30870 26280 36502
rect 26344 35766 26372 41386
rect 26424 40928 26476 40934
rect 26424 40870 26476 40876
rect 26332 35760 26384 35766
rect 26332 35702 26384 35708
rect 26436 33046 26464 40870
rect 26424 33040 26476 33046
rect 26424 32982 26476 32988
rect 26240 30864 26292 30870
rect 26240 30806 26292 30812
rect 26528 30802 26556 53382
rect 26700 42628 26752 42634
rect 26700 42570 26752 42576
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 26712 14618 26740 42570
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 24676 12718 24728 12724
rect 25594 12744 25650 12753
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24688 11150 24716 12718
rect 25594 12679 25650 12688
rect 24950 12200 25006 12209
rect 24950 12135 24952 12144
rect 25004 12135 25006 12144
rect 24952 12106 25004 12112
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24044 7970 24072 10746
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 10266 24624 10610
rect 24780 10606 24808 11319
rect 24872 10674 24900 11494
rect 25042 10704 25098 10713
rect 24860 10668 24912 10674
rect 25042 10639 25098 10648
rect 24860 10610 24912 10616
rect 24768 10600 24820 10606
rect 24674 10568 24730 10577
rect 24768 10542 24820 10548
rect 24674 10503 24730 10512
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24136 8090 24164 9522
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24216 8016 24268 8022
rect 24044 7942 24164 7970
rect 24216 7958 24268 7964
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7002 24072 7686
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24044 6186 24072 6598
rect 24032 6180 24084 6186
rect 24032 6122 24084 6128
rect 24136 5234 24164 7942
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24228 4622 24256 7958
rect 24412 4690 24440 9658
rect 24688 9518 24716 10503
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24596 6322 24624 8774
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24688 3534 24716 9046
rect 24780 8430 24808 9687
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24766 6488 24822 6497
rect 24766 6423 24822 6432
rect 24780 5166 24808 6423
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24872 4758 24900 7210
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24320 800 24348 2994
rect 24872 2038 24900 3402
rect 24964 2650 24992 6598
rect 25056 5710 25084 10639
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25134 7304 25190 7313
rect 25134 7239 25190 7248
rect 25148 6390 25176 7239
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 21836 734 22048 762
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25148 785 25176 3674
rect 25134 776 25190 785
rect 25134 711 25190 720
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3514 8744 3570 8800
rect 3422 6432 3478 6488
rect 3882 4120 3938 4176
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3422 1844 3424 1864
rect 3424 1844 3476 1864
rect 3476 1844 3478 1864
rect 3422 1808 3478 1844
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7746 12824 7802 12880
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 9034 18128 9090 18184
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13358 15544 13414 15600
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13634 15408 13690 15464
rect 14830 25064 14886 25120
rect 13450 12960 13506 13016
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12438 4120 12494 4176
rect 12714 8336 12770 8392
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13726 12960 13782 13016
rect 13634 8880 13690 8936
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13174 3052 13230 3088
rect 13174 3032 13176 3052
rect 13176 3032 13228 3052
rect 13228 3032 13230 3052
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 12898 2488 12954 2544
rect 16762 25880 16818 25936
rect 15014 12980 15070 13016
rect 15014 12960 15016 12980
rect 15016 12960 15068 12980
rect 15068 12960 15070 12980
rect 15106 12860 15108 12880
rect 15108 12860 15160 12880
rect 15160 12860 15162 12880
rect 15106 12824 15162 12860
rect 13910 8472 13966 8528
rect 13818 8336 13874 8392
rect 14462 7828 14464 7848
rect 14464 7828 14516 7848
rect 14516 7828 14518 7848
rect 14462 7792 14518 7828
rect 14830 8200 14886 8256
rect 15658 12980 15714 13016
rect 15658 12960 15660 12980
rect 15660 12960 15712 12980
rect 15712 12960 15714 12980
rect 16026 12824 16082 12880
rect 15934 10684 15936 10704
rect 15936 10684 15988 10704
rect 15988 10684 15990 10704
rect 15934 10648 15990 10684
rect 15566 6840 15622 6896
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17314 27956 17316 27976
rect 17316 27956 17368 27976
rect 17368 27956 17370 27976
rect 17314 27920 17370 27956
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 23294 56072 23350 56128
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17314 19352 17370 19408
rect 16946 17448 17002 17504
rect 17222 18264 17278 18320
rect 17130 16632 17186 16688
rect 16762 12708 16818 12744
rect 16762 12688 16764 12708
rect 16764 12688 16816 12708
rect 16816 12688 16818 12708
rect 16946 10104 17002 10160
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17130 9016 17186 9072
rect 17130 8492 17186 8528
rect 17130 8472 17132 8492
rect 17132 8472 17184 8492
rect 17184 8472 17186 8492
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18142 15972 18198 16008
rect 18142 15952 18144 15972
rect 18144 15952 18196 15972
rect 18196 15952 18198 15972
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17866 13640 17922 13696
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18326 12688 18382 12744
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17498 9460 17500 9480
rect 17500 9460 17552 9480
rect 17552 9460 17554 9480
rect 17498 9424 17554 9460
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18694 15952 18750 16008
rect 18234 10140 18236 10160
rect 18236 10140 18288 10160
rect 18288 10140 18290 10160
rect 18234 10104 18290 10140
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17498 9324 17500 9344
rect 17500 9324 17552 9344
rect 17552 9324 17554 9344
rect 17498 9288 17554 9324
rect 18326 9424 18382 9480
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 23386 55392 23442 55448
rect 23754 54576 23810 54632
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 19982 24248 20038 24304
rect 18602 3848 18658 3904
rect 19246 18128 19302 18184
rect 19062 9324 19064 9344
rect 19064 9324 19116 9344
rect 19116 9324 19118 9344
rect 19062 9288 19118 9324
rect 19062 8200 19118 8256
rect 19706 13812 19708 13832
rect 19708 13812 19760 13832
rect 19760 13812 19762 13832
rect 19706 13776 19762 13812
rect 19246 9016 19302 9072
rect 19246 8780 19248 8800
rect 19248 8780 19300 8800
rect 19300 8780 19302 8800
rect 19246 8744 19302 8780
rect 19522 9016 19578 9072
rect 18878 5344 18934 5400
rect 21086 22480 21142 22536
rect 20350 8744 20406 8800
rect 21086 12688 21142 12744
rect 20902 8916 20904 8936
rect 20904 8916 20956 8936
rect 20956 8916 20958 8936
rect 20626 8336 20682 8392
rect 20074 3168 20130 3224
rect 20442 5772 20498 5808
rect 20442 5752 20444 5772
rect 20444 5752 20496 5772
rect 20496 5752 20498 5772
rect 20902 8880 20958 8916
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22190 26016 22246 26072
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22006 21428 22008 21448
rect 22008 21428 22060 21448
rect 22060 21428 22062 21448
rect 22006 21392 22062 21428
rect 22098 20340 22100 20360
rect 22100 20340 22152 20360
rect 22152 20340 22154 20360
rect 22098 20304 22154 20340
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 25042 53760 25098 53816
rect 25042 52944 25098 53000
rect 24950 52128 25006 52184
rect 24950 51332 25006 51368
rect 24950 51312 24952 51332
rect 24952 51312 25004 51332
rect 25004 51312 25006 51332
rect 24950 50496 25006 50552
rect 24858 49680 24914 49736
rect 25134 48864 25190 48920
rect 25134 48068 25190 48104
rect 25134 48048 25136 48068
rect 25136 48048 25188 48068
rect 25188 48048 25190 48068
rect 24766 43968 24822 44024
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 25134 43152 25190 43208
rect 25134 42336 25190 42392
rect 25226 41656 25282 41712
rect 25134 41540 25190 41576
rect 25134 41520 25136 41540
rect 25136 41520 25188 41540
rect 25188 41520 25190 41540
rect 25226 41420 25228 41440
rect 25228 41420 25280 41440
rect 25280 41420 25282 41440
rect 25226 41384 25282 41420
rect 25318 40704 25374 40760
rect 25318 39888 25374 39944
rect 25318 39072 25374 39128
rect 25318 38292 25320 38312
rect 25320 38292 25372 38312
rect 25372 38292 25374 38312
rect 25134 37440 25190 37496
rect 25134 36624 25190 36680
rect 25318 38256 25374 38292
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34176 25374 34232
rect 25318 33360 25374 33416
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23386 23568 23442 23624
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 24030 27648 24086 27704
rect 23846 19488 23902 19544
rect 21454 10648 21510 10704
rect 20718 3304 20774 3360
rect 21270 6740 21272 6760
rect 21272 6740 21324 6760
rect 21324 6740 21326 6760
rect 21270 6704 21326 6740
rect 21914 5072 21970 5128
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22190 5752 22246 5808
rect 22282 3848 22338 3904
rect 21822 2352 21878 2408
rect 22098 1536 22154 1592
rect 22466 5344 22522 5400
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 23294 9016 23350 9072
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23294 5616 23350 5672
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22834 3984 22890 4040
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23662 6740 23664 6760
rect 23664 6740 23716 6760
rect 23716 6740 23718 6760
rect 23662 6704 23718 6740
rect 24766 28464 24822 28520
rect 24766 24384 24822 24440
rect 25410 32544 25466 32600
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30912 25374 30968
rect 25318 30096 25374 30152
rect 25410 29280 25466 29336
rect 24950 25220 25006 25256
rect 24950 25200 24952 25220
rect 24952 25200 25004 25220
rect 25004 25200 25006 25220
rect 24858 22752 24914 22808
rect 25318 26832 25374 26888
rect 25134 21936 25190 21992
rect 24766 18672 24822 18728
rect 24858 17856 24914 17912
rect 24858 17040 24914 17096
rect 24858 16224 24914 16280
rect 24766 15408 24822 15464
rect 25134 14592 25190 14648
rect 24858 13812 24860 13832
rect 24860 13812 24912 13832
rect 24912 13812 24914 13832
rect 24858 13776 24914 13812
rect 24950 12960 25006 13016
rect 25594 12688 25650 12744
rect 24950 12164 25006 12200
rect 24950 12144 24952 12164
rect 24952 12144 25004 12164
rect 25004 12144 25006 12164
rect 24766 11328 24822 11384
rect 25042 10648 25098 10704
rect 24674 10512 24730 10568
rect 24766 9696 24822 9752
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24766 6432 24822 6488
rect 25134 8064 25190 8120
rect 25134 7248 25190 7304
rect 25134 720 25190 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23289 56130 23355 56133
rect 23430 56130 23490 56206
rect 26200 56176 27000 56206
rect 23289 56128 23490 56130
rect 23289 56072 23294 56128
rect 23350 56072 23490 56128
rect 23289 56070 23490 56072
rect 23289 56067 23355 56070
rect 23381 55450 23447 55453
rect 26200 55450 27000 55480
rect 23381 55448 27000 55450
rect 23381 55392 23386 55448
rect 23442 55392 27000 55448
rect 23381 55390 27000 55392
rect 23381 55387 23447 55390
rect 26200 55360 27000 55390
rect 23749 54634 23815 54637
rect 26200 54634 27000 54664
rect 23749 54632 27000 54634
rect 23749 54576 23754 54632
rect 23810 54576 27000 54632
rect 23749 54574 27000 54576
rect 23749 54571 23815 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 25037 53818 25103 53821
rect 26200 53818 27000 53848
rect 25037 53816 27000 53818
rect 25037 53760 25042 53816
rect 25098 53760 27000 53816
rect 25037 53758 27000 53760
rect 25037 53755 25103 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 24945 51370 25011 51373
rect 26200 51370 27000 51400
rect 24945 51368 27000 51370
rect 24945 51312 24950 51368
rect 25006 51312 27000 51368
rect 24945 51310 27000 51312
rect 24945 51307 25011 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 24945 50554 25011 50557
rect 26200 50554 27000 50584
rect 24945 50552 27000 50554
rect 24945 50496 24950 50552
rect 25006 50496 27000 50552
rect 24945 50494 27000 50496
rect 24945 50491 25011 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 24853 49738 24919 49741
rect 26200 49738 27000 49768
rect 24853 49736 27000 49738
rect 24853 49680 24858 49736
rect 24914 49680 27000 49736
rect 24853 49678 27000 49680
rect 24853 49675 24919 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25129 48922 25195 48925
rect 26200 48922 27000 48952
rect 25129 48920 27000 48922
rect 25129 48864 25134 48920
rect 25190 48864 27000 48920
rect 25129 48862 27000 48864
rect 25129 48859 25195 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25129 48106 25195 48109
rect 26200 48106 27000 48136
rect 25129 48104 27000 48106
rect 25129 48048 25134 48104
rect 25190 48048 27000 48104
rect 25129 48046 27000 48048
rect 25129 48043 25195 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24761 44026 24827 44029
rect 26200 44026 27000 44056
rect 24761 44024 27000 44026
rect 24761 43968 24766 44024
rect 24822 43968 27000 44024
rect 24761 43966 27000 43968
rect 24761 43963 24827 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25129 43210 25195 43213
rect 26200 43210 27000 43240
rect 25129 43208 27000 43210
rect 25129 43152 25134 43208
rect 25190 43152 27000 43208
rect 25129 43150 27000 43152
rect 25129 43147 25195 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25129 42394 25195 42397
rect 26200 42394 27000 42424
rect 25129 42392 27000 42394
rect 25129 42336 25134 42392
rect 25190 42336 27000 42392
rect 25129 42334 27000 42336
rect 25129 42331 25195 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 19190 41652 19196 41716
rect 19260 41714 19266 41716
rect 25221 41714 25287 41717
rect 19260 41712 25287 41714
rect 19260 41656 25226 41712
rect 25282 41656 25287 41712
rect 19260 41654 25287 41656
rect 19260 41652 19266 41654
rect 25221 41651 25287 41654
rect 25129 41578 25195 41581
rect 26200 41578 27000 41608
rect 25129 41576 27000 41578
rect 25129 41520 25134 41576
rect 25190 41520 27000 41576
rect 25129 41518 27000 41520
rect 25129 41515 25195 41518
rect 26200 41488 27000 41518
rect 19926 41380 19932 41444
rect 19996 41442 20002 41444
rect 25221 41442 25287 41445
rect 19996 41440 25287 41442
rect 19996 41384 25226 41440
rect 25282 41384 25287 41440
rect 19996 41382 25287 41384
rect 19996 41380 20002 41382
rect 25221 41379 25287 41382
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25313 39946 25379 39949
rect 26200 39946 27000 39976
rect 25313 39944 27000 39946
rect 25313 39888 25318 39944
rect 25374 39888 27000 39944
rect 25313 39886 27000 39888
rect 25313 39883 25379 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25129 37498 25195 37501
rect 26200 37498 27000 37528
rect 25129 37496 27000 37498
rect 25129 37440 25134 37496
rect 25190 37440 27000 37496
rect 25129 37438 27000 37440
rect 25129 37435 25195 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 25129 36682 25195 36685
rect 26200 36682 27000 36712
rect 25129 36680 27000 36682
rect 25129 36624 25134 36680
rect 25190 36624 27000 36680
rect 25129 36622 27000 36624
rect 25129 36619 25195 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 25405 32602 25471 32605
rect 26200 32602 27000 32632
rect 25405 32600 27000 32602
rect 25405 32544 25410 32600
rect 25466 32544 27000 32600
rect 25405 32542 27000 32544
rect 25405 32539 25471 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 25405 29338 25471 29341
rect 26200 29338 27000 29368
rect 25405 29336 27000 29338
rect 25405 29280 25410 29336
rect 25466 29280 27000 29336
rect 25405 29278 27000 29280
rect 25405 29275 25471 29278
rect 26200 29248 27000 29278
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24761 28522 24827 28525
rect 26200 28522 27000 28552
rect 24761 28520 27000 28522
rect 24761 28464 24766 28520
rect 24822 28464 27000 28520
rect 24761 28462 27000 28464
rect 24761 28459 24827 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 17309 27980 17375 27981
rect 17309 27978 17356 27980
rect 17264 27976 17356 27978
rect 17264 27920 17314 27976
rect 17264 27918 17356 27920
rect 17309 27916 17356 27918
rect 17420 27916 17426 27980
rect 17309 27915 17375 27916
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24025 27706 24091 27709
rect 26200 27706 27000 27736
rect 24025 27704 27000 27706
rect 24025 27648 24030 27704
rect 24086 27648 27000 27704
rect 24025 27646 27000 27648
rect 24025 27643 24091 27646
rect 26200 27616 27000 27646
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25313 26890 25379 26893
rect 26200 26890 27000 26920
rect 25313 26888 27000 26890
rect 25313 26832 25318 26888
rect 25374 26832 27000 26888
rect 25313 26830 27000 26832
rect 25313 26827 25379 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 22185 26074 22251 26077
rect 26200 26074 27000 26104
rect 22185 26072 27000 26074
rect 22185 26016 22190 26072
rect 22246 26016 27000 26072
rect 22185 26014 27000 26016
rect 22185 26011 22251 26014
rect 26200 25984 27000 26014
rect 16757 25940 16823 25941
rect 16757 25936 16804 25940
rect 16868 25938 16874 25940
rect 16757 25880 16762 25936
rect 16757 25876 16804 25880
rect 16868 25878 16914 25938
rect 16868 25876 16874 25878
rect 16757 25875 16823 25876
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 24945 25258 25011 25261
rect 26200 25258 27000 25288
rect 24945 25256 27000 25258
rect 24945 25200 24950 25256
rect 25006 25200 27000 25256
rect 24945 25198 27000 25200
rect 24945 25195 25011 25198
rect 26200 25168 27000 25198
rect 14825 25124 14891 25125
rect 14774 25122 14780 25124
rect 14734 25062 14780 25122
rect 14844 25120 14891 25124
rect 14886 25064 14891 25120
rect 14774 25060 14780 25062
rect 14844 25060 14891 25064
rect 14825 25059 14891 25060
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24761 24442 24827 24445
rect 26200 24442 27000 24472
rect 24761 24440 27000 24442
rect 24761 24384 24766 24440
rect 24822 24384 27000 24440
rect 24761 24382 27000 24384
rect 24761 24379 24827 24382
rect 26200 24352 27000 24382
rect 15694 24244 15700 24308
rect 15764 24306 15770 24308
rect 19977 24306 20043 24309
rect 15764 24304 20043 24306
rect 15764 24248 19982 24304
rect 20038 24248 20043 24304
rect 15764 24246 20043 24248
rect 15764 24244 15770 24246
rect 19977 24243 20043 24246
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 23381 23626 23447 23629
rect 26200 23626 27000 23656
rect 23381 23624 27000 23626
rect 23381 23568 23386 23624
rect 23442 23568 27000 23624
rect 23381 23566 27000 23568
rect 23381 23563 23447 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 24853 22810 24919 22813
rect 26200 22810 27000 22840
rect 24853 22808 27000 22810
rect 24853 22752 24858 22808
rect 24914 22752 27000 22808
rect 24853 22750 27000 22752
rect 24853 22747 24919 22750
rect 26200 22720 27000 22750
rect 20846 22476 20852 22540
rect 20916 22538 20922 22540
rect 21081 22538 21147 22541
rect 20916 22536 21147 22538
rect 20916 22480 21086 22536
rect 21142 22480 21147 22536
rect 20916 22478 21147 22480
rect 20916 22476 20922 22478
rect 21081 22475 21147 22478
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 25129 21994 25195 21997
rect 26200 21994 27000 22024
rect 25129 21992 27000 21994
rect 25129 21936 25134 21992
rect 25190 21936 27000 21992
rect 25129 21934 27000 21936
rect 25129 21931 25195 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 22001 21450 22067 21453
rect 22001 21448 23674 21450
rect 22001 21392 22006 21448
rect 22062 21392 23674 21448
rect 22001 21390 23674 21392
rect 22001 21387 22067 21390
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 23614 21178 23674 21390
rect 26200 21178 27000 21208
rect 23614 21118 27000 21178
rect 26200 21088 27000 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 22093 20362 22159 20365
rect 26200 20362 27000 20392
rect 22093 20360 27000 20362
rect 22093 20304 22098 20360
rect 22154 20304 27000 20360
rect 22093 20302 27000 20304
rect 22093 20299 22159 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23841 19546 23907 19549
rect 26200 19546 27000 19576
rect 23841 19544 27000 19546
rect 23841 19488 23846 19544
rect 23902 19488 27000 19544
rect 23841 19486 27000 19488
rect 23841 19483 23907 19486
rect 26200 19456 27000 19486
rect 17309 19410 17375 19413
rect 17534 19410 17540 19412
rect 17309 19408 17540 19410
rect 17309 19352 17314 19408
rect 17370 19352 17540 19408
rect 17309 19350 17540 19352
rect 17309 19347 17375 19350
rect 17534 19348 17540 19350
rect 17604 19348 17610 19412
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 20846 18730 20852 18732
rect 16530 18670 20852 18730
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 9029 18186 9095 18189
rect 16530 18186 16590 18670
rect 20846 18668 20852 18670
rect 20916 18668 20922 18732
rect 24761 18730 24827 18733
rect 26200 18730 27000 18760
rect 24761 18728 27000 18730
rect 24761 18672 24766 18728
rect 24822 18672 27000 18728
rect 24761 18670 27000 18672
rect 24761 18667 24827 18670
rect 26200 18640 27000 18670
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 17217 18322 17283 18325
rect 17718 18322 17724 18324
rect 17217 18320 17724 18322
rect 17217 18264 17222 18320
rect 17278 18264 17724 18320
rect 17217 18262 17724 18264
rect 17217 18259 17283 18262
rect 17718 18260 17724 18262
rect 17788 18260 17794 18324
rect 9029 18184 16590 18186
rect 9029 18128 9034 18184
rect 9090 18128 16590 18184
rect 9029 18126 16590 18128
rect 19241 18186 19307 18189
rect 19926 18186 19932 18188
rect 19241 18184 19932 18186
rect 19241 18128 19246 18184
rect 19302 18128 19932 18184
rect 19241 18126 19932 18128
rect 9029 18123 9095 18126
rect 19241 18123 19307 18126
rect 19926 18124 19932 18126
rect 19996 18124 20002 18188
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 16798 17444 16804 17508
rect 16868 17506 16874 17508
rect 16941 17506 17007 17509
rect 16868 17504 17007 17506
rect 16868 17448 16946 17504
rect 17002 17448 17007 17504
rect 16868 17446 17007 17448
rect 16868 17444 16874 17446
rect 16941 17443 17007 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24853 17098 24919 17101
rect 26200 17098 27000 17128
rect 24853 17096 27000 17098
rect 24853 17040 24858 17096
rect 24914 17040 27000 17096
rect 24853 17038 27000 17040
rect 24853 17035 24919 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 17125 16692 17191 16693
rect 17125 16688 17172 16692
rect 17236 16690 17242 16692
rect 17125 16632 17130 16688
rect 17125 16628 17172 16632
rect 17236 16630 17282 16690
rect 17236 16628 17242 16630
rect 17125 16627 17191 16628
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 24853 16282 24919 16285
rect 26200 16282 27000 16312
rect 24853 16280 27000 16282
rect 24853 16224 24858 16280
rect 24914 16224 27000 16280
rect 24853 16222 27000 16224
rect 24853 16219 24919 16222
rect 26200 16192 27000 16222
rect 18137 16010 18203 16013
rect 18689 16010 18755 16013
rect 19190 16010 19196 16012
rect 18137 16008 19196 16010
rect 18137 15952 18142 16008
rect 18198 15952 18694 16008
rect 18750 15952 19196 16008
rect 18137 15950 19196 15952
rect 18137 15947 18203 15950
rect 18689 15947 18755 15950
rect 19190 15948 19196 15950
rect 19260 15948 19266 16012
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 13353 15602 13419 15605
rect 13353 15600 13554 15602
rect 13353 15544 13358 15600
rect 13414 15544 13554 15600
rect 13353 15542 13554 15544
rect 13353 15539 13419 15542
rect 13494 15466 13554 15542
rect 13629 15466 13695 15469
rect 13494 15464 13695 15466
rect 13494 15408 13634 15464
rect 13690 15408 13695 15464
rect 13494 15406 13695 15408
rect 13629 15403 13695 15406
rect 24761 15466 24827 15469
rect 26200 15466 27000 15496
rect 24761 15464 27000 15466
rect 24761 15408 24766 15464
rect 24822 15408 27000 15464
rect 24761 15406 27000 15408
rect 24761 15403 24827 15406
rect 26200 15376 27000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 15878 13772 15884 13836
rect 15948 13834 15954 13836
rect 19701 13834 19767 13837
rect 15948 13832 19767 13834
rect 15948 13776 19706 13832
rect 19762 13776 19767 13832
rect 15948 13774 19767 13776
rect 15948 13772 15954 13774
rect 19701 13771 19767 13774
rect 24853 13834 24919 13837
rect 26200 13834 27000 13864
rect 24853 13832 27000 13834
rect 24853 13776 24858 13832
rect 24914 13776 27000 13832
rect 24853 13774 27000 13776
rect 24853 13771 24919 13774
rect 26200 13744 27000 13774
rect 17718 13636 17724 13700
rect 17788 13698 17794 13700
rect 17861 13698 17927 13701
rect 17788 13696 17927 13698
rect 17788 13640 17866 13696
rect 17922 13640 17927 13696
rect 17788 13638 17927 13640
rect 17788 13636 17794 13638
rect 17861 13635 17927 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 13445 13018 13511 13021
rect 13721 13018 13787 13021
rect 13445 13016 13787 13018
rect 13445 12960 13450 13016
rect 13506 12960 13726 13016
rect 13782 12960 13787 13016
rect 13445 12958 13787 12960
rect 13445 12955 13511 12958
rect 13721 12955 13787 12958
rect 15009 13018 15075 13021
rect 15653 13018 15719 13021
rect 15009 13016 15719 13018
rect 15009 12960 15014 13016
rect 15070 12960 15658 13016
rect 15714 12960 15719 13016
rect 15009 12958 15719 12960
rect 15009 12955 15075 12958
rect 15653 12955 15719 12958
rect 24945 13018 25011 13021
rect 26200 13018 27000 13048
rect 24945 13016 27000 13018
rect 24945 12960 24950 13016
rect 25006 12960 27000 13016
rect 24945 12958 27000 12960
rect 24945 12955 25011 12958
rect 26200 12928 27000 12958
rect 7741 12882 7807 12885
rect 15101 12882 15167 12885
rect 16021 12882 16087 12885
rect 7741 12880 16087 12882
rect 7741 12824 7746 12880
rect 7802 12824 15106 12880
rect 15162 12824 16026 12880
rect 16082 12824 16087 12880
rect 7741 12822 16087 12824
rect 7741 12819 7807 12822
rect 15101 12819 15167 12822
rect 16021 12819 16087 12822
rect 16757 12746 16823 12749
rect 17534 12746 17540 12748
rect 16757 12744 17540 12746
rect 16757 12688 16762 12744
rect 16818 12688 17540 12744
rect 16757 12686 17540 12688
rect 16757 12683 16823 12686
rect 17534 12684 17540 12686
rect 17604 12746 17610 12748
rect 18321 12746 18387 12749
rect 17604 12744 18387 12746
rect 17604 12688 18326 12744
rect 18382 12688 18387 12744
rect 17604 12686 18387 12688
rect 17604 12684 17610 12686
rect 18321 12683 18387 12686
rect 21081 12746 21147 12749
rect 25589 12746 25655 12749
rect 21081 12744 25655 12746
rect 21081 12688 21086 12744
rect 21142 12688 25594 12744
rect 25650 12688 25655 12744
rect 21081 12686 25655 12688
rect 21081 12683 21147 12686
rect 25589 12683 25655 12686
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 24945 12202 25011 12205
rect 26200 12202 27000 12232
rect 24945 12200 27000 12202
rect 24945 12144 24950 12200
rect 25006 12144 27000 12200
rect 24945 12142 27000 12144
rect 24945 12139 25011 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24761 11386 24827 11389
rect 26200 11386 27000 11416
rect 24761 11384 27000 11386
rect 24761 11328 24766 11384
rect 24822 11328 27000 11384
rect 24761 11326 27000 11328
rect 24761 11323 24827 11326
rect 26200 11296 27000 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 15929 10706 15995 10709
rect 21449 10706 21515 10709
rect 25037 10706 25103 10709
rect 15929 10704 25103 10706
rect 15929 10648 15934 10704
rect 15990 10648 21454 10704
rect 21510 10648 25042 10704
rect 25098 10648 25103 10704
rect 15929 10646 25103 10648
rect 15929 10643 15995 10646
rect 21449 10643 21515 10646
rect 25037 10643 25103 10646
rect 24669 10570 24735 10573
rect 26200 10570 27000 10600
rect 24669 10568 27000 10570
rect 24669 10512 24674 10568
rect 24730 10512 27000 10568
rect 24669 10510 27000 10512
rect 24669 10507 24735 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 16941 10162 17007 10165
rect 17350 10162 17356 10164
rect 16941 10160 17356 10162
rect 16941 10104 16946 10160
rect 17002 10104 17356 10160
rect 16941 10102 17356 10104
rect 16941 10099 17007 10102
rect 17350 10100 17356 10102
rect 17420 10162 17426 10164
rect 18229 10162 18295 10165
rect 17420 10160 18295 10162
rect 17420 10104 18234 10160
rect 18290 10104 18295 10160
rect 17420 10102 18295 10104
rect 17420 10100 17426 10102
rect 18229 10099 18295 10102
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24761 9754 24827 9757
rect 26200 9754 27000 9784
rect 24761 9752 27000 9754
rect 24761 9696 24766 9752
rect 24822 9696 27000 9752
rect 24761 9694 27000 9696
rect 24761 9691 24827 9694
rect 26200 9664 27000 9694
rect 17493 9482 17559 9485
rect 18321 9482 18387 9485
rect 17493 9480 18387 9482
rect 17493 9424 17498 9480
rect 17554 9424 18326 9480
rect 18382 9424 18387 9480
rect 17493 9422 18387 9424
rect 17493 9419 17559 9422
rect 18321 9419 18387 9422
rect 17493 9346 17559 9349
rect 19057 9346 19123 9349
rect 17493 9344 19123 9346
rect 17493 9288 17498 9344
rect 17554 9288 19062 9344
rect 19118 9288 19123 9344
rect 17493 9286 19123 9288
rect 17493 9283 17559 9286
rect 19057 9283 19123 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 17125 9074 17191 9077
rect 19241 9074 19307 9077
rect 17125 9072 19307 9074
rect 17125 9016 17130 9072
rect 17186 9016 19246 9072
rect 19302 9016 19307 9072
rect 17125 9014 19307 9016
rect 17125 9011 17191 9014
rect 19241 9011 19307 9014
rect 19517 9074 19583 9077
rect 23289 9074 23355 9077
rect 19517 9072 23355 9074
rect 19517 9016 19522 9072
rect 19578 9016 23294 9072
rect 23350 9016 23355 9072
rect 19517 9014 23355 9016
rect 19517 9011 19583 9014
rect 23289 9011 23355 9014
rect 13629 8938 13695 8941
rect 20897 8938 20963 8941
rect 13629 8936 20963 8938
rect 13629 8880 13634 8936
rect 13690 8880 20902 8936
rect 20958 8880 20963 8936
rect 13629 8878 20963 8880
rect 13629 8875 13695 8878
rect 20897 8875 20963 8878
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 3509 8802 3575 8805
rect 0 8800 3575 8802
rect 0 8744 3514 8800
rect 3570 8744 3575 8800
rect 0 8742 3575 8744
rect 0 8712 800 8742
rect 3509 8739 3575 8742
rect 19241 8802 19307 8805
rect 20345 8802 20411 8805
rect 20662 8802 20668 8804
rect 19241 8800 20668 8802
rect 19241 8744 19246 8800
rect 19302 8744 20350 8800
rect 20406 8744 20668 8800
rect 19241 8742 20668 8744
rect 19241 8739 19307 8742
rect 20345 8739 20411 8742
rect 20662 8740 20668 8742
rect 20732 8740 20738 8804
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 13905 8530 13971 8533
rect 17125 8530 17191 8533
rect 13905 8528 17191 8530
rect 13905 8472 13910 8528
rect 13966 8472 17130 8528
rect 17186 8472 17191 8528
rect 13905 8470 17191 8472
rect 13905 8467 13971 8470
rect 17125 8467 17191 8470
rect 12709 8394 12775 8397
rect 13813 8394 13879 8397
rect 20621 8394 20687 8397
rect 12709 8392 20687 8394
rect 12709 8336 12714 8392
rect 12770 8336 13818 8392
rect 13874 8336 20626 8392
rect 20682 8336 20687 8392
rect 12709 8334 20687 8336
rect 12709 8331 12775 8334
rect 13813 8331 13879 8334
rect 20621 8331 20687 8334
rect 14825 8258 14891 8261
rect 19057 8258 19123 8261
rect 14825 8256 19123 8258
rect 14825 8200 14830 8256
rect 14886 8200 19062 8256
rect 19118 8200 19123 8256
rect 14825 8198 19123 8200
rect 14825 8195 14891 8198
rect 19057 8195 19123 8198
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 14457 7850 14523 7853
rect 14774 7850 14780 7852
rect 14457 7848 14780 7850
rect 14457 7792 14462 7848
rect 14518 7792 14780 7848
rect 14457 7790 14780 7792
rect 14457 7787 14523 7790
rect 14774 7788 14780 7790
rect 14844 7788 14850 7852
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 25129 7306 25195 7309
rect 26200 7306 27000 7336
rect 25129 7304 27000 7306
rect 25129 7248 25134 7304
rect 25190 7248 27000 7304
rect 25129 7246 27000 7248
rect 25129 7243 25195 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 14774 6972 14780 7036
rect 14844 7034 14850 7036
rect 14844 6974 15210 7034
rect 14844 6972 14850 6974
rect 15150 6898 15210 6974
rect 15561 6898 15627 6901
rect 15150 6896 15627 6898
rect 15150 6840 15566 6896
rect 15622 6840 15627 6896
rect 15150 6838 15627 6840
rect 15561 6835 15627 6838
rect 21265 6762 21331 6765
rect 23657 6762 23723 6765
rect 21265 6760 23723 6762
rect 21265 6704 21270 6760
rect 21326 6704 23662 6760
rect 23718 6704 23723 6760
rect 21265 6702 23723 6704
rect 21265 6699 21331 6702
rect 23657 6699 23723 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3417 6490 3483 6493
rect 0 6488 3483 6490
rect 0 6432 3422 6488
rect 3478 6432 3483 6488
rect 0 6430 3483 6432
rect 0 6400 800 6430
rect 3417 6427 3483 6430
rect 24761 6490 24827 6493
rect 26200 6490 27000 6520
rect 24761 6488 27000 6490
rect 24761 6432 24766 6488
rect 24822 6432 27000 6488
rect 24761 6430 27000 6432
rect 24761 6427 24827 6430
rect 26200 6400 27000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 20437 5810 20503 5813
rect 22185 5810 22251 5813
rect 20437 5808 22251 5810
rect 20437 5752 20442 5808
rect 20498 5752 22190 5808
rect 22246 5752 22251 5808
rect 20437 5750 22251 5752
rect 20437 5747 20503 5750
rect 22185 5747 22251 5750
rect 23289 5674 23355 5677
rect 26200 5674 27000 5704
rect 23289 5672 27000 5674
rect 23289 5616 23294 5672
rect 23350 5616 27000 5672
rect 23289 5614 27000 5616
rect 23289 5611 23355 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 18873 5402 18939 5405
rect 22461 5402 22527 5405
rect 18873 5400 22527 5402
rect 18873 5344 18878 5400
rect 18934 5344 22466 5400
rect 22522 5344 22527 5400
rect 18873 5342 22527 5344
rect 18873 5339 18939 5342
rect 22461 5339 22527 5342
rect 21909 5130 21975 5133
rect 21909 5128 24226 5130
rect 21909 5072 21914 5128
rect 21970 5072 24226 5128
rect 21909 5070 24226 5072
rect 21909 5067 21975 5070
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24166 4858 24226 5070
rect 26200 4858 27000 4888
rect 24166 4798 27000 4858
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4178 800 4208
rect 3877 4178 3943 4181
rect 0 4176 3943 4178
rect 0 4120 3882 4176
rect 3938 4120 3943 4176
rect 0 4118 3943 4120
rect 0 4088 800 4118
rect 3877 4115 3943 4118
rect 12433 4178 12499 4181
rect 15878 4178 15884 4180
rect 12433 4176 15884 4178
rect 12433 4120 12438 4176
rect 12494 4120 15884 4176
rect 12433 4118 15884 4120
rect 12433 4115 12499 4118
rect 15878 4116 15884 4118
rect 15948 4116 15954 4180
rect 22829 4042 22895 4045
rect 26200 4042 27000 4072
rect 22829 4040 27000 4042
rect 22829 3984 22834 4040
rect 22890 3984 27000 4040
rect 22829 3982 27000 3984
rect 22829 3979 22895 3982
rect 26200 3952 27000 3982
rect 18597 3906 18663 3909
rect 22277 3906 22343 3909
rect 18597 3904 22343 3906
rect 18597 3848 18602 3904
rect 18658 3848 22282 3904
rect 22338 3848 22343 3904
rect 18597 3846 22343 3848
rect 18597 3843 18663 3846
rect 22277 3843 22343 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 20713 3364 20779 3365
rect 20662 3362 20668 3364
rect 20622 3302 20668 3362
rect 20732 3360 20779 3364
rect 20774 3304 20779 3360
rect 20662 3300 20668 3302
rect 20732 3300 20779 3304
rect 20713 3299 20779 3300
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 20069 3226 20135 3229
rect 26200 3226 27000 3256
rect 20069 3224 27000 3226
rect 20069 3168 20074 3224
rect 20130 3168 27000 3224
rect 20069 3166 27000 3168
rect 20069 3163 20135 3166
rect 26200 3136 27000 3166
rect 13169 3090 13235 3093
rect 17166 3090 17172 3092
rect 13169 3088 17172 3090
rect 13169 3032 13174 3088
rect 13230 3032 17172 3088
rect 13169 3030 17172 3032
rect 13169 3027 13235 3030
rect 17166 3028 17172 3030
rect 17236 3028 17242 3092
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 12893 2546 12959 2549
rect 15694 2546 15700 2548
rect 12893 2544 15700 2546
rect 12893 2488 12898 2544
rect 12954 2488 15700 2544
rect 12893 2486 15700 2488
rect 12893 2483 12959 2486
rect 15694 2484 15700 2486
rect 15764 2484 15770 2548
rect 21817 2410 21883 2413
rect 26200 2410 27000 2440
rect 21817 2408 27000 2410
rect 21817 2352 21822 2408
rect 21878 2352 27000 2408
rect 21817 2350 27000 2352
rect 21817 2347 21883 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 800 1806
rect 3417 1803 3483 1806
rect 22093 1594 22159 1597
rect 26200 1594 27000 1624
rect 22093 1592 27000 1594
rect 22093 1536 22098 1592
rect 22154 1536 27000 1592
rect 22093 1534 27000 1536
rect 22093 1531 22159 1534
rect 26200 1504 27000 1534
rect 25129 778 25195 781
rect 26200 778 27000 808
rect 25129 776 27000 778
rect 25129 720 25134 776
rect 25190 720 27000 776
rect 25129 718 27000 720
rect 25129 715 25195 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 19196 41652 19260 41716
rect 19932 41380 19996 41444
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 17356 27976 17420 27980
rect 17356 27920 17370 27976
rect 17370 27920 17420 27976
rect 17356 27916 17420 27920
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 16804 25936 16868 25940
rect 16804 25880 16818 25936
rect 16818 25880 16868 25936
rect 16804 25876 16868 25880
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 14780 25120 14844 25124
rect 14780 25064 14830 25120
rect 14830 25064 14844 25120
rect 14780 25060 14844 25064
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 15700 24244 15764 24308
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 20852 22476 20916 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 17540 19348 17604 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 20852 18668 20916 18732
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 17724 18260 17788 18324
rect 19932 18124 19996 18188
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 16804 17444 16868 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 17172 16688 17236 16692
rect 17172 16632 17186 16688
rect 17186 16632 17236 16688
rect 17172 16628 17236 16632
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 19196 15948 19260 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 15884 13772 15948 13836
rect 17724 13636 17788 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 17540 12684 17604 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 17356 10100 17420 10164
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 20668 8740 20732 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 14780 7788 14844 7852
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 14780 6972 14844 7036
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 15884 4116 15948 4180
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 20668 3360 20732 3364
rect 20668 3304 20718 3360
rect 20718 3304 20732 3360
rect 20668 3300 20732 3304
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 17172 3028 17236 3092
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 15700 2484 15764 2548
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 19195 41716 19261 41717
rect 19195 41652 19196 41716
rect 19260 41652 19261 41716
rect 19195 41651 19261 41652
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17355 27980 17421 27981
rect 17355 27916 17356 27980
rect 17420 27916 17421 27980
rect 17355 27915 17421 27916
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 16803 25940 16869 25941
rect 16803 25876 16804 25940
rect 16868 25876 16869 25940
rect 16803 25875 16869 25876
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 14779 25124 14845 25125
rect 14779 25060 14780 25124
rect 14844 25060 14845 25124
rect 14779 25059 14845 25060
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 14782 7853 14842 25059
rect 15699 24308 15765 24309
rect 15699 24244 15700 24308
rect 15764 24244 15765 24308
rect 15699 24243 15765 24244
rect 14779 7852 14845 7853
rect 14779 7788 14780 7852
rect 14844 7788 14845 7852
rect 14779 7787 14845 7788
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 14782 7037 14842 7787
rect 14779 7036 14845 7037
rect 14779 6972 14780 7036
rect 14844 6972 14845 7036
rect 14779 6971 14845 6972
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 15702 2549 15762 24243
rect 16806 17509 16866 25875
rect 16803 17508 16869 17509
rect 16803 17444 16804 17508
rect 16868 17444 16869 17508
rect 16803 17443 16869 17444
rect 17171 16692 17237 16693
rect 17171 16628 17172 16692
rect 17236 16628 17237 16692
rect 17171 16627 17237 16628
rect 15883 13836 15949 13837
rect 15883 13772 15884 13836
rect 15948 13772 15949 13836
rect 15883 13771 15949 13772
rect 15886 4181 15946 13771
rect 15883 4180 15949 4181
rect 15883 4116 15884 4180
rect 15948 4116 15949 4180
rect 15883 4115 15949 4116
rect 17174 3093 17234 16627
rect 17358 10165 17418 27915
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17542 12749 17602 19347
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17723 18324 17789 18325
rect 17723 18260 17724 18324
rect 17788 18260 17789 18324
rect 17723 18259 17789 18260
rect 17726 13701 17786 18259
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 19198 16013 19258 41651
rect 19931 41444 19997 41445
rect 19931 41380 19932 41444
rect 19996 41380 19997 41444
rect 19931 41379 19997 41380
rect 19934 18189 19994 41379
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 20851 22540 20917 22541
rect 20851 22476 20852 22540
rect 20916 22476 20917 22540
rect 20851 22475 20917 22476
rect 20854 18733 20914 22475
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 20851 18732 20917 18733
rect 20851 18668 20852 18732
rect 20916 18668 20917 18732
rect 20851 18667 20917 18668
rect 19931 18188 19997 18189
rect 19931 18124 19932 18188
rect 19996 18124 19997 18188
rect 19931 18123 19997 18124
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 19195 16012 19261 16013
rect 19195 15948 19196 16012
rect 19260 15948 19261 16012
rect 19195 15947 19261 15948
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17723 13700 17789 13701
rect 17723 13636 17724 13700
rect 17788 13636 17789 13700
rect 17723 13635 17789 13636
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17539 12748 17605 12749
rect 17539 12684 17540 12748
rect 17604 12684 17605 12748
rect 17539 12683 17605 12684
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17355 10164 17421 10165
rect 17355 10100 17356 10164
rect 17420 10100 17421 10164
rect 17355 10099 17421 10100
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 20667 8804 20733 8805
rect 20667 8740 20668 8804
rect 20732 8740 20733 8804
rect 20667 8739 20733 8740
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 20670 3365 20730 8739
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 20667 3364 20733 3365
rect 20667 3300 20668 3364
rect 20732 3300 20733 3364
rect 20667 3299 20733 3300
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17171 3092 17237 3093
rect 17171 3028 17172 3092
rect 17236 3028 17237 3092
rect 17171 3027 17237 3028
rect 15699 2548 15765 2549
rect 15699 2484 15700 2548
rect 15764 2484 15765 2548
rect 15699 2483 15765 2484
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _108_
timestamp 1676037725
transform 1 0 13432 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_
timestamp 1676037725
transform 1 0 18400 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1676037725
transform 1 0 12880 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1676037725
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1676037725
transform 1 0 21620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1676037725
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1676037725
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 16928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1676037725
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 14904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1676037725
transform 1 0 5152 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 6624 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 7544 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 8280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 9384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 11408 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 15916 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6440 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7268 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6348 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15180 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9752 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1676037725
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14720 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 14444 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 12512 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 10212 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 14260 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 11592 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 12144 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 10304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 7544 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8096 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17204 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17480 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 14260 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 14628 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 15364 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 22172 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 19964 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1676037725
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1676037725
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_238
timestamp 1676037725
transform 1 0 23000 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1676037725
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1676037725
transform 1 0 6532 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1676037725
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1676037725
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_259
timestamp 1676037725
transform 1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1676037725
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_62
timestamp 1676037725
transform 1 0 6808 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_74
timestamp 1676037725
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_86
timestamp 1676037725
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_98
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1676037725
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1676037725
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1676037725
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1676037725
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_243
timestamp 1676037725
transform 1 0 23460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1676037725
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_150
timestamp 1676037725
transform 1 0 14904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1676037725
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1676037725
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_116
timestamp 1676037725
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_128
timestamp 1676037725
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1676037725
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1676037725
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_203
timestamp 1676037725
transform 1 0 19780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1676037725
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_144
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_152
timestamp 1676037725
transform 1 0 15088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1676037725
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_198
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1676037725
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1676037725
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1676037725
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_224
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1676037725
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1676037725
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_124
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1676037725
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_176
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_200
timestamp 1676037725
transform 1 0 19504 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1676037725
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1676037725
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_179
timestamp 1676037725
transform 1 0 17572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_203
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_226
timestamp 1676037725
transform 1 0 21896 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_124
timestamp 1676037725
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1676037725
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_148
timestamp 1676037725
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_180
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_197
timestamp 1676037725
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_201
timestamp 1676037725
transform 1 0 19596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_113
timestamp 1676037725
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_183
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1676037725
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_139
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1676037725
transform 1 0 17296 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1676037725
transform 1 0 19504 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_167
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_224
timestamp 1676037725
transform 1 0 21712 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_120
timestamp 1676037725
transform 1 0 12144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_146
timestamp 1676037725
transform 1 0 14536 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_154
timestamp 1676037725
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1676037725
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1676037725
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1676037725
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1676037725
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_231
timestamp 1676037725
transform 1 0 22356 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_258
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_87
timestamp 1676037725
transform 1 0 9108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1676037725
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_153
timestamp 1676037725
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1676037725
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_232
timestamp 1676037725
transform 1 0 22448 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_238
timestamp 1676037725
transform 1 0 23000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_259
timestamp 1676037725
transform 1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1676037725
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1676037725
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp 1676037725
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1676037725
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1676037725
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207
timestamp 1676037725
transform 1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_57
timestamp 1676037725
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1676037725
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1676037725
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1676037725
transform 1 0 21620 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_258
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1676037725
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1676037725
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1676037725
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_223
timestamp 1676037725
transform 1 0 21620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_258
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_96
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_108
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_124
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1676037725
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_161
timestamp 1676037725
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_79
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_91
timestamp 1676037725
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1676037725
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1676037725
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1676037725
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_110
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1676037725
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1676037725
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1676037725
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_224
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1676037725
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1676037725
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1676037725
transform 1 0 17940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_206
timestamp 1676037725
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_212
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1676037725
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_157
timestamp 1676037725
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_161
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_172
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_180
timestamp 1676037725
transform 1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_219
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_225
timestamp 1676037725
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1676037725
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_133
timestamp 1676037725
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_146
timestamp 1676037725
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1676037725
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_203
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1676037725
transform 1 0 20608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_129
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1676037725
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1676037725
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_143
timestamp 1676037725
transform 1 0 14260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_182
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1676037725
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1676037725
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_95
timestamp 1676037725
transform 1 0 9844 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_231
timestamp 1676037725
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_61
timestamp 1676037725
transform 1 0 6716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_100
timestamp 1676037725
transform 1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_185
timestamp 1676037725
transform 1 0 18124 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1676037725
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_98
timestamp 1676037725
transform 1 0 10120 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_126
timestamp 1676037725
transform 1 0 12696 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1676037725
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1676037725
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_95
timestamp 1676037725
transform 1 0 9844 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1676037725
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_154
timestamp 1676037725
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1676037725
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_204
timestamp 1676037725
transform 1 0 19872 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1676037725
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_212
timestamp 1676037725
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_96
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_119
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_163
timestamp 1676037725
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_175
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1676037725
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_216
timestamp 1676037725
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1676037725
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1676037725
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_195
timestamp 1676037725
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_207
timestamp 1676037725
transform 1 0 20148 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1676037725
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_232
timestamp 1676037725
transform 1 0 22448 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_260
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_105
timestamp 1676037725
transform 1 0 10764 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_126
timestamp 1676037725
transform 1 0 12696 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_219
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1676037725
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_112
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_152
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_158
timestamp 1676037725
transform 1 0 15640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_190
timestamp 1676037725
transform 1 0 18584 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1676037725
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_218
timestamp 1676037725
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1676037725
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_128
timestamp 1676037725
transform 1 0 12880 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_134
timestamp 1676037725
transform 1 0 13432 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1676037725
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_174
timestamp 1676037725
transform 1 0 17112 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_191
timestamp 1676037725
transform 1 0 18676 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_199
timestamp 1676037725
transform 1 0 19412 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_152
timestamp 1676037725
transform 1 0 15088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_166
timestamp 1676037725
transform 1 0 16376 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_178
timestamp 1676037725
transform 1 0 17480 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_219
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1676037725
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_87
timestamp 1676037725
transform 1 0 9108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1676037725
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_129
timestamp 1676037725
transform 1 0 12972 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1676037725
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_203
timestamp 1676037725
transform 1 0 19780 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_211
timestamp 1676037725
transform 1 0 20516 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1676037725
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_265
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_122
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_128
timestamp 1676037725
transform 1 0 12880 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_162
timestamp 1676037725
transform 1 0 16008 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_174
timestamp 1676037725
transform 1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_182
timestamp 1676037725
transform 1 0 17848 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1676037725
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1676037725
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_225
timestamp 1676037725
transform 1 0 21804 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1676037725
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1676037725
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_133
timestamp 1676037725
transform 1 0 13340 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_145
timestamp 1676037725
transform 1 0 14444 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_157
timestamp 1676037725
transform 1 0 15548 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1676037725
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1676037725
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1676037725
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1676037725
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_147
timestamp 1676037725
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_157
timestamp 1676037725
transform 1 0 15548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_170
timestamp 1676037725
transform 1 0 16744 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1676037725
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_205
timestamp 1676037725
transform 1 0 19964 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_231
timestamp 1676037725
transform 1 0 22356 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1676037725
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1676037725
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1676037725
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_188
timestamp 1676037725
transform 1 0 18400 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_206
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1676037725
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_129
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1676037725
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_162
timestamp 1676037725
transform 1 0 16008 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_170
timestamp 1676037725
transform 1 0 16744 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1676037725
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_87
timestamp 1676037725
transform 1 0 9108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_99
timestamp 1676037725
transform 1 0 10212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1676037725
transform 1 0 13524 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_154
timestamp 1676037725
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1676037725
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_201
timestamp 1676037725
transform 1 0 19596 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_212
timestamp 1676037725
transform 1 0 20608 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_218
timestamp 1676037725
transform 1 0 21160 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1676037725
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1676037725
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_114
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_154
timestamp 1676037725
transform 1 0 15272 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_166
timestamp 1676037725
transform 1 0 16376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1676037725
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_208
timestamp 1676037725
transform 1 0 20240 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_232
timestamp 1676037725
transform 1 0 22448 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1676037725
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_131
timestamp 1676037725
transform 1 0 13156 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_153
timestamp 1676037725
transform 1 0 15180 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_180
timestamp 1676037725
transform 1 0 17664 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_192
timestamp 1676037725
transform 1 0 18768 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_204
timestamp 1676037725
transform 1 0 19872 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1676037725
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_251
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_259
timestamp 1676037725
transform 1 0 24932 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1676037725
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_232
timestamp 1676037725
transform 1 0 22448 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_175
timestamp 1676037725
transform 1 0 17204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_196
timestamp 1676037725
transform 1 0 19136 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1676037725
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1676037725
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_216
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_228
timestamp 1676037725
transform 1 0 22080 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1676037725
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1676037725
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1676037725
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1676037725
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1676037725
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1676037725
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_158
timestamp 1676037725
transform 1 0 15640 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_170
timestamp 1676037725
transform 1 0 16744 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_182
timestamp 1676037725
transform 1 0 17848 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1676037725
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1676037725
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_248
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_257
timestamp 1676037725
transform 1 0 24748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1676037725
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1676037725
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_257
timestamp 1676037725
transform 1 0 24748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_265
timestamp 1676037725
transform 1 0 25484 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_106
timestamp 1676037725
transform 1 0 10856 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_118
timestamp 1676037725
transform 1 0 11960 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_130
timestamp 1676037725
transform 1 0 13064 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_138
timestamp 1676037725
transform 1 0 13800 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_265
timestamp 1676037725
transform 1 0 25484 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_100
timestamp 1676037725
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_112
timestamp 1676037725
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_124
timestamp 1676037725
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1676037725
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_259
timestamp 1676037725
transform 1 0 24932 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1676037725
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_230
timestamp 1676037725
transform 1 0 22264 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_242
timestamp 1676037725
transform 1 0 23368 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1676037725
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1676037725
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_257
timestamp 1676037725
transform 1 0 24748 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_119
timestamp 1676037725
transform 1 0 12052 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_131
timestamp 1676037725
transform 1 0 13156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_265
timestamp 1676037725
transform 1 0 25484 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_127
timestamp 1676037725
transform 1 0 12788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_131
timestamp 1676037725
transform 1 0 13156 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1676037725
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_157
timestamp 1676037725
transform 1 0 15548 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_179
timestamp 1676037725
transform 1 0 17572 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1676037725
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_75
timestamp 1676037725
transform 1 0 8004 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_84
timestamp 1676037725
transform 1 0 8832 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_96
timestamp 1676037725
transform 1 0 9936 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 1676037725
transform 1 0 12052 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_141
timestamp 1676037725
transform 1 0 14076 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1676037725
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_117
timestamp 1676037725
transform 1 0 11868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1676037725
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1676037725
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_164
timestamp 1676037725
transform 1 0 16192 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_176
timestamp 1676037725
transform 1 0 17296 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1676037725
transform 1 0 18400 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1676037725
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_96
timestamp 1676037725
transform 1 0 9936 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_108
timestamp 1676037725
transform 1 0 11040 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_103
timestamp 1676037725
transform 1 0 10580 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1676037725
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1676037725
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_80
timestamp 1676037725
transform 1 0 8464 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_92
timestamp 1676037725
transform 1 0 9568 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_104
timestamp 1676037725
transform 1 0 10672 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_265
timestamp 1676037725
transform 1 0 25484 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_105
timestamp 1676037725
transform 1 0 10764 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1676037725
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_116
timestamp 1676037725
transform 1 0 11776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_128
timestamp 1676037725
transform 1 0 12880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_259
timestamp 1676037725
transform 1 0 24932 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1676037725
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_69
timestamp 1676037725
transform 1 0 7452 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_76
timestamp 1676037725
transform 1 0 8096 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_89
timestamp 1676037725
transform 1 0 9292 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_94
timestamp 1676037725
transform 1 0 9752 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1676037725
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1676037725
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_130
timestamp 1676037725
transform 1 0 13064 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_138
timestamp 1676037725
transform 1 0 13800 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1676037725
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1676037725
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_257
timestamp 1676037725
transform 1 0 24748 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1676037725
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1676037725
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1676037725
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_257
timestamp 1676037725
transform 1 0 24748 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_63
timestamp 1676037725
transform 1 0 6900 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_75
timestamp 1676037725
transform 1 0 8004 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_87
timestamp 1676037725
transform 1 0 9108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_99
timestamp 1676037725
transform 1 0 10212 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1676037725
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_257
timestamp 1676037725
transform 1 0 24748 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1676037725
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1676037725
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1676037725
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_43
timestamp 1676037725
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1676037725
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_249
timestamp 1676037725
transform 1 0 24012 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1676037725
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1676037725
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_47
timestamp 1676037725
transform 1 0 5428 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_59
timestamp 1676037725
transform 1 0 6532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_76
timestamp 1676037725
transform 1 0 8096 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_237
timestamp 1676037725
transform 1 0 22908 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_259
timestamp 1676037725
transform 1 0 24932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1676037725
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_106
timestamp 1676037725
transform 1 0 10856 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_136
timestamp 1676037725
transform 1 0 13616 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_146
timestamp 1676037725
transform 1 0 14536 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_174
timestamp 1676037725
transform 1 0 17112 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1676037725
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_209
timestamp 1676037725
transform 1 0 20332 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_239
timestamp 1676037725
transform 1 0 23092 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_244
timestamp 1676037725
transform 1 0 23552 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_259
timestamp 1676037725
transform 1 0 24932 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_265
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1676037725
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 11040 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 24288 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 23000 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 20700 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 22080 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 20792 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 20056 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 17480 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 22172 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20424 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 6624 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 9384 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 10764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19964 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17940 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16744 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17296 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20516 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20424 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13248 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10488 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10396 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9200 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11960 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10856 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8740 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9292 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12420 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9936 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23092 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17664 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22080 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 19688 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19320 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22172 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1676037725
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 17940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 19688 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 23368 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20976 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19780 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 18584 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13616 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14720 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15916 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 9844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10304 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13616 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17756 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18400 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 23368 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20884 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22724 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1676037725
transform 1 0 17020 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 9890 29070 9890 29070 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9706 41582 9706 41582 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9246 42670 9246 42670 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9062 34170 9062 34170 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8280 37978 8280 37978 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 8970 19210 8970 19210 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 15226 12750 15226 12750 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 6831 13226 6831 13226 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 9660 15538 9660 15538 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 8096 17714 8096 17714 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal2 13662 14654 13662 14654 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13524 10098 13524 10098 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 9890 13362 9890 13362 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 8326 20366 8326 20366 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 13938 16082 13938 16082 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 11822 18326 11822 18326 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 10994 20400 10994 20400 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 9890 17714 9890 17714 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 13478 25721 13478 25721 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 10442 25330 10442 25330 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 14306 8840 14306 8840 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9154 17510 9154 17510 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9062 30702 9062 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 14030 9146 14030 9146 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14582 10914 14582 10914 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13708 12614 13708 12614 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9522 12784 9522 12784 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11132 14994 11132 14994 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11270 15062 11270 15062 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9338 12954 9338 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10442 12920 10442 12920 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10120 16932 10120 16932 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 16652 8058 16652 8058 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8740 17578 8740 17578 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7774 17850 7774 17850 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13386 8942 13386 8942 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15226 10200 15226 10200 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13570 11118 13570 11118 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12880 14246 12880 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 10718 10574 10718 10574 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10626 11696 10626 11696 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9798 13430 9798 13430 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11500 12682 11500 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9154 17510 9154 17510 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13570 13158 13570 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 20570 9982 20570 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 33966 9200 33966 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15364 10778 15364 10778 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13754 10880 13754 10880 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12558 11458 12558 11458 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13110 15946 13110 15946 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12098 13498 12098 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11132 16490 11132 16490 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10350 20502 10350 20502 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12788 20570 12788 20570 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9660 16422 9660 16422 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14306 11866 14306 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10488 25466 10488 25466 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 37842 9200 37842 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13478 16218 13478 16218 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12512 15334 12512 15334 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12374 15402 12374 15402 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12144 18394 12144 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11546 21386 11546 21386 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11684 19108 11684 19108 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10442 18938 10442 18938 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 13294 25806 13294 25806 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 21658 10350 21658 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 10718 43146 10718 43146 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 11040 44166 11040 44166 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 10856 41786 10856 41786 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 14651 45866 14651 45866 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9568 44778 9568 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 10672 46682 10672 46682 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 10212 42738 10212 42738 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 13685 46138 13685 46138 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10166 45050 10166 45050 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9200 44370 9200 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 9568 50286 9568 50286 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 13133 46954 13133 46954 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 7912 50422 7912 50422 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 8510 48892 8510 48892 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 12374 47294 12374 47294 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25622 51986 25622 51986 0 ccff_head
rlabel metal2 1518 2438 1518 2438 0 ccff_head_0
rlabel metal3 25768 748 25768 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal2 22218 26197 22218 26197 0 chanx_right_in[0]
rlabel metal2 25346 34391 25346 34391 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal2 25346 35989 25346 35989 0 chanx_right_in[12]
rlabel metal2 25162 36703 25162 36703 0 chanx_right_in[13]
rlabel metal2 25162 37655 25162 37655 0 chanx_right_in[14]
rlabel via2 25346 38301 25346 38301 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal2 25346 39967 25346 39967 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25162 41531 25162 41531 0 chanx_right_in[19]
rlabel metal2 25346 26061 25346 26061 0 chanx_right_in[1]
rlabel metal2 25162 42483 25162 42483 0 chanx_right_in[20]
rlabel metal2 25162 43231 25162 43231 0 chanx_right_in[21]
rlabel metal1 24978 44370 24978 44370 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25162 48059 25162 48059 0 chanx_right_in[27]
rlabel metal2 25162 49011 25162 49011 0 chanx_right_in[28]
rlabel metal1 24702 49810 24702 49810 0 chanx_right_in[29]
rlabel metal2 24058 27013 24058 27013 0 chanx_right_in[2]
rlabel metal1 24886 29138 24886 29138 0 chanx_right_in[3]
rlabel metal1 25392 30702 25392 30702 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel metal2 25346 31127 25346 31127 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal1 25392 33490 25392 33490 0 chanx_right_in[8]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[9]
rlabel metal2 22126 1751 22126 1751 0 chanx_right_out[0]
rlabel metal2 24794 9061 24794 9061 0 chanx_right_out[10]
rlabel metal2 24702 10013 24702 10013 0 chanx_right_out[11]
rlabel metal2 24794 10965 24794 10965 0 chanx_right_out[12]
rlabel metal3 25676 12172 25676 12172 0 chanx_right_out[13]
rlabel metal3 25676 12988 25676 12988 0 chanx_right_out[14]
rlabel metal1 24104 13838 24104 13838 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal2 24794 15181 24794 15181 0 chanx_right_out[17]
rlabel metal1 24380 16490 24380 16490 0 chanx_right_out[18]
rlabel metal1 24104 17238 24104 17238 0 chanx_right_out[19]
rlabel metal3 24112 2380 24112 2380 0 chanx_right_out[1]
rlabel metal1 24380 17714 24380 17714 0 chanx_right_out[20]
rlabel metal2 24794 17901 24794 17901 0 chanx_right_out[21]
rlabel metal2 23874 19159 23874 19159 0 chanx_right_out[22]
rlabel metal1 21712 20366 21712 20366 0 chanx_right_out[23]
rlabel metal1 21666 21454 21666 21454 0 chanx_right_out[24]
rlabel metal1 24518 20842 24518 20842 0 chanx_right_out[25]
rlabel metal1 24104 22678 24104 22678 0 chanx_right_out[26]
rlabel metal1 23460 23154 23460 23154 0 chanx_right_out[27]
rlabel metal2 24794 23477 24794 23477 0 chanx_right_out[28]
rlabel metal3 25676 25228 25676 25228 0 chanx_right_out[29]
rlabel metal1 16790 5780 16790 5780 0 chanx_right_out[2]
rlabel metal2 20470 6392 20470 6392 0 chanx_right_out[3]
rlabel metal2 21942 6205 21942 6205 0 chanx_right_out[4]
rlabel metal2 23322 6477 23322 6477 0 chanx_right_out[5]
rlabel metal2 24794 5797 24794 5797 0 chanx_right_out[6]
rlabel metal2 25162 6817 25162 6817 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal2 1886 2438 1886 2438 0 chany_bottom_in_0[0]
rlabel metal2 5566 1622 5566 1622 0 chany_bottom_in_0[10]
rlabel metal1 6348 4114 6348 4114 0 chany_bottom_in_0[11]
rlabel metal2 6302 1554 6302 1554 0 chany_bottom_in_0[12]
rlabel metal1 6808 3502 6808 3502 0 chany_bottom_in_0[13]
rlabel metal1 7176 3026 7176 3026 0 chany_bottom_in_0[14]
rlabel metal2 7406 1588 7406 1588 0 chany_bottom_in_0[15]
rlabel metal2 7774 1588 7774 1588 0 chany_bottom_in_0[16]
rlabel metal2 8142 823 8142 823 0 chany_bottom_in_0[17]
rlabel metal1 8234 3026 8234 3026 0 chany_bottom_in_0[18]
rlabel metal1 8740 3026 8740 3026 0 chany_bottom_in_0[19]
rlabel metal2 2254 2132 2254 2132 0 chany_bottom_in_0[1]
rlabel metal2 9246 1894 9246 1894 0 chany_bottom_in_0[20]
rlabel metal1 9752 3502 9752 3502 0 chany_bottom_in_0[21]
rlabel metal2 9982 1554 9982 1554 0 chany_bottom_in_0[22]
rlabel metal1 10120 3026 10120 3026 0 chany_bottom_in_0[23]
rlabel metal1 10672 3502 10672 3502 0 chany_bottom_in_0[24]
rlabel metal1 10810 3026 10810 3026 0 chany_bottom_in_0[25]
rlabel metal1 11592 2958 11592 2958 0 chany_bottom_in_0[26]
rlabel metal1 11500 3026 11500 3026 0 chany_bottom_in_0[27]
rlabel metal2 12190 1588 12190 1588 0 chany_bottom_in_0[28]
rlabel metal2 12558 2166 12558 2166 0 chany_bottom_in_0[29]
rlabel metal2 2622 1894 2622 1894 0 chany_bottom_in_0[2]
rlabel metal2 2990 1622 2990 1622 0 chany_bottom_in_0[3]
rlabel metal1 3404 2958 3404 2958 0 chany_bottom_in_0[4]
rlabel metal2 3726 1299 3726 1299 0 chany_bottom_in_0[5]
rlabel metal1 4232 4114 4232 4114 0 chany_bottom_in_0[6]
rlabel metal2 4462 2132 4462 2132 0 chany_bottom_in_0[7]
rlabel metal1 4876 3502 4876 3502 0 chany_bottom_in_0[8]
rlabel metal2 5198 1860 5198 1860 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal1 17894 3094 17894 3094 0 chany_bottom_out_0[10]
rlabel metal1 18446 2890 18446 2890 0 chany_bottom_out_0[11]
rlabel metal2 17342 1503 17342 1503 0 chany_bottom_out_0[12]
rlabel metal1 18860 3570 18860 3570 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal1 22310 2482 22310 2482 0 chany_bottom_out_0[15]
rlabel metal1 19366 3638 19366 3638 0 chany_bottom_out_0[16]
rlabel metal1 20470 3434 20470 3434 0 chany_bottom_out_0[17]
rlabel metal1 20332 3366 20332 3366 0 chany_bottom_out_0[18]
rlabel metal2 19918 1435 19918 1435 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal2 20286 1761 20286 1761 0 chany_bottom_out_0[20]
rlabel metal1 20976 2890 20976 2890 0 chany_bottom_out_0[21]
rlabel metal2 21022 2336 21022 2336 0 chany_bottom_out_0[22]
rlabel metal2 21390 1826 21390 1826 0 chany_bottom_out_0[23]
rlabel metal2 21758 823 21758 823 0 chany_bottom_out_0[24]
rlabel metal2 22126 1095 22126 1095 0 chany_bottom_out_0[25]
rlabel metal2 22494 1761 22494 1761 0 chany_bottom_out_0[26]
rlabel metal2 22862 1554 22862 1554 0 chany_bottom_out_0[27]
rlabel metal2 23230 1690 23230 1690 0 chany_bottom_out_0[28]
rlabel metal1 23460 9486 23460 9486 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal1 16238 2822 16238 2822 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16606 2958 16606 2958 0 chany_bottom_out_0[8]
rlabel metal1 16790 4046 16790 4046 0 chany_bottom_out_0[9]
rlabel metal1 18630 13294 18630 13294 0 clknet_0_prog_clk
rlabel metal2 6394 14688 6394 14688 0 clknet_4_0_0_prog_clk
rlabel metal1 6670 48586 6670 48586 0 clknet_4_10_0_prog_clk
rlabel metal1 14490 32334 14490 32334 0 clknet_4_11_0_prog_clk
rlabel metal1 18124 20570 18124 20570 0 clknet_4_12_0_prog_clk
rlabel metal1 23276 21522 23276 21522 0 clknet_4_13_0_prog_clk
rlabel metal1 19504 32402 19504 32402 0 clknet_4_14_0_prog_clk
rlabel metal1 20010 43758 20010 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 13294 12886 13294 12886 0 clknet_4_1_0_prog_clk
rlabel metal1 6624 18734 6624 18734 0 clknet_4_2_0_prog_clk
rlabel via1 12742 21522 12742 21522 0 clknet_4_3_0_prog_clk
rlabel metal2 16882 4896 16882 4896 0 clknet_4_4_0_prog_clk
rlabel metal1 22954 12750 22954 12750 0 clknet_4_5_0_prog_clk
rlabel metal1 18906 16626 18906 16626 0 clknet_4_6_0_prog_clk
rlabel metal1 20102 19890 20102 19890 0 clknet_4_7_0_prog_clk
rlabel metal1 13386 29172 13386 29172 0 clknet_4_8_0_prog_clk
rlabel metal2 15134 29342 15134 29342 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal1 4140 53618 4140 53618 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 5198 55158 5198 55158 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6578 54920 6578 54920 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 13662 56236 13662 56236 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal1 9614 54094 9614 54094 0 gfpga_pad_io_soc_out[1]
rlabel metal1 10718 53652 10718 53652 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54162 19228 54162 0 isol_n
rlabel metal1 22448 43826 22448 43826 0 net1
rlabel metal1 22310 31790 22310 31790 0 net10
rlabel metal1 22172 22950 22172 22950 0 net100
rlabel metal2 23782 22406 23782 22406 0 net101
rlabel metal2 22678 23290 22678 23290 0 net102
rlabel metal2 23966 23970 23966 23970 0 net103
rlabel metal1 21574 25160 21574 25160 0 net104
rlabel metal2 16146 4828 16146 4828 0 net105
rlabel metal1 17710 6800 17710 6800 0 net106
rlabel metal1 13800 6290 13800 6290 0 net107
rlabel metal2 20746 7888 20746 7888 0 net108
rlabel metal1 18722 10710 18722 10710 0 net109
rlabel metal1 23230 31790 23230 31790 0 net11
rlabel metal1 24380 6290 24380 6290 0 net110
rlabel metal2 15778 7684 15778 7684 0 net111
rlabel via2 20930 8925 20930 8925 0 net112
rlabel via2 19734 13821 19734 13821 0 net113
rlabel metal1 18630 3026 18630 3026 0 net114
rlabel metal1 19274 2414 19274 2414 0 net115
rlabel metal1 18216 4590 18216 4590 0 net116
rlabel metal1 19688 3502 19688 3502 0 net117
rlabel metal1 17986 4114 17986 4114 0 net118
rlabel metal1 22034 2482 22034 2482 0 net119
rlabel metal1 25070 32980 25070 32980 0 net12
rlabel metal1 19734 4590 19734 4590 0 net120
rlabel metal1 21022 3502 21022 3502 0 net121
rlabel metal2 22724 13906 22724 13906 0 net122
rlabel metal1 22586 17034 22586 17034 0 net123
rlabel metal1 12742 2414 12742 2414 0 net124
rlabel metal2 20378 5882 20378 5882 0 net125
rlabel metal2 20654 5372 20654 5372 0 net126
rlabel metal1 23874 4182 23874 4182 0 net127
rlabel metal1 17526 5678 17526 5678 0 net128
rlabel metal1 21896 6290 21896 6290 0 net129
rlabel metal3 19619 18156 19619 18156 0 net13
rlabel metal1 20470 3162 20470 3162 0 net130
rlabel metal2 18906 4437 18906 4437 0 net131
rlabel metal1 18170 5678 18170 5678 0 net132
rlabel metal2 20654 7548 20654 7548 0 net133
rlabel metal1 22862 9554 22862 9554 0 net134
rlabel via3 17181 16660 17181 16660 0 net135
rlabel metal1 16836 15878 16836 15878 0 net136
rlabel metal1 14352 2414 14352 2414 0 net137
rlabel metal1 14490 3026 14490 3026 0 net138
rlabel metal1 16836 2414 16836 2414 0 net139
rlabel metal1 21482 22678 21482 22678 0 net14
rlabel metal1 16376 3502 16376 3502 0 net140
rlabel metal1 18308 13226 18308 13226 0 net141
rlabel metal1 17664 13158 17664 13158 0 net142
rlabel metal1 4646 53210 4646 53210 0 net143
rlabel metal2 6670 52836 6670 52836 0 net144
rlabel metal2 4830 52768 4830 52768 0 net145
rlabel metal1 8556 51510 8556 51510 0 net146
rlabel metal1 7866 51578 7866 51578 0 net147
rlabel metal2 9614 52326 9614 52326 0 net148
rlabel metal2 10718 51442 10718 51442 0 net149
rlabel metal1 26036 42602 26036 42602 0 net15
rlabel metal2 11730 51748 11730 51748 0 net150
rlabel metal1 18354 26010 18354 26010 0 net151
rlabel metal1 18308 27642 18308 27642 0 net152
rlabel metal1 24840 17510 24840 17510 0 net153
rlabel metal1 19780 28730 19780 28730 0 net154
rlabel metal1 24104 27642 24104 27642 0 net155
rlabel metal1 24150 28526 24150 28526 0 net156
rlabel metal1 21942 30226 21942 30226 0 net157
rlabel metal2 20194 30498 20194 30498 0 net158
rlabel metal1 19182 29138 19182 29138 0 net159
rlabel metal3 22241 41684 22241 41684 0 net16
rlabel metal1 22034 19278 22034 19278 0 net160
rlabel metal1 22954 16762 22954 16762 0 net161
rlabel metal1 19826 23834 19826 23834 0 net162
rlabel metal2 22218 21284 22218 21284 0 net163
rlabel metal1 7728 17306 7728 17306 0 net164
rlabel metal1 7314 12410 7314 12410 0 net165
rlabel metal1 8280 12886 8280 12886 0 net166
rlabel metal1 12420 17306 12420 17306 0 net167
rlabel metal1 13432 17306 13432 17306 0 net168
rlabel metal1 15824 16082 15824 16082 0 net169
rlabel metal2 22034 18530 22034 18530 0 net17
rlabel metal2 9890 21454 9890 21454 0 net170
rlabel metal2 12006 10234 12006 10234 0 net171
rlabel metal1 12926 6290 12926 6290 0 net172
rlabel metal2 14674 8092 14674 8092 0 net173
rlabel metal1 17296 14382 17296 14382 0 net174
rlabel metal1 14260 15130 14260 15130 0 net175
rlabel metal1 16008 17646 16008 17646 0 net176
rlabel metal1 15916 15130 15916 15130 0 net177
rlabel metal2 13386 8058 13386 8058 0 net178
rlabel metal1 15226 4794 15226 4794 0 net179
rlabel metal1 25070 44710 25070 44710 0 net18
rlabel metal2 19274 5916 19274 5916 0 net180
rlabel metal1 11500 21522 11500 21522 0 net181
rlabel metal1 13386 7378 13386 7378 0 net182
rlabel metal2 21298 10608 21298 10608 0 net183
rlabel metal2 19642 11526 19642 11526 0 net184
rlabel metal1 19734 12954 19734 12954 0 net185
rlabel metal2 21666 11526 21666 11526 0 net186
rlabel metal1 17250 9588 17250 9588 0 net187
rlabel metal1 24886 2618 24886 2618 0 net188
rlabel metal1 21206 2618 21206 2618 0 net189
rlabel metal1 25484 45798 25484 45798 0 net19
rlabel metal2 20010 9146 20010 9146 0 net190
rlabel metal1 11638 8466 11638 8466 0 net191
rlabel metal1 11822 19346 11822 19346 0 net192
rlabel metal2 9430 17476 9430 17476 0 net193
rlabel metal1 10948 12954 10948 12954 0 net194
rlabel metal2 11178 10200 11178 10200 0 net195
rlabel metal1 15502 23086 15502 23086 0 net196
rlabel metal1 15732 25874 15732 25874 0 net197
rlabel metal1 19734 21658 19734 21658 0 net198
rlabel metal1 24978 22032 24978 22032 0 net199
rlabel metal2 5382 4216 5382 4216 0 net2
rlabel metal1 25622 46342 25622 46342 0 net20
rlabel metal1 24472 24378 24472 24378 0 net200
rlabel metal2 20930 23562 20930 23562 0 net201
rlabel metal1 18722 24174 18722 24174 0 net202
rlabel metal1 25300 47430 25300 47430 0 net21
rlabel metal1 17434 16150 17434 16150 0 net22
rlabel metal3 16905 17476 16905 17476 0 net23
rlabel metal1 22310 49742 22310 49742 0 net24
rlabel metal1 25024 20910 25024 20910 0 net25
rlabel metal1 24978 23154 24978 23154 0 net26
rlabel metal1 22632 26010 22632 26010 0 net27
rlabel metal1 23874 26282 23874 26282 0 net28
rlabel metal1 25024 26418 25024 26418 0 net29
rlabel metal1 20608 13974 20608 13974 0 net3
rlabel metal1 25116 31926 25116 31926 0 net30
rlabel metal1 25530 33286 25530 33286 0 net31
rlabel metal1 21482 27098 21482 27098 0 net32
rlabel metal2 2254 6188 2254 6188 0 net33
rlabel metal1 13386 14246 13386 14246 0 net34
rlabel metal1 12834 13838 12834 13838 0 net35
rlabel metal1 7544 2278 7544 2278 0 net36
rlabel metal2 6762 5610 6762 5610 0 net37
rlabel metal1 13938 12818 13938 12818 0 net38
rlabel metal1 8096 2618 8096 2618 0 net39
rlabel metal1 24334 34714 24334 34714 0 net4
rlabel metal1 7866 2482 7866 2482 0 net40
rlabel metal1 15272 12886 15272 12886 0 net41
rlabel metal2 12742 5304 12742 5304 0 net42
rlabel metal1 12903 6698 12903 6698 0 net43
rlabel metal1 5750 17102 5750 17102 0 net44
rlabel metal1 15318 6630 15318 6630 0 net45
rlabel metal1 14076 10574 14076 10574 0 net46
rlabel metal1 9936 2618 9936 2618 0 net47
rlabel metal1 15180 9962 15180 9962 0 net48
rlabel metal1 17250 12716 17250 12716 0 net49
rlabel metal1 23920 17782 23920 17782 0 net5
rlabel metal1 17572 9010 17572 9010 0 net50
rlabel metal1 17710 13294 17710 13294 0 net51
rlabel metal1 16560 8806 16560 8806 0 net52
rlabel metal1 14444 2618 14444 2618 0 net53
rlabel metal1 14858 11696 14858 11696 0 net54
rlabel metal1 10212 18734 10212 18734 0 net55
rlabel metal1 4876 2618 4876 2618 0 net56
rlabel metal1 11868 19686 11868 19686 0 net57
rlabel metal1 1886 3604 1886 3604 0 net58
rlabel metal1 5658 12750 5658 12750 0 net59
rlabel metal1 24196 18394 24196 18394 0 net6
rlabel metal1 7406 12716 7406 12716 0 net60
rlabel metal1 12466 17204 12466 17204 0 net61
rlabel metal1 13478 17170 13478 17170 0 net62
rlabel metal1 12328 46478 12328 46478 0 net63
rlabel metal1 14628 47090 14628 47090 0 net64
rlabel metal2 16146 50286 16146 50286 0 net65
rlabel metal2 17710 49980 17710 49980 0 net66
rlabel metal1 19734 54196 19734 54196 0 net67
rlabel metal1 20983 17578 20983 17578 0 net68
rlabel metal1 21344 50694 21344 50694 0 net69
rlabel metal1 23138 13430 23138 13430 0 net7
rlabel metal2 24978 45540 24978 45540 0 net70
rlabel metal1 25668 52462 25668 52462 0 net71
rlabel metal1 17434 19482 17434 19482 0 net72
rlabel metal2 19642 21964 19642 21964 0 net73
rlabel metal1 20194 21998 20194 21998 0 net74
rlabel metal1 22264 52870 22264 52870 0 net75
rlabel metal1 17158 19414 17158 19414 0 net76
rlabel metal1 18814 33082 18814 33082 0 net77
rlabel metal1 19918 22066 19918 22066 0 net78
rlabel metal1 21022 54298 21022 54298 0 net79
rlabel metal3 23368 12716 23368 12716 0 net8
rlabel metal2 17250 20383 17250 20383 0 net80
rlabel metal1 22816 17102 22816 17102 0 net81
rlabel metal1 1794 53516 1794 53516 0 net82
rlabel metal2 9890 2210 9890 2210 0 net83
rlabel metal2 23506 6018 23506 6018 0 net84
rlabel metal1 24426 8058 24426 8058 0 net85
rlabel metal2 24610 10438 24610 10438 0 net86
rlabel metal1 22862 12240 22862 12240 0 net87
rlabel metal1 23460 13294 23460 13294 0 net88
rlabel metal1 22310 13940 22310 13940 0 net89
rlabel metal2 24932 32300 24932 32300 0 net9
rlabel metal2 24150 14076 24150 14076 0 net90
rlabel metal1 22310 12954 22310 12954 0 net91
rlabel metal1 22540 16558 22540 16558 0 net92
rlabel metal1 22264 15130 22264 15130 0 net93
rlabel metal1 15778 5100 15778 5100 0 net94
rlabel metal1 22632 17646 22632 17646 0 net95
rlabel metal2 24150 17884 24150 17884 0 net96
rlabel metal2 22678 19482 22678 19482 0 net97
rlabel metal1 21436 18938 21436 18938 0 net98
rlabel metal2 22126 20740 22126 20740 0 net99
rlabel metal1 23046 21114 23046 21114 0 prog_clk
rlabel metal1 23966 3026 23966 3026 0 prog_reset_bottom_in
rlabel metal2 24978 50711 24978 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 24978 51323 24978 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52275 24978 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25070 53669 25070 53669 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 23782 54077 23782 54077 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 24894 55420 24894 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 23391 56100 23391 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20562 56236 20562 56236 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21896 54162 21896 54162 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 23184 54162 23184 54162 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24564 54162 24564 54162 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 2062 1836 2062 1836 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 25116 20774 25116 20774 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 18630 46954 18630 46954 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 19412 21522 19412 21522 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 19366 17578 19366 17578 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal1 21666 19720 21666 19720 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal2 20194 18802 20194 18802 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 23092 21590 23092 21590 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 25300 24718 25300 24718 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 25070 23834 25070 23834 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 22678 26350 22678 26350 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal2 25254 26758 25254 26758 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20332 26418 20332 26418 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal2 22862 27676 22862 27676 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal2 19734 27200 19734 27200 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal1 21298 26860 21298 26860 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal2 18814 30192 18814 30192 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 18906 29172 18906 29172 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 18400 31994 18400 31994 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 17756 31858 17756 31858 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 19924 25162 19924 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal2 23874 20502 23874 20502 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal2 20930 29852 20930 29852 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal2 19090 32062 19090 32062 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 23644 30158 23644 30158 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 23138 31858 23138 31858 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 25024 32538 25024 32538 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24472 32334 24472 32334 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 22011 33898 22011 33898 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 22356 33422 22356 33422 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 20654 33286 20654 33286 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal1 19826 33592 19826 33592 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 21068 32198 21068 32198 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 33184 21206 33184 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal1 23460 21658 23460 21658 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 24472 21454 24472 21454 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 23644 18326 23644 18326 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 20838 24242 20838 24242 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 20010 23596 20010 23596 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 22310 25568 22310 25568 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 10856 26010 10856 26010 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 17526 31280 17526 31280 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 8648 17102 8648 17102 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal1 12466 22100 12466 22100 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8786 19142 8786 19142 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal1 10994 21318 10994 21318 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 9982 21658 9982 21658 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal2 10902 19244 10902 19244 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 9328 20026 9328 20026 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 13754 21454 13754 21454 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 12558 20978 12558 20978 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 14490 19754 14490 19754 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 14904 21454 14904 21454 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal1 14352 16626 14352 16626 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 14306 16762 14306 16762 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal1 11040 27098 11040 27098 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 15962 28594 15962 28594 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal2 13570 27030 13570 27030 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 10304 10982 10304 10982 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 10718 11186 10718 11186 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 10856 7514 10856 7514 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal2 10902 7616 10902 7616 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal2 12558 8160 12558 8160 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal2 11086 7072 11086 7072 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 15134 17102 15134 17102 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal1 14207 13702 14207 13702 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 15916 20026 15916 20026 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 14582 19720 14582 19720 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal2 17158 21182 17158 21182 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal2 17066 21590 17066 21590 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal2 18630 17884 18630 17884 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 17894 18190 17894 18190 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal1 16422 11254 16422 11254 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 17618 18802 17618 18802 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal2 14858 5780 14858 5780 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 13662 6868 13662 6868 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 17112 5270 17112 5270 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15502 5678 15502 5678 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13708 28390 13708 28390 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal1 16054 29682 16054 29682 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 14812 30022 14812 30022 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal1 18492 7310 18492 7310 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal2 17158 5678 17158 5678 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal1 21114 10574 21114 10574 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 19826 10710 19826 10710 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal2 20102 15470 20102 15470 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal1 19780 20978 19780 20978 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal1 22632 15538 22632 15538 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 21022 15878 21022 15878 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal2 23322 13566 23322 13566 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal1 21804 20978 21804 20978 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal1 24058 10574 24058 10574 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 22448 13362 22448 13362 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal2 24058 7344 24058 7344 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal2 22862 9690 22862 9690 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal2 21482 6018 21482 6018 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 19780 5134 19780 5134 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal2 20194 9248 20194 9248 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel via1 20003 8262 20003 8262 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 17480 19210 17480 19210 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 13340 24718 13340 24718 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 14398 29070 14398 29070 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 15870 26860 15870 26860 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal2 14766 24480 14766 24480 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal1 9154 17170 9154 17170 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 18768 14790 18768 14790 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20470 20400 20470 20400 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20148 16116 20148 16116 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 15962 10693 15962 10693 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24840 26554 24840 26554 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22816 19210 22816 19210 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 16456 20838 16456 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 23046 24786 23046 24786 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 20196 22218 20196 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18492 15878 18492 15878 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal1 21436 23834 21436 23834 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19964 16422 19964 16422 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17342 15878 17342 15878 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal2 18630 25500 18630 25500 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18216 16082 18216 16082 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16790 17510 16790 17510 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal2 18354 27846 18354 27846 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16928 17646 16928 17646 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 18598 15870 18598 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal2 18538 29648 18538 29648 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17687 18870 17687 18870 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18400 7854 18400 7854 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal1 25024 17714 25024 17714 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23736 17510 23736 17510 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18952 19686 18952 19686 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal1 20700 31994 20700 31994 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19044 19822 19044 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20976 18054 20976 18054 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 23230 31926 23230 31926 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22724 18190 22724 18190 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 18598 20838 18598 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 24104 33014 24104 33014 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21298 18734 21298 18734 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19136 18598 19136 18598 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal1 22632 34918 22632 34918 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 18666 20792 18666 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18354 13838 18354 13838 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 21160 35802 21160 35802 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19550 30022 19550 30022 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 21386 15226 21386 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 20332 35462 20332 35462 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15916 21522 15916 21522 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22080 3094 22080 3094 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 23644 19482 23644 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 19482 21528 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19918 13056 19918 13056 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal1 22770 17306 22770 17306 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20608 16966 20608 16966 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17986 16830 17986 16830 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 20378 23086 20378 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19918 23290 19918 23290 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18400 17238 18400 17238 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20148 14246 20148 14246 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22494 21386 22494 21386 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20102 21386 20102 21386 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21390 25262 21390 25262 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14858 31926 14858 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14306 28118 14306 28118 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12190 26316 12190 26316 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7590 17034 7590 17034 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13754 24922 13754 24922 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19458 19992 19458 19992 0 sb_0__8_.mux_right_track_10.out
rlabel metal1 13570 25160 13570 25160 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11730 23018 11730 23018 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10810 22950 10810 22950 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10212 17068 10212 17068 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12512 18122 12512 18122 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19366 19414 19366 19414 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12282 18666 12282 18666 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7912 18598 7912 18598 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16698 19380 16698 19380 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22770 20434 22770 20434 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15548 22134 15548 22134 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12328 17034 12328 17034 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17503 21522 17503 21522 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24196 18734 24196 18734 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 16192 24582 16192 24582 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 16966 14122 16966 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17802 19788 17802 19788 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19688 17306 19688 17306 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 14720 16218 14720 16218 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 17136 19090 17136 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 25500 20930 25500 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 14122 27438 14122 27438 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13616 27370 13616 27370 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 26656 12558 26656 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10994 21114 10994 21114 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17066 25908 17066 25908 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18354 12954 18354 12954 0 sb_0__8_.mux_right_track_20.out
rlabel metal1 11776 10098 11776 10098 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17848 12818 17848 12818 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17526 9792 17526 9792 0 sb_0__8_.mux_right_track_22.out
rlabel metal1 12190 7718 12190 7718 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13754 9044 13754 9044 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17342 11322 17342 11322 0 sb_0__8_.mux_right_track_24.out
rlabel metal2 14766 7616 14766 7616 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15088 8058 15088 8058 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22494 14042 22494 14042 0 sb_0__8_.mux_right_track_26.out
rlabel metal2 16698 13600 16698 13600 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20378 14110 20378 14110 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 17034 20930 17034 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 16192 19414 16192 19414 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13892 19482 13892 19482 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 19380 17526 19380 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21850 18122 21850 18122 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 17940 19822 17940 19822 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17894 18122 17894 18122 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19918 18258 19918 18258 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24794 13328 24794 13328 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 18124 23018 18124 23018 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18630 17578 18630 17578 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21482 17578 21482 17578 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23874 10642 23874 10642 0 sb_0__8_.mux_right_track_34.out
rlabel metal2 16882 14484 16882 14484 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12972 7718 12972 7718 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20654 11118 20654 11118 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14398 6732 14398 6732 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 14536 6358 14536 6358 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15318 6596 15318 6596 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23230 3332 23230 3332 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 15916 6698 15916 6698 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 3060 21482 3060 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19826 24446 19826 24446 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15640 29274 15640 29274 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 30158 15962 30158 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14628 26010 14628 26010 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10718 21896 10718 21896 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17802 25296 17802 25296 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12926 4556 12926 4556 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 17894 8602 17894 8602 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18676 8262 18676 8262 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16882 4760 16882 4760 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 21298 10098 21298 10098 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20930 9928 20930 9928 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 8942 23782 8942 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 19734 20842 19734 20842 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 14994 19642 14994 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 14858 20746 14858 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18446 10370 18446 10370 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 20194 21930 20194 21930 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18722 12920 18722 12920 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22172 14790 22172 14790 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23966 11322 23966 11322 0 sb_0__8_.mux_right_track_48.out
rlabel metal1 20976 21046 20976 21046 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20930 12818 20930 12818 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23920 12750 23920 12750 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18630 2312 18630 2312 0 sb_0__8_.mux_right_track_50.out
rlabel metal1 21022 13158 21022 13158 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23920 2414 23920 2414 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 2380 17526 2380 0 sb_0__8_.mux_right_track_52.out
rlabel metal2 21758 7888 21758 7888 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18998 6120 18998 6120 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17158 3706 17158 3706 0 sb_0__8_.mux_right_track_54.out
rlabel metal2 21022 6052 21022 6052 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18170 3706 18170 3706 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16192 5202 16192 5202 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 19780 9010 19780 9010 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19458 6630 19458 6630 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24702 6290 24702 6290 0 sb_0__8_.mux_right_track_58.out
rlabel metal2 16744 18700 16744 18700 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12098 12750 12098 12750 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 12614 17894 12614 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23644 21998 23644 21998 0 sb_0__8_.mux_right_track_6.out
rlabel metal2 15778 28016 15778 28016 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 27098 16284 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 25296 14950 25296 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12650 20026 12650 20026 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 23630 18262 23630 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19366 22746 19366 22746 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 13754 23562 13754 23562 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14122 23834 14122 23834 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12328 22066 12328 22066 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9200 17306 9200 17306 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11914 21896 11914 21896 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
